magic
tech sky130A
magscale 1 2
timestamp 1621206590
<< locali >>
rect 74733 19159 74767 19465
rect 43361 6647 43395 6749
rect 83105 5695 83139 5865
rect 85957 5627 85991 5797
rect 69213 5015 69247 5321
rect 13553 3995 13587 4165
rect 104725 3927 104759 4097
rect 10241 3383 10275 3689
rect 14197 3383 14231 3553
rect 24685 3451 24719 3689
rect 81081 3587 81115 3689
rect 9873 2975 9907 3077
rect 27261 2907 27295 3145
rect 48605 1615 48639 1989
rect 61209 1683 61243 2057
rect 77125 1479 77159 2057
rect 87061 1547 87095 1649
rect 88625 1547 88659 1853
rect 90281 1751 90315 2057
rect 90189 1547 90223 1717
<< viali >>
rect 2605 117249 2639 117283
rect 4537 117249 4571 117283
rect 7297 117249 7331 117283
rect 8677 117249 8711 117283
rect 12541 117249 12575 117283
rect 13553 117249 13587 117283
rect 16681 117249 16715 117283
rect 18245 117249 18279 117283
rect 21373 117249 21407 117283
rect 23213 117249 23247 117283
rect 26065 117249 26099 117283
rect 27353 117249 27387 117283
rect 31217 117249 31251 117283
rect 32321 117249 32355 117283
rect 35357 117249 35391 117283
rect 37013 117249 37047 117283
rect 40141 117249 40175 117283
rect 41889 117249 41923 117283
rect 44833 117249 44867 117283
rect 47225 117249 47259 117283
rect 49893 117249 49927 117283
rect 51089 117249 51123 117283
rect 54033 117249 54067 117283
rect 55781 117249 55815 117283
rect 58909 117249 58943 117283
rect 60565 117249 60599 117283
rect 63601 117249 63635 117283
rect 65901 117249 65935 117283
rect 68569 117249 68603 117283
rect 69857 117249 69891 117283
rect 72709 117249 72743 117283
rect 74549 117249 74583 117283
rect 77677 117249 77711 117283
rect 79241 117249 79275 117283
rect 82369 117249 82403 117283
rect 84577 117249 84611 117283
rect 87245 117249 87279 117283
rect 88625 117249 88659 117283
rect 92581 117249 92615 117283
rect 93409 117249 93443 117283
rect 96537 117249 96571 117283
rect 97825 117249 97859 117283
rect 101229 117249 101263 117283
rect 103253 117249 103287 117283
rect 105921 117249 105955 117283
rect 107393 117249 107427 117283
rect 111257 117249 111291 117283
rect 112177 117249 112211 117283
rect 115305 117249 115339 117283
rect 116869 117249 116903 117283
rect 119997 117249 120031 117283
rect 121929 117249 121963 117283
rect 124689 117249 124723 117283
rect 126069 117249 126103 117283
rect 129933 117249 129967 117283
rect 130945 117249 130979 117283
rect 134073 117249 134107 117283
rect 135637 117249 135671 117283
rect 138765 117249 138799 117283
rect 140605 117249 140639 117283
rect 143457 117249 143491 117283
rect 144745 117249 144779 117283
rect 148609 117249 148643 117283
rect 149713 117249 149747 117283
rect 152749 117249 152783 117283
rect 154405 117249 154439 117283
rect 157533 117249 157567 117283
rect 159281 117249 159315 117283
rect 162225 117249 162259 117283
rect 164617 117249 164651 117283
rect 167285 117249 167319 117283
rect 168481 117249 168515 117283
rect 171425 117249 171459 117283
rect 173173 117249 173207 117283
rect 176301 117249 176335 117283
rect 177957 117249 177991 117283
rect 1409 117181 1443 117215
rect 5457 117181 5491 117215
rect 10149 117181 10183 117215
rect 14933 117181 14967 117215
rect 20269 117181 20303 117215
rect 24225 117181 24259 117215
rect 28917 117181 28951 117215
rect 33609 117181 33643 117215
rect 35173 117181 35207 117215
rect 38945 117181 38979 117215
rect 42993 117181 43027 117215
rect 47685 117181 47719 117215
rect 52377 117181 52411 117215
rect 57621 117181 57655 117215
rect 61761 117181 61795 117215
rect 66453 117181 66487 117215
rect 71145 117181 71179 117215
rect 76297 117181 76331 117215
rect 80529 117181 80563 117215
rect 84393 117181 84427 117215
rect 85221 117181 85255 117215
rect 89913 117181 89947 117215
rect 94973 117181 95007 117215
rect 98009 117181 98043 117215
rect 99205 117181 99239 117215
rect 104081 117181 104115 117215
rect 108773 117181 108807 117215
rect 113649 117181 113683 117215
rect 118985 117181 119019 117215
rect 122849 117181 122883 117215
rect 127541 117181 127575 117215
rect 132325 117181 132359 117215
rect 137661 117181 137695 117215
rect 141617 117181 141651 117215
rect 146309 117181 146343 117215
rect 151001 117181 151035 117215
rect 156337 117181 156371 117215
rect 160385 117181 160419 117215
rect 165077 117181 165111 117215
rect 169769 117181 169803 117215
rect 173909 117181 173943 117215
rect 175565 117181 175599 117215
rect 2421 117113 2455 117147
rect 4353 117113 4387 117147
rect 7113 117113 7147 117147
rect 8493 117113 8527 117147
rect 12357 117113 12391 117147
rect 13369 117113 13403 117147
rect 16497 117113 16531 117147
rect 18061 117113 18095 117147
rect 21189 117113 21223 117147
rect 23029 117113 23063 117147
rect 25881 117113 25915 117147
rect 27169 117113 27203 117147
rect 31033 117113 31067 117147
rect 32137 117113 32171 117147
rect 36829 117113 36863 117147
rect 39957 117113 39991 117147
rect 41705 117113 41739 117147
rect 44649 117113 44683 117147
rect 47041 117113 47075 117147
rect 49709 117113 49743 117147
rect 50905 117113 50939 117147
rect 53849 117113 53883 117147
rect 55597 117113 55631 117147
rect 58725 117113 58759 117147
rect 60381 117113 60415 117147
rect 63417 117113 63451 117147
rect 65717 117113 65751 117147
rect 68385 117113 68419 117147
rect 69673 117113 69707 117147
rect 72525 117113 72559 117147
rect 74365 117113 74399 117147
rect 77493 117113 77527 117147
rect 79057 117113 79091 117147
rect 82185 117113 82219 117147
rect 87061 117113 87095 117147
rect 88441 117113 88475 117147
rect 92397 117113 92431 117147
rect 93225 117113 93259 117147
rect 96353 117113 96387 117147
rect 101045 117113 101079 117147
rect 103069 117113 103103 117147
rect 105737 117113 105771 117147
rect 107209 117113 107243 117147
rect 111073 117113 111107 117147
rect 111993 117113 112027 117147
rect 115121 117113 115155 117147
rect 116685 117113 116719 117147
rect 119813 117113 119847 117147
rect 121745 117113 121779 117147
rect 124505 117113 124539 117147
rect 125885 117113 125919 117147
rect 129749 117113 129783 117147
rect 130761 117113 130795 117147
rect 133889 117113 133923 117147
rect 135453 117113 135487 117147
rect 138581 117113 138615 117147
rect 140421 117113 140455 117147
rect 143273 117113 143307 117147
rect 144561 117113 144595 117147
rect 148425 117113 148459 117147
rect 149529 117113 149563 117147
rect 152565 117113 152599 117147
rect 154221 117113 154255 117147
rect 157349 117113 157383 117147
rect 159097 117113 159131 117147
rect 162041 117113 162075 117147
rect 164433 117113 164467 117147
rect 167101 117113 167135 117147
rect 168297 117113 168331 117147
rect 171241 117113 171275 117147
rect 172989 117113 173023 117147
rect 175381 117113 175415 117147
rect 176117 117113 176151 117147
rect 177773 117113 177807 117147
rect 97641 117045 97675 117079
rect 58265 116841 58299 116875
rect 158637 116841 158671 116875
rect 58449 116705 58483 116739
rect 158821 116705 158855 116739
rect 7941 116297 7975 116331
rect 12081 116297 12115 116331
rect 14749 116297 14783 116331
rect 18521 116297 18555 116331
rect 22569 116297 22603 116331
rect 26617 116297 26651 116331
rect 30849 116297 30883 116331
rect 35265 116297 35299 116331
rect 39773 116297 39807 116331
rect 44373 116297 44407 116331
rect 48973 116297 49007 116331
rect 54033 116297 54067 116331
rect 62957 116297 62991 116331
rect 77125 116297 77159 116331
rect 81817 116297 81851 116331
rect 86601 116297 86635 116331
rect 91385 116297 91419 116331
rect 96077 116297 96111 116331
rect 101229 116297 101263 116331
rect 105369 116297 105403 116331
rect 110245 116297 110279 116331
rect 114937 116297 114971 116331
rect 119629 116297 119663 116331
rect 124321 116297 124355 116331
rect 128921 116297 128955 116331
rect 133521 116297 133555 116331
rect 138029 116297 138063 116331
rect 143181 116297 143215 116331
rect 146769 116297 146803 116331
rect 150909 116297 150943 116331
rect 154129 116297 154163 116331
rect 154865 116297 154899 116331
rect 159097 116297 159131 116331
rect 162133 116297 162167 116331
rect 164341 116297 164375 116331
rect 168205 116297 168239 116331
rect 172897 116297 172931 116331
rect 176025 116297 176059 116331
rect 176945 116297 176979 116331
rect 177589 116297 177623 116331
rect 67649 116229 67683 116263
rect 72433 116229 72467 116263
rect 8125 116093 8159 116127
rect 12265 116093 12299 116127
rect 14933 116093 14967 116127
rect 18705 116093 18739 116127
rect 22753 116093 22787 116127
rect 26801 116093 26835 116127
rect 31033 116093 31067 116127
rect 35449 116093 35483 116127
rect 39957 116093 39991 116127
rect 44557 116093 44591 116127
rect 49157 116093 49191 116127
rect 54217 116093 54251 116127
rect 56793 116093 56827 116127
rect 57989 116093 58023 116127
rect 63141 116093 63175 116127
rect 67833 116093 67867 116127
rect 72617 116093 72651 116127
rect 77309 116093 77343 116127
rect 82001 116093 82035 116127
rect 86785 116093 86819 116127
rect 91569 116093 91603 116127
rect 96261 116093 96295 116127
rect 101413 116093 101447 116127
rect 105553 116093 105587 116127
rect 110429 116093 110463 116127
rect 115121 116093 115155 116127
rect 119813 116093 119847 116127
rect 124505 116093 124539 116127
rect 129105 116093 129139 116127
rect 133705 116093 133739 116127
rect 138213 116093 138247 116127
rect 143365 116093 143399 116127
rect 146953 116093 146987 116127
rect 151093 116093 151127 116127
rect 155049 116093 155083 116127
rect 162317 116093 162351 116127
rect 1869 60129 1903 60163
rect 177957 60129 177991 60163
rect 2053 59993 2087 60027
rect 178141 59993 178175 60027
rect 3065 59721 3099 59755
rect 176945 59721 176979 59755
rect 32781 24225 32815 24259
rect 32965 24225 32999 24259
rect 32873 24021 32907 24055
rect 26433 23137 26467 23171
rect 26617 23137 26651 23171
rect 26525 22933 26559 22967
rect 33149 22593 33183 22627
rect 33517 22525 33551 22559
rect 33634 22457 33668 22491
rect 33425 22389 33459 22423
rect 33793 22389 33827 22423
rect 29101 22117 29135 22151
rect 29306 22117 29340 22151
rect 29469 21913 29503 21947
rect 29285 21845 29319 21879
rect 27997 21437 28031 21471
rect 28089 21301 28123 21335
rect 29009 21029 29043 21063
rect 29193 20961 29227 20995
rect 29285 20961 29319 20995
rect 29009 20757 29043 20791
rect 28181 20417 28215 20451
rect 27997 20349 28031 20383
rect 28273 20349 28307 20383
rect 76113 20349 76147 20383
rect 27813 20213 27847 20247
rect 75745 20213 75779 20247
rect 76021 20213 76055 20247
rect 29101 20009 29135 20043
rect 29098 19873 29132 19907
rect 29469 19873 29503 19907
rect 31217 19873 31251 19907
rect 31401 19873 31435 19907
rect 29561 19805 29595 19839
rect 28917 19669 28951 19703
rect 31309 19669 31343 19703
rect 74733 19465 74767 19499
rect 75193 19465 75227 19499
rect 37013 19261 37047 19295
rect 37197 19261 37231 19295
rect 57161 19261 57195 19295
rect 59277 19261 59311 19295
rect 60197 19261 60231 19295
rect 61025 19261 61059 19295
rect 65257 19261 65291 19295
rect 73445 19261 73479 19295
rect 73353 19193 73387 19227
rect 75161 19193 75195 19227
rect 75331 19193 75365 19227
rect 37197 19125 37231 19159
rect 57253 19125 57287 19159
rect 59369 19125 59403 19159
rect 60289 19125 60323 19159
rect 61117 19125 61151 19159
rect 65349 19125 65383 19159
rect 73077 19125 73111 19159
rect 74733 19125 74767 19159
rect 74825 19125 74859 19159
rect 75009 19125 75043 19159
rect 75561 19125 75595 19159
rect 46857 18853 46891 18887
rect 47062 18853 47096 18887
rect 74181 18853 74215 18887
rect 74391 18853 74425 18887
rect 31769 18785 31803 18819
rect 42625 18785 42659 18819
rect 44005 18785 44039 18819
rect 66085 18785 66119 18819
rect 67833 18785 67867 18819
rect 68477 18785 68511 18819
rect 72433 18785 72467 18819
rect 73077 18785 73111 18819
rect 74089 18785 74123 18819
rect 74273 18785 74307 18819
rect 75009 18785 75043 18819
rect 75193 18785 75227 18819
rect 74549 18717 74583 18751
rect 75101 18717 75135 18751
rect 31953 18649 31987 18683
rect 46765 18649 46799 18683
rect 68569 18649 68603 18683
rect 73169 18649 73203 18683
rect 42717 18581 42751 18615
rect 44097 18581 44131 18615
rect 47041 18581 47075 18615
rect 47225 18581 47259 18615
rect 66177 18581 66211 18615
rect 67925 18581 67959 18615
rect 72525 18581 72559 18615
rect 73905 18581 73939 18615
rect 31861 18377 31895 18411
rect 31493 18241 31527 18275
rect 30665 18173 30699 18207
rect 30849 18173 30883 18207
rect 31677 18173 31711 18207
rect 31953 18173 31987 18207
rect 39129 18173 39163 18207
rect 39221 18173 39255 18207
rect 40785 18173 40819 18207
rect 41061 18173 41095 18207
rect 46121 18173 46155 18207
rect 49433 18173 49467 18207
rect 49617 18173 49651 18207
rect 54033 18173 54067 18207
rect 54217 18173 54251 18207
rect 72157 18173 72191 18207
rect 73537 18173 73571 18207
rect 30757 18105 30791 18139
rect 41153 18105 41187 18139
rect 54401 18105 54435 18139
rect 46213 18037 46247 18071
rect 49617 18037 49651 18071
rect 72249 18037 72283 18071
rect 73629 18037 73663 18071
rect 51549 17833 51583 17867
rect 60381 17765 60415 17799
rect 31769 17697 31803 17731
rect 37473 17697 37507 17731
rect 37749 17697 37783 17731
rect 51457 17697 51491 17731
rect 59461 17697 59495 17731
rect 59737 17697 59771 17731
rect 60197 17697 60231 17731
rect 37657 17629 37691 17663
rect 37289 17561 37323 17595
rect 59645 17561 59679 17595
rect 31861 17493 31895 17527
rect 59277 17493 59311 17527
rect 60565 17493 60599 17527
rect 45661 17289 45695 17323
rect 49433 17289 49467 17323
rect 59442 17289 59476 17323
rect 65882 17289 65916 17323
rect 67281 17289 67315 17323
rect 70041 17289 70075 17323
rect 72341 17289 72375 17323
rect 43729 17221 43763 17255
rect 57713 17221 57747 17255
rect 59553 17221 59587 17255
rect 64613 17221 64647 17255
rect 65993 17221 66027 17255
rect 59645 17153 59679 17187
rect 66085 17153 66119 17187
rect 34989 17085 35023 17119
rect 35265 17085 35299 17119
rect 35449 17085 35483 17119
rect 43637 17085 43671 17119
rect 43913 17085 43947 17119
rect 44373 17085 44407 17119
rect 45569 17085 45603 17119
rect 49249 17085 49283 17119
rect 49525 17085 49559 17119
rect 57621 17085 57655 17119
rect 57897 17085 57931 17119
rect 58357 17085 58391 17119
rect 64521 17085 64555 17119
rect 64797 17085 64831 17119
rect 65717 17085 65751 17119
rect 66913 17085 66947 17119
rect 67097 17085 67131 17119
rect 69857 17085 69891 17119
rect 70041 17085 70075 17119
rect 71145 17085 71179 17119
rect 71329 17085 71363 17119
rect 72249 17085 72283 17119
rect 73077 17085 73111 17119
rect 73261 17085 73295 17119
rect 73353 17085 73387 17119
rect 59277 17017 59311 17051
rect 65257 17017 65291 17051
rect 34805 16949 34839 16983
rect 49065 16949 49099 16983
rect 59921 16949 59955 16983
rect 66361 16949 66395 16983
rect 70225 16949 70259 16983
rect 71513 16949 71547 16983
rect 72893 16949 72927 16983
rect 32235 16745 32269 16779
rect 42901 16745 42935 16779
rect 32321 16677 32355 16711
rect 43821 16677 43855 16711
rect 59645 16677 59679 16711
rect 70409 16677 70443 16711
rect 32137 16609 32171 16643
rect 32413 16609 32447 16643
rect 40969 16609 41003 16643
rect 41153 16609 41187 16643
rect 42533 16609 42567 16643
rect 42993 16609 43027 16643
rect 43453 16609 43487 16643
rect 43637 16609 43671 16643
rect 46213 16609 46247 16643
rect 46397 16609 46431 16643
rect 47225 16609 47259 16643
rect 47409 16609 47443 16643
rect 47685 16609 47719 16643
rect 47869 16609 47903 16643
rect 52745 16609 52779 16643
rect 52929 16609 52963 16643
rect 53205 16609 53239 16643
rect 56701 16609 56735 16643
rect 56885 16609 56919 16643
rect 58541 16609 58575 16643
rect 58725 16609 58759 16643
rect 58817 16609 58851 16643
rect 59093 16609 59127 16643
rect 59553 16609 59587 16643
rect 65809 16609 65843 16643
rect 65993 16609 66027 16643
rect 68937 16609 68971 16643
rect 69121 16609 69155 16643
rect 70556 16609 70590 16643
rect 72433 16609 72467 16643
rect 72617 16609 72651 16643
rect 72893 16609 72927 16643
rect 73077 16609 73111 16643
rect 41337 16541 41371 16575
rect 41429 16541 41463 16575
rect 46305 16541 46339 16575
rect 53113 16541 53147 16575
rect 66269 16541 66303 16575
rect 70777 16541 70811 16575
rect 71145 16541 71179 16575
rect 70685 16473 70719 16507
rect 42717 16405 42751 16439
rect 56701 16405 56735 16439
rect 59001 16405 59035 16439
rect 66177 16405 66211 16439
rect 68937 16405 68971 16439
rect 32045 16201 32079 16235
rect 33241 16201 33275 16235
rect 33425 16201 33459 16235
rect 71145 16201 71179 16235
rect 71881 16201 71915 16235
rect 31493 16133 31527 16167
rect 44097 16133 44131 16167
rect 45845 16133 45879 16167
rect 57437 16065 57471 16099
rect 65717 16065 65751 16099
rect 31674 15997 31708 16031
rect 32137 15997 32171 16031
rect 44373 15997 44407 16031
rect 45845 15997 45879 16031
rect 46121 15997 46155 16031
rect 57253 15997 57287 16031
rect 57529 15997 57563 16031
rect 63417 15997 63451 16031
rect 63601 15997 63635 16031
rect 65441 15997 65475 16031
rect 65533 15997 65567 16031
rect 65809 15997 65843 16031
rect 66269 15997 66303 16031
rect 70317 15997 70351 16031
rect 70501 15997 70535 16031
rect 70685 15997 70719 16031
rect 71421 15997 71455 16031
rect 71881 15997 71915 16031
rect 72065 15997 72099 16031
rect 33057 15929 33091 15963
rect 44097 15929 44131 15963
rect 44281 15929 44315 15963
rect 46029 15929 46063 15963
rect 66361 15929 66395 15963
rect 71145 15929 71179 15963
rect 71329 15929 71363 15963
rect 31677 15861 31711 15895
rect 33262 15861 33296 15895
rect 57069 15861 57103 15895
rect 63509 15861 63543 15895
rect 65257 15861 65291 15895
rect 29285 15657 29319 15691
rect 31953 15657 31987 15691
rect 56885 15657 56919 15691
rect 62681 15657 62715 15691
rect 70225 15657 70259 15691
rect 71145 15657 71179 15691
rect 56701 15589 56735 15623
rect 62497 15589 62531 15623
rect 70961 15589 70995 15623
rect 29193 15521 29227 15555
rect 31861 15521 31895 15555
rect 33701 15521 33735 15555
rect 33885 15521 33919 15555
rect 56977 15521 57011 15555
rect 62773 15521 62807 15555
rect 63877 15521 63911 15555
rect 64061 15521 64095 15555
rect 64153 15521 64187 15555
rect 69121 15521 69155 15555
rect 69857 15521 69891 15555
rect 70317 15521 70351 15555
rect 71237 15521 71271 15555
rect 29469 15453 29503 15487
rect 32045 15453 32079 15487
rect 69305 15453 69339 15487
rect 69397 15453 69431 15487
rect 28825 15317 28859 15351
rect 31493 15317 31527 15351
rect 33701 15317 33735 15351
rect 56701 15317 56735 15351
rect 62497 15317 62531 15351
rect 63693 15317 63727 15351
rect 68937 15317 68971 15351
rect 70041 15317 70075 15351
rect 70961 15317 70995 15351
rect 30665 15045 30699 15079
rect 31125 14977 31159 15011
rect 31217 14977 31251 15011
rect 65993 14977 66027 15011
rect 33517 14909 33551 14943
rect 33793 14909 33827 14943
rect 59921 14909 59955 14943
rect 65809 14909 65843 14943
rect 68385 14909 68419 14943
rect 35173 14841 35207 14875
rect 59737 14841 59771 14875
rect 60105 14841 60139 14875
rect 65625 14841 65659 14875
rect 68109 14841 68143 14875
rect 31033 14773 31067 14807
rect 68207 14773 68241 14807
rect 68293 14773 68327 14807
rect 33241 14569 33275 14603
rect 68661 14569 68695 14603
rect 31861 14501 31895 14535
rect 34069 14501 34103 14535
rect 46857 14501 46891 14535
rect 69857 14501 69891 14535
rect 31125 14433 31159 14467
rect 33149 14433 33183 14467
rect 68569 14433 68603 14467
rect 69765 14433 69799 14467
rect 33425 14365 33459 14399
rect 68845 14365 68879 14399
rect 70041 14365 70075 14399
rect 34253 14297 34287 14331
rect 32781 14229 32815 14263
rect 46949 14229 46983 14263
rect 68201 14229 68235 14263
rect 69397 14229 69431 14263
rect 30481 14025 30515 14059
rect 40693 14025 40727 14059
rect 46857 14025 46891 14059
rect 60565 14025 60599 14059
rect 65073 14025 65107 14059
rect 33425 13957 33459 13991
rect 35909 13957 35943 13991
rect 38393 13957 38427 13991
rect 48789 13957 48823 13991
rect 59277 13957 59311 13991
rect 66269 13957 66303 13991
rect 68109 13957 68143 13991
rect 69765 13957 69799 13991
rect 29101 13889 29135 13923
rect 33885 13889 33919 13923
rect 34069 13889 34103 13923
rect 36369 13889 36403 13923
rect 36461 13889 36495 13923
rect 38853 13889 38887 13923
rect 39037 13889 39071 13923
rect 41153 13889 41187 13923
rect 41337 13889 41371 13923
rect 44925 13889 44959 13923
rect 47317 13889 47351 13923
rect 47501 13889 47535 13923
rect 49249 13889 49283 13923
rect 49433 13889 49467 13923
rect 59737 13889 59771 13923
rect 59921 13889 59955 13923
rect 61209 13889 61243 13923
rect 65533 13889 65567 13923
rect 65717 13889 65751 13923
rect 66821 13889 66855 13923
rect 68753 13889 68787 13923
rect 70317 13889 70351 13923
rect 29377 13821 29411 13855
rect 39681 13821 39715 13855
rect 39865 13821 39899 13855
rect 44741 13821 44775 13855
rect 55229 13821 55263 13855
rect 55413 13821 55447 13855
rect 56977 13821 57011 13855
rect 61025 13821 61059 13855
rect 66729 13821 66763 13855
rect 68569 13821 68603 13855
rect 70133 13821 70167 13855
rect 70225 13821 70259 13855
rect 36277 13753 36311 13787
rect 38761 13753 38795 13787
rect 41061 13753 41095 13787
rect 47225 13753 47259 13787
rect 33793 13685 33827 13719
rect 49157 13685 49191 13719
rect 56793 13685 56827 13719
rect 59645 13685 59679 13719
rect 60933 13685 60967 13719
rect 65441 13685 65475 13719
rect 66637 13685 66671 13719
rect 68477 13685 68511 13719
rect 32229 13481 32263 13515
rect 33425 13481 33459 13515
rect 43545 13481 43579 13515
rect 44741 13481 44775 13515
rect 47593 13481 47627 13515
rect 51917 13481 51951 13515
rect 55321 13481 55355 13515
rect 57621 13481 57655 13515
rect 63325 13481 63359 13515
rect 71237 13481 71271 13515
rect 42625 13413 42659 13447
rect 43453 13413 43487 13447
rect 44649 13413 44683 13447
rect 30849 13345 30883 13379
rect 33149 13345 33183 13379
rect 33609 13345 33643 13379
rect 33977 13345 34011 13379
rect 46213 13345 46247 13379
rect 48513 13345 48547 13379
rect 51825 13345 51859 13379
rect 55229 13345 55263 13379
rect 57529 13345 57563 13379
rect 58633 13345 58667 13379
rect 63233 13345 63267 13379
rect 69489 13345 69523 13379
rect 71145 13345 71179 13379
rect 31125 13277 31159 13311
rect 33057 13277 33091 13311
rect 36277 13277 36311 13311
rect 36553 13277 36587 13311
rect 40969 13277 41003 13311
rect 41245 13277 41279 13311
rect 43637 13277 43671 13311
rect 44833 13277 44867 13311
rect 46489 13277 46523 13311
rect 48881 13277 48915 13311
rect 52101 13277 52135 13311
rect 55505 13277 55539 13311
rect 57805 13277 57839 13311
rect 58357 13277 58391 13311
rect 60013 13277 60047 13311
rect 63417 13277 63451 13311
rect 64613 13277 64647 13311
rect 64889 13277 64923 13311
rect 67189 13277 67223 13311
rect 67465 13277 67499 13311
rect 70133 13277 70167 13311
rect 71421 13277 71455 13311
rect 43085 13209 43119 13243
rect 37657 13141 37691 13175
rect 44281 13141 44315 13175
rect 51457 13141 51491 13175
rect 54861 13141 54895 13175
rect 57161 13141 57195 13175
rect 62865 13141 62899 13175
rect 66177 13141 66211 13175
rect 68753 13141 68787 13175
rect 70777 13141 70811 13175
rect 32045 12937 32079 12971
rect 34621 12937 34655 12971
rect 36829 12937 36863 12971
rect 39865 12937 39899 12971
rect 41981 12937 42015 12971
rect 45661 12937 45695 12971
rect 56425 12937 56459 12971
rect 61669 12937 61703 12971
rect 69765 12937 69799 12971
rect 30481 12801 30515 12835
rect 33057 12801 33091 12835
rect 35449 12801 35483 12835
rect 38485 12801 38519 12835
rect 40601 12801 40635 12835
rect 44281 12801 44315 12835
rect 46857 12801 46891 12835
rect 47041 12801 47075 12835
rect 49065 12801 49099 12835
rect 54861 12801 54895 12835
rect 57437 12801 57471 12835
rect 57621 12801 57655 12835
rect 59553 12801 59587 12835
rect 62313 12801 62347 12835
rect 63417 12801 63451 12835
rect 66637 12801 66671 12835
rect 68293 12801 68327 12835
rect 70363 12801 70397 12835
rect 30757 12733 30791 12767
rect 33333 12733 33367 12767
rect 35725 12733 35759 12767
rect 38761 12733 38795 12767
rect 40877 12733 40911 12767
rect 44557 12733 44591 12767
rect 46765 12733 46799 12767
rect 48789 12733 48823 12767
rect 50905 12733 50939 12767
rect 51181 12733 51215 12767
rect 55137 12733 55171 12767
rect 59829 12733 59863 12767
rect 62037 12733 62071 12767
rect 62129 12733 62163 12767
rect 64521 12733 64555 12767
rect 64797 12733 64831 12767
rect 66913 12733 66947 12767
rect 70133 12733 70167 12767
rect 50445 12665 50479 12699
rect 61209 12665 61243 12699
rect 63325 12665 63359 12699
rect 70225 12665 70259 12699
rect 46397 12597 46431 12631
rect 52285 12597 52319 12631
rect 56977 12597 57011 12631
rect 57345 12597 57379 12631
rect 62865 12597 62899 12631
rect 63233 12597 63267 12631
rect 66085 12597 66119 12631
rect 36185 12393 36219 12427
rect 38393 12393 38427 12427
rect 60381 12393 60415 12427
rect 36093 12257 36127 12291
rect 37013 12257 37047 12291
rect 46857 12257 46891 12291
rect 56701 12257 56735 12291
rect 59093 12257 59127 12291
rect 36369 12189 36403 12223
rect 37289 12189 37323 12223
rect 47133 12189 47167 12223
rect 56977 12189 57011 12223
rect 61945 12189 61979 12223
rect 62221 12189 62255 12223
rect 64061 12189 64095 12223
rect 64337 12189 64371 12223
rect 67281 12189 67315 12223
rect 67557 12189 67591 12223
rect 69397 12189 69431 12223
rect 69673 12189 69707 12223
rect 35725 12053 35759 12087
rect 48421 12053 48455 12087
rect 58081 12053 58115 12087
rect 63509 12053 63543 12087
rect 65441 12053 65475 12087
rect 68661 12053 68695 12087
rect 70961 12053 70995 12087
rect 61669 11849 61703 11883
rect 59277 11713 59311 11747
rect 65349 11713 65383 11747
rect 67465 11713 67499 11747
rect 59553 11645 59587 11679
rect 61853 11645 61887 11679
rect 65073 11645 65107 11679
rect 67189 11645 67223 11679
rect 60841 11509 60875 11543
rect 66453 11509 66487 11543
rect 68569 11509 68603 11543
rect 68937 11305 68971 11339
rect 67373 11169 67407 11203
rect 67649 11101 67683 11135
rect 33425 10761 33459 10795
rect 34529 10761 34563 10795
rect 33241 10557 33275 10591
rect 34345 10557 34379 10591
rect 60381 10557 60415 10591
rect 60657 10557 60691 10591
rect 33057 10489 33091 10523
rect 34161 10489 34195 10523
rect 31401 10149 31435 10183
rect 31769 10149 31803 10183
rect 32965 10149 32999 10183
rect 33793 10149 33827 10183
rect 39957 10149 39991 10183
rect 41613 10149 41647 10183
rect 45293 10149 45327 10183
rect 46581 10149 46615 10183
rect 47961 10149 47995 10183
rect 62773 10149 62807 10183
rect 66269 10149 66303 10183
rect 31585 10081 31619 10115
rect 32597 10081 32631 10115
rect 32781 10081 32815 10115
rect 33425 10081 33459 10115
rect 33609 10081 33643 10115
rect 39589 10081 39623 10115
rect 39773 10081 39807 10115
rect 41245 10081 41279 10115
rect 41429 10081 41463 10115
rect 44925 10081 44959 10115
rect 45109 10081 45143 10115
rect 46213 10081 46247 10115
rect 46397 10081 46431 10115
rect 47593 10081 47627 10115
rect 47777 10081 47811 10115
rect 56701 10081 56735 10115
rect 58725 10081 58759 10115
rect 62405 10081 62439 10115
rect 62589 10081 62623 10115
rect 65901 10081 65935 10115
rect 66085 10081 66119 10115
rect 58909 9945 58943 9979
rect 56885 9877 56919 9911
rect 37381 9605 37415 9639
rect 38669 9605 38703 9639
rect 40877 9605 40911 9639
rect 42441 9605 42475 9639
rect 47225 9605 47259 9639
rect 49157 9605 49191 9639
rect 55229 9605 55263 9639
rect 57437 9605 57471 9639
rect 58357 9605 58391 9639
rect 56609 9537 56643 9571
rect 63601 9537 63635 9571
rect 65625 9537 65659 9571
rect 66453 9537 66487 9571
rect 67281 9537 67315 9571
rect 37197 9469 37231 9503
rect 38485 9469 38519 9503
rect 40693 9469 40727 9503
rect 42257 9469 42291 9503
rect 47041 9469 47075 9503
rect 48973 9469 49007 9503
rect 55045 9469 55079 9503
rect 56425 9469 56459 9503
rect 57253 9469 57287 9503
rect 58173 9469 58207 9503
rect 62037 9469 62071 9503
rect 63417 9469 63451 9503
rect 65441 9469 65475 9503
rect 66269 9469 66303 9503
rect 67097 9469 67131 9503
rect 37013 9401 37047 9435
rect 38301 9401 38335 9435
rect 40509 9401 40543 9435
rect 42073 9401 42107 9435
rect 46857 9401 46891 9435
rect 48789 9401 48823 9435
rect 54861 9401 54895 9435
rect 56241 9401 56275 9435
rect 57069 9401 57103 9435
rect 57989 9401 58023 9435
rect 61853 9401 61887 9435
rect 62221 9401 62255 9435
rect 63233 9401 63267 9435
rect 65257 9401 65291 9435
rect 66085 9401 66119 9435
rect 66913 9401 66947 9435
rect 32781 9061 32815 9095
rect 63693 9061 63727 9095
rect 65993 9061 66027 9095
rect 32597 8993 32631 9027
rect 32873 8993 32907 9027
rect 32965 8993 32999 9027
rect 55413 8993 55447 9027
rect 55597 8993 55631 9027
rect 60565 8993 60599 9027
rect 60749 8993 60783 9027
rect 61945 8993 61979 9027
rect 62129 8993 62163 9027
rect 63325 8993 63359 9027
rect 63509 8993 63543 9027
rect 65625 8993 65659 9027
rect 65809 8993 65843 9027
rect 55781 8925 55815 8959
rect 60933 8925 60967 8959
rect 62313 8925 62347 8959
rect 33149 8789 33183 8823
rect 41429 8585 41463 8619
rect 33793 8517 33827 8551
rect 33241 8381 33275 8415
rect 33425 8381 33459 8415
rect 33609 8381 33643 8415
rect 35173 8381 35207 8415
rect 35357 8381 35391 8415
rect 40877 8381 40911 8415
rect 41061 8381 41095 8415
rect 41153 8381 41187 8415
rect 41245 8381 41279 8415
rect 45937 8381 45971 8415
rect 46121 8381 46155 8415
rect 46305 8381 46339 8415
rect 33517 8313 33551 8347
rect 35909 8313 35943 8347
rect 36093 8313 36127 8347
rect 46213 8313 46247 8347
rect 46489 8245 46523 8279
rect 33609 8041 33643 8075
rect 33793 8041 33827 8075
rect 64429 8041 64463 8075
rect 21005 7973 21039 8007
rect 21097 7973 21131 8007
rect 25789 7973 25823 8007
rect 27813 7973 27847 8007
rect 30665 7973 30699 8007
rect 31861 7973 31895 8007
rect 32505 7973 32539 8007
rect 32781 7973 32815 8007
rect 33241 7973 33275 8007
rect 38301 7973 38335 8007
rect 39681 7973 39715 8007
rect 41889 7973 41923 8007
rect 41981 7973 42015 8007
rect 48605 7973 48639 8007
rect 48697 7973 48731 8007
rect 20821 7905 20855 7939
rect 21189 7905 21223 7939
rect 25605 7905 25639 7939
rect 25881 7905 25915 7939
rect 25973 7905 26007 7939
rect 27629 7905 27663 7939
rect 27905 7905 27939 7939
rect 27997 7905 28031 7939
rect 28733 7905 28767 7939
rect 30481 7905 30515 7939
rect 30757 7905 30791 7939
rect 30849 7905 30883 7939
rect 31677 7905 31711 7939
rect 32873 7905 32907 7939
rect 36461 7905 36495 7939
rect 39497 7905 39531 7939
rect 39773 7905 39807 7939
rect 39865 7905 39899 7939
rect 40969 7905 41003 7939
rect 41705 7905 41739 7939
rect 42073 7905 42107 7939
rect 44557 7905 44591 7939
rect 46397 7905 46431 7939
rect 46581 7905 46615 7939
rect 46673 7905 46707 7939
rect 46811 7905 46845 7939
rect 47409 7905 47443 7939
rect 47547 7905 47581 7939
rect 47685 7905 47719 7939
rect 47777 7905 47811 7939
rect 48421 7905 48455 7939
rect 48789 7905 48823 7939
rect 62589 7905 62623 7939
rect 63527 7905 63561 7939
rect 63626 7905 63660 7939
rect 28917 7837 28951 7871
rect 36645 7837 36679 7871
rect 62773 7837 62807 7871
rect 63785 7837 63819 7871
rect 38485 7769 38519 7803
rect 41153 7769 41187 7803
rect 63233 7769 63267 7803
rect 21373 7701 21407 7735
rect 26157 7701 26191 7735
rect 28181 7701 28215 7735
rect 31033 7701 31067 7735
rect 40049 7701 40083 7735
rect 42257 7701 42291 7735
rect 44373 7701 44407 7735
rect 46949 7701 46983 7735
rect 47961 7701 47995 7735
rect 48973 7701 49007 7735
rect 29653 7497 29687 7531
rect 35817 7497 35851 7531
rect 40877 7497 40911 7531
rect 56701 7497 56735 7531
rect 61485 7497 61519 7531
rect 64613 7497 64647 7531
rect 31033 7429 31067 7463
rect 44189 7429 44223 7463
rect 46397 7429 46431 7463
rect 45017 7361 45051 7395
rect 54861 7361 54895 7395
rect 55045 7361 55079 7395
rect 55505 7361 55539 7395
rect 55919 7361 55953 7395
rect 62267 7361 62301 7395
rect 62681 7361 62715 7395
rect 63325 7361 63359 7395
rect 18613 7293 18647 7327
rect 18797 7293 18831 7327
rect 18981 7293 19015 7327
rect 20177 7293 20211 7327
rect 20361 7293 20395 7327
rect 20545 7293 20579 7327
rect 23029 7293 23063 7327
rect 23305 7293 23339 7327
rect 23397 7293 23431 7327
rect 26341 7293 26375 7327
rect 26525 7293 26559 7327
rect 26709 7293 26743 7327
rect 28457 7293 28491 7327
rect 28595 7293 28629 7327
rect 28871 7293 28905 7327
rect 30941 7293 30975 7327
rect 31217 7293 31251 7327
rect 33333 7293 33367 7327
rect 33517 7293 33551 7327
rect 33701 7293 33735 7327
rect 34897 7293 34931 7327
rect 35265 7293 35299 7327
rect 36369 7293 36403 7327
rect 36553 7293 36587 7327
rect 36737 7293 36771 7327
rect 38301 7293 38335 7327
rect 38485 7293 38519 7327
rect 38669 7293 38703 7327
rect 39221 7293 39255 7327
rect 41705 7293 41739 7327
rect 41889 7293 41923 7327
rect 42073 7293 42107 7327
rect 43637 7293 43671 7327
rect 43913 7293 43947 7327
rect 44005 7293 44039 7327
rect 45284 7293 45318 7327
rect 47041 7293 47075 7327
rect 48789 7293 48823 7327
rect 48973 7293 49007 7327
rect 49157 7293 49191 7327
rect 49801 7293 49835 7327
rect 49985 7293 50019 7327
rect 50169 7293 50203 7327
rect 55799 7293 55833 7327
rect 56057 7293 56091 7327
rect 62129 7293 62163 7327
rect 62386 7293 62420 7327
rect 63141 7293 63175 7327
rect 18889 7225 18923 7259
rect 20453 7225 20487 7259
rect 23213 7225 23247 7259
rect 24869 7225 24903 7259
rect 26617 7225 26651 7259
rect 28733 7225 28767 7259
rect 29561 7225 29595 7259
rect 33609 7225 33643 7259
rect 34483 7225 34517 7259
rect 34805 7225 34839 7259
rect 36645 7225 36679 7259
rect 38577 7225 38611 7259
rect 39589 7225 39623 7259
rect 39865 7225 39899 7259
rect 39957 7225 39991 7259
rect 40325 7225 40359 7259
rect 40693 7225 40727 7259
rect 41981 7225 42015 7259
rect 43821 7225 43855 7259
rect 47685 7225 47719 7259
rect 49065 7225 49099 7259
rect 50077 7225 50111 7259
rect 65165 7225 65199 7259
rect 65533 7225 65567 7259
rect 65625 7225 65659 7259
rect 19165 7157 19199 7191
rect 20729 7157 20763 7191
rect 23581 7157 23615 7191
rect 24961 7157 24995 7191
rect 26893 7157 26927 7191
rect 29009 7157 29043 7191
rect 31401 7157 31435 7191
rect 33885 7157 33919 7191
rect 34161 7157 34195 7191
rect 35633 7157 35667 7191
rect 36921 7157 36955 7191
rect 38853 7157 38887 7191
rect 42257 7157 42291 7191
rect 49341 7157 49375 7191
rect 50353 7157 50387 7191
rect 61393 7157 61427 7191
rect 64429 7157 64463 7191
rect 64797 7157 64831 7191
rect 65901 7157 65935 7191
rect 21097 6953 21131 6987
rect 41153 6953 41187 6987
rect 63509 6953 63543 6987
rect 21741 6885 21775 6919
rect 31401 6885 31435 6919
rect 31656 6885 31690 6919
rect 31769 6885 31803 6919
rect 32505 6885 32539 6919
rect 33425 6885 33459 6919
rect 34529 6885 34563 6919
rect 39773 6885 39807 6919
rect 42257 6885 42291 6919
rect 46765 6885 46799 6919
rect 50169 6885 50203 6919
rect 16672 6817 16706 6851
rect 18521 6817 18555 6851
rect 18705 6817 18739 6851
rect 18797 6817 18831 6851
rect 18889 6817 18923 6851
rect 20545 6817 20579 6851
rect 20729 6817 20763 6851
rect 20821 6817 20855 6851
rect 20913 6817 20947 6851
rect 21557 6817 21591 6851
rect 21829 6817 21863 6851
rect 21949 6817 21983 6851
rect 25513 6817 25547 6851
rect 28549 6817 28583 6851
rect 29377 6817 29411 6851
rect 30573 6817 30607 6851
rect 32137 6817 32171 6851
rect 33701 6817 33735 6851
rect 33793 6817 33827 6851
rect 34161 6817 34195 6851
rect 36001 6817 36035 6851
rect 36645 6817 36679 6851
rect 37682 6817 37716 6851
rect 39589 6817 39623 6851
rect 41429 6817 41463 6851
rect 41521 6817 41555 6851
rect 41889 6817 41923 6851
rect 44490 6817 44524 6851
rect 44649 6817 44683 6851
rect 45293 6817 45327 6851
rect 46489 6817 46523 6851
rect 46673 6817 46707 6851
rect 46857 6817 46891 6851
rect 48630 6817 48664 6851
rect 49433 6817 49467 6851
rect 49893 6817 49927 6851
rect 50077 6817 50111 6851
rect 50261 6817 50295 6851
rect 52837 6817 52871 6851
rect 53481 6817 53515 6851
rect 54978 6817 55012 6851
rect 55781 6817 55815 6851
rect 57069 6817 57103 6851
rect 59185 6817 59219 6851
rect 60105 6817 60139 6851
rect 62129 6817 62163 6851
rect 62957 6817 62991 6851
rect 63693 6817 63727 6851
rect 65533 6817 65567 6851
rect 80529 6817 80563 6851
rect 82921 6817 82955 6851
rect 16405 6749 16439 6783
rect 36829 6749 36863 6783
rect 37289 6749 37323 6783
rect 37565 6749 37599 6783
rect 37841 6749 37875 6783
rect 38485 6749 38519 6783
rect 43361 6749 43395 6783
rect 43453 6749 43487 6783
rect 43637 6749 43671 6783
rect 44373 6749 44407 6783
rect 47593 6749 47627 6783
rect 47777 6749 47811 6783
rect 48513 6749 48547 6783
rect 48789 6749 48823 6783
rect 51641 6749 51675 6783
rect 51825 6749 51859 6783
rect 52561 6749 52595 6783
rect 52699 6749 52733 6783
rect 53941 6749 53975 6783
rect 54125 6749 54159 6783
rect 54861 6749 54895 6783
rect 55137 6749 55171 6783
rect 58909 6749 58943 6783
rect 59047 6749 59081 6783
rect 59921 6749 59955 6783
rect 64337 6749 64371 6783
rect 64475 6749 64509 6783
rect 64613 6749 64647 6783
rect 65349 6749 65383 6783
rect 22109 6681 22143 6715
rect 25697 6681 25731 6715
rect 32689 6681 32723 6715
rect 34713 6681 34747 6715
rect 36185 6681 36219 6715
rect 42441 6681 42475 6715
rect 44097 6681 44131 6715
rect 48237 6681 48271 6715
rect 52285 6681 52319 6715
rect 54585 6681 54619 6715
rect 59461 6681 59495 6715
rect 64889 6681 64923 6715
rect 17785 6613 17819 6647
rect 19073 6613 19107 6647
rect 28641 6613 28675 6647
rect 29469 6613 29503 6647
rect 30665 6613 30699 6647
rect 31033 6613 31067 6647
rect 36461 6613 36495 6647
rect 43361 6613 43395 6647
rect 47041 6613 47075 6647
rect 50445 6613 50479 6647
rect 56885 6613 56919 6647
rect 58081 6613 58115 6647
rect 58265 6613 58299 6647
rect 61945 6613 61979 6647
rect 62773 6613 62807 6647
rect 80713 6613 80747 6647
rect 83105 6613 83139 6647
rect 34529 6409 34563 6443
rect 37381 6409 37415 6443
rect 39773 6409 39807 6443
rect 42533 6409 42567 6443
rect 45569 6409 45603 6443
rect 57989 6409 58023 6443
rect 61117 6409 61151 6443
rect 83657 6409 83691 6443
rect 29193 6341 29227 6375
rect 31309 6341 31343 6375
rect 46029 6341 46063 6375
rect 47225 6341 47259 6375
rect 62957 6341 62991 6375
rect 64521 6341 64555 6375
rect 80897 6341 80931 6375
rect 35541 6273 35575 6307
rect 36185 6273 36219 6307
rect 36578 6273 36612 6307
rect 36737 6273 36771 6307
rect 43729 6273 43763 6307
rect 43913 6273 43947 6307
rect 44373 6273 44407 6307
rect 44787 6273 44821 6307
rect 46673 6273 46707 6307
rect 46832 6273 46866 6307
rect 47869 6273 47903 6307
rect 56149 6273 56183 6307
rect 56793 6273 56827 6307
rect 57207 6273 57241 6307
rect 57345 6273 57379 6307
rect 59277 6273 59311 6307
rect 59921 6273 59955 6307
rect 60197 6273 60231 6307
rect 60473 6273 60507 6307
rect 62405 6273 62439 6307
rect 62564 6273 62598 6307
rect 63417 6273 63451 6307
rect 64429 6273 64463 6307
rect 65165 6273 65199 6307
rect 65324 6273 65358 6307
rect 65717 6273 65751 6307
rect 66361 6273 66395 6307
rect 82369 6273 82403 6307
rect 17325 6205 17359 6239
rect 17592 6205 17626 6239
rect 19165 6205 19199 6239
rect 19432 6205 19466 6239
rect 21005 6205 21039 6239
rect 21281 6205 21315 6239
rect 21373 6205 21407 6239
rect 23765 6205 23799 6239
rect 24032 6205 24066 6239
rect 27813 6205 27847 6239
rect 33977 6205 34011 6239
rect 35725 6205 35759 6239
rect 36461 6205 36495 6239
rect 39221 6205 39255 6239
rect 41981 6205 42015 6239
rect 44649 6205 44683 6239
rect 44925 6205 44959 6239
rect 46949 6205 46983 6239
rect 47685 6205 47719 6239
rect 48789 6205 48823 6239
rect 49061 6205 49095 6239
rect 49203 6205 49237 6239
rect 49985 6205 50019 6239
rect 50629 6205 50663 6239
rect 51273 6205 51307 6239
rect 54225 6205 54259 6239
rect 56333 6205 56367 6239
rect 57069 6205 57103 6239
rect 59461 6205 59495 6239
rect 60335 6205 60369 6239
rect 61761 6205 61795 6239
rect 62681 6205 62715 6239
rect 63601 6205 63635 6239
rect 65441 6205 65475 6239
rect 66177 6205 66211 6239
rect 67005 6205 67039 6239
rect 68109 6205 68143 6239
rect 70317 6205 70351 6239
rect 71329 6205 71363 6239
rect 75193 6205 75227 6239
rect 77217 6205 77251 6239
rect 78321 6205 78355 6239
rect 80253 6205 80287 6239
rect 81081 6205 81115 6239
rect 81541 6205 81575 6239
rect 83013 6205 83047 6239
rect 83473 6205 83507 6239
rect 84117 6205 84151 6239
rect 21189 6137 21223 6171
rect 28080 6137 28114 6171
rect 31125 6137 31159 6171
rect 33241 6137 33275 6171
rect 33517 6137 33551 6171
rect 33609 6137 33643 6171
rect 38485 6137 38519 6171
rect 38761 6137 38795 6171
rect 38853 6137 38887 6171
rect 41245 6137 41279 6171
rect 41521 6137 41555 6171
rect 41613 6137 41647 6171
rect 42349 6137 42383 6171
rect 48973 6137 49007 6171
rect 18705 6069 18739 6103
rect 20545 6069 20579 6103
rect 21557 6069 21591 6103
rect 25145 6069 25179 6103
rect 34345 6069 34379 6103
rect 35357 6069 35391 6103
rect 39589 6069 39623 6103
rect 45937 6069 45971 6103
rect 49341 6069 49375 6103
rect 49801 6069 49835 6103
rect 50445 6069 50479 6103
rect 51089 6069 51123 6103
rect 54033 6069 54067 6103
rect 61669 6069 61703 6103
rect 66453 6069 66487 6103
rect 66821 6069 66855 6103
rect 67925 6069 67959 6103
rect 70133 6069 70167 6103
rect 71145 6069 71179 6103
rect 75009 6069 75043 6103
rect 77401 6069 77435 6103
rect 78505 6069 78539 6103
rect 80437 6069 80471 6103
rect 81725 6069 81759 6103
rect 82829 6069 82863 6103
rect 84301 6069 84335 6103
rect 17049 5865 17083 5899
rect 31861 5865 31895 5899
rect 34805 5865 34839 5899
rect 46213 5865 46247 5899
rect 55045 5865 55079 5899
rect 59369 5865 59403 5899
rect 63325 5865 63359 5899
rect 72433 5865 72467 5899
rect 77677 5865 77711 5899
rect 83105 5865 83139 5899
rect 15936 5797 15970 5831
rect 23112 5797 23146 5831
rect 25504 5797 25538 5831
rect 27344 5797 27378 5831
rect 42156 5797 42190 5831
rect 46121 5797 46155 5831
rect 48780 5797 48814 5831
rect 15669 5729 15703 5763
rect 17776 5729 17810 5763
rect 20904 5729 20938 5763
rect 22845 5729 22879 5763
rect 25237 5729 25271 5763
rect 27077 5729 27111 5763
rect 30481 5729 30515 5763
rect 30748 5729 30782 5763
rect 32588 5729 32622 5763
rect 34621 5729 34655 5763
rect 35909 5729 35943 5763
rect 36461 5729 36495 5763
rect 37105 5729 37139 5763
rect 39405 5729 39439 5763
rect 41429 5729 41463 5763
rect 43996 5729 44030 5763
rect 46857 5729 46891 5763
rect 47133 5729 47167 5763
rect 48053 5729 48087 5763
rect 52101 5729 52135 5763
rect 53205 5729 53239 5763
rect 53389 5729 53423 5763
rect 54263 5729 54297 5763
rect 55689 5729 55723 5763
rect 57529 5729 57563 5763
rect 58566 5729 58600 5763
rect 58725 5729 58759 5763
rect 60013 5729 60047 5763
rect 60665 5729 60699 5763
rect 64220 5729 64254 5763
rect 65901 5729 65935 5763
rect 69029 5729 69063 5763
rect 72617 5729 72651 5763
rect 73261 5729 73295 5763
rect 74089 5729 74123 5763
rect 77861 5729 77895 5763
rect 79701 5729 79735 5763
rect 80345 5729 80379 5763
rect 81725 5729 81759 5763
rect 85957 5797 85991 5831
rect 83197 5729 83231 5763
rect 84485 5729 84519 5763
rect 85129 5729 85163 5763
rect 17509 5661 17543 5695
rect 20637 5661 20671 5695
rect 32321 5661 32355 5695
rect 37381 5661 37415 5695
rect 41889 5661 41923 5695
rect 43729 5661 43763 5695
rect 47016 5661 47050 5695
rect 47869 5661 47903 5695
rect 48513 5661 48547 5695
rect 53849 5661 53883 5695
rect 54125 5661 54159 5695
rect 54399 5661 54433 5695
rect 57713 5661 57747 5695
rect 58449 5661 58483 5695
rect 64061 5661 64095 5695
rect 64337 5661 64371 5695
rect 65073 5661 65107 5695
rect 65257 5661 65291 5695
rect 83105 5661 83139 5695
rect 84025 5661 84059 5695
rect 86049 5729 86083 5763
rect 177957 5729 177991 5763
rect 28457 5593 28491 5627
rect 43269 5593 43303 5627
rect 47409 5593 47443 5627
rect 58173 5593 58207 5627
rect 64613 5593 64647 5627
rect 79517 5593 79551 5627
rect 80161 5593 80195 5627
rect 85313 5593 85347 5627
rect 85957 5593 85991 5627
rect 86233 5593 86267 5627
rect 18889 5525 18923 5559
rect 22017 5525 22051 5559
rect 24225 5525 24259 5559
rect 26617 5525 26651 5559
rect 33701 5525 33735 5559
rect 35725 5525 35759 5559
rect 36645 5525 36679 5559
rect 38669 5525 38703 5559
rect 39221 5525 39255 5559
rect 41245 5525 41279 5559
rect 45109 5525 45143 5559
rect 49893 5525 49927 5559
rect 51917 5525 51951 5559
rect 55505 5525 55539 5559
rect 59829 5525 59863 5559
rect 60473 5525 60507 5559
rect 63417 5525 63451 5559
rect 65717 5525 65751 5559
rect 68845 5525 68879 5559
rect 73077 5525 73111 5559
rect 73905 5525 73939 5559
rect 79057 5525 79091 5559
rect 81265 5525 81299 5559
rect 81909 5525 81943 5559
rect 83381 5525 83415 5559
rect 84669 5525 84703 5559
rect 34437 5321 34471 5355
rect 41521 5321 41555 5355
rect 42441 5321 42475 5355
rect 63141 5321 63175 5355
rect 69213 5321 69247 5355
rect 78229 5321 78263 5355
rect 78873 5321 78907 5355
rect 82277 5321 82311 5355
rect 18705 5253 18739 5287
rect 20545 5253 20579 5287
rect 39681 5253 39715 5287
rect 17325 5185 17359 5219
rect 19165 5185 19199 5219
rect 23857 5185 23891 5219
rect 29285 5185 29319 5219
rect 33057 5185 33091 5219
rect 34897 5185 34931 5219
rect 40141 5185 40175 5219
rect 45385 5185 45419 5219
rect 61301 5185 61335 5219
rect 61485 5185 61519 5219
rect 61945 5185 61979 5219
rect 62359 5185 62393 5219
rect 19432 5117 19466 5151
rect 33324 5117 33358 5151
rect 35164 5117 35198 5151
rect 37381 5117 37415 5151
rect 38301 5117 38335 5151
rect 42625 5117 42659 5151
rect 43545 5117 43579 5151
rect 47409 5117 47443 5151
rect 62221 5117 62255 5151
rect 62497 5117 62531 5151
rect 64705 5117 64739 5151
rect 17592 5049 17626 5083
rect 29552 5049 29586 5083
rect 38546 5049 38580 5083
rect 40408 5049 40442 5083
rect 43812 5049 43846 5083
rect 45652 5049 45686 5083
rect 82093 5253 82127 5287
rect 86969 5253 87003 5287
rect 82645 5185 82679 5219
rect 85681 5185 85715 5219
rect 75837 5117 75871 5151
rect 76665 5117 76699 5151
rect 77585 5117 77619 5151
rect 78045 5117 78079 5151
rect 78689 5117 78723 5151
rect 80437 5117 80471 5151
rect 81449 5117 81483 5151
rect 83105 5117 83139 5151
rect 83473 5117 83507 5151
rect 84117 5117 84151 5151
rect 86141 5117 86175 5151
rect 86785 5117 86819 5151
rect 87429 5117 87463 5151
rect 177313 5117 177347 5151
rect 177957 5117 177991 5151
rect 82001 5049 82035 5083
rect 82277 5049 82311 5083
rect 24869 4981 24903 5015
rect 30665 4981 30699 5015
rect 36277 4981 36311 5015
rect 37197 4981 37231 5015
rect 44925 4981 44959 5015
rect 46765 4981 46799 5015
rect 47225 4981 47259 5015
rect 64521 4981 64555 5015
rect 69213 4981 69247 5015
rect 76021 4981 76055 5015
rect 76481 4981 76515 5015
rect 81633 4981 81667 5015
rect 83289 4981 83323 5015
rect 83381 4981 83415 5015
rect 83657 4981 83691 5015
rect 84301 4981 84335 5015
rect 86325 4981 86359 5015
rect 87613 4981 87647 5015
rect 28365 4777 28399 4811
rect 33425 4777 33459 4811
rect 37013 4777 37047 4811
rect 39589 4777 39623 4811
rect 45201 4777 45235 4811
rect 79333 4777 79367 4811
rect 83933 4777 83967 4811
rect 89637 4777 89671 4811
rect 102793 4777 102827 4811
rect 36001 4709 36035 4743
rect 38476 4709 38510 4743
rect 44088 4709 44122 4743
rect 78045 4709 78079 4743
rect 80253 4709 80287 4743
rect 80989 4709 81023 4743
rect 82001 4709 82035 4743
rect 84853 4709 84887 4743
rect 85129 4709 85163 4743
rect 11805 4641 11839 4675
rect 38209 4641 38243 4675
rect 43821 4641 43855 4675
rect 46480 4641 46514 4675
rect 70593 4641 70627 4675
rect 72433 4641 72467 4675
rect 73077 4641 73111 4675
rect 74733 4641 74767 4675
rect 75561 4641 75595 4675
rect 79149 4641 79183 4675
rect 81817 4641 81851 4675
rect 83105 4641 83139 4675
rect 83197 4641 83231 4675
rect 83473 4641 83507 4675
rect 84117 4641 84151 4675
rect 84209 4641 84243 4675
rect 84485 4641 84519 4675
rect 88165 4641 88199 4675
rect 88809 4641 88843 4675
rect 89453 4641 89487 4675
rect 93777 4641 93811 4675
rect 102609 4641 102643 4675
rect 175381 4641 175415 4675
rect 176209 4641 176243 4675
rect 177313 4641 177347 4675
rect 177957 4641 177991 4675
rect 27353 4573 27387 4607
rect 32413 4573 32447 4607
rect 36645 4573 36679 4607
rect 46213 4573 46247 4607
rect 81633 4573 81667 4607
rect 83381 4573 83415 4607
rect 84393 4573 84427 4607
rect 75377 4505 75411 4539
rect 81173 4505 81207 4539
rect 84945 4505 84979 4539
rect 85497 4505 85531 4539
rect 88349 4505 88383 4539
rect 88993 4505 89027 4539
rect 93961 4505 93995 4539
rect 11989 4437 12023 4471
rect 47593 4437 47627 4471
rect 74917 4437 74951 4471
rect 76757 4437 76791 4471
rect 78137 4437 78171 4471
rect 80345 4437 80379 4471
rect 82921 4437 82955 4471
rect 85129 4437 85163 4471
rect 86141 4437 86175 4471
rect 86785 4437 86819 4471
rect 78321 4233 78355 4267
rect 81725 4233 81759 4267
rect 82921 4233 82955 4267
rect 86233 4233 86267 4267
rect 88625 4233 88659 4267
rect 88809 4233 88843 4267
rect 89453 4233 89487 4267
rect 13553 4165 13587 4199
rect 39681 4165 39715 4199
rect 51641 4165 51675 4199
rect 84577 4165 84611 4199
rect 87797 4165 87831 4199
rect 90925 4165 90959 4199
rect 94329 4165 94363 4199
rect 1409 4029 1443 4063
rect 2053 4029 2087 4063
rect 12567 4029 12601 4063
rect 36001 4097 36035 4131
rect 38301 4097 38335 4131
rect 77677 4097 77711 4131
rect 79149 4097 79183 4131
rect 83381 4097 83415 4131
rect 104725 4097 104759 4131
rect 13645 4029 13679 4063
rect 15853 4029 15887 4063
rect 20269 4029 20303 4063
rect 38568 4029 38602 4063
rect 45753 4029 45787 4063
rect 50629 4029 50663 4063
rect 51733 4029 51767 4063
rect 56977 4029 57011 4063
rect 59277 4029 59311 4063
rect 66177 4029 66211 4063
rect 67281 4029 67315 4063
rect 68385 4029 68419 4063
rect 69765 4029 69799 4063
rect 70501 4029 70535 4063
rect 71237 4029 71271 4063
rect 72065 4029 72099 4063
rect 73169 4029 73203 4063
rect 73905 4029 73939 4063
rect 75193 4029 75227 4063
rect 76021 4029 76055 4063
rect 76757 4029 76791 4063
rect 77493 4029 77527 4063
rect 80345 4029 80379 4063
rect 81357 4029 81391 4063
rect 83105 4029 83139 4063
rect 83197 4029 83231 4063
rect 83473 4029 83507 4063
rect 84209 4029 84243 4063
rect 84393 4029 84427 4063
rect 85865 4029 85899 4063
rect 86969 4029 87003 4063
rect 88257 4029 88291 4063
rect 90741 4029 90775 4063
rect 91569 4029 91603 4063
rect 92397 4029 92431 4063
rect 93041 4029 93075 4063
rect 94145 4029 94179 4063
rect 94881 4029 94915 4063
rect 95985 4029 96019 4063
rect 97089 4029 97123 4063
rect 98193 4029 98227 4063
rect 99297 4029 99331 4063
rect 101229 4029 101263 4063
rect 101873 4029 101907 4063
rect 102977 4029 103011 4063
rect 103713 4029 103747 4063
rect 13553 3961 13587 3995
rect 36268 3961 36302 3995
rect 46020 3961 46054 3995
rect 57161 3961 57195 3995
rect 78229 3961 78263 3995
rect 78965 3961 78999 3995
rect 80529 3961 80563 3995
rect 84025 3961 84059 3995
rect 88625 3961 88659 3995
rect 104817 4029 104851 4063
rect 106473 4029 106507 4063
rect 107117 4029 107151 4063
rect 111717 4029 111751 4063
rect 112545 4029 112579 4063
rect 113649 4029 113683 4063
rect 114753 4029 114787 4063
rect 115857 4029 115891 4063
rect 116961 4029 116995 4063
rect 118065 4029 118099 4063
rect 119169 4029 119203 4063
rect 120181 4029 120215 4063
rect 121101 4029 121135 4063
rect 122389 4029 122423 4063
rect 123493 4029 123527 4063
rect 124597 4029 124631 4063
rect 125701 4029 125735 4063
rect 127449 4029 127483 4063
rect 128093 4029 128127 4063
rect 131221 4029 131255 4063
rect 133429 4029 133463 4063
rect 134533 4029 134567 4063
rect 136741 4029 136775 4063
rect 137937 4029 137971 4063
rect 138949 4029 138983 4063
rect 140053 4029 140087 4063
rect 141157 4029 141191 4063
rect 142077 4029 142111 4063
rect 143365 4029 143399 4063
rect 144469 4029 144503 4063
rect 145573 4029 145607 4063
rect 146677 4029 146711 4063
rect 148425 4029 148459 4063
rect 149069 4029 149103 4063
rect 152197 4029 152231 4063
rect 153669 4029 153703 4063
rect 154405 4029 154439 4063
rect 155509 4029 155543 4063
rect 157717 4029 157751 4063
rect 158913 4029 158947 4063
rect 159925 4029 159959 4063
rect 161029 4029 161063 4063
rect 162133 4029 162167 4063
rect 165445 4029 165479 4063
rect 166549 4029 166583 4063
rect 167653 4029 167687 4063
rect 169401 4029 169435 4063
rect 170045 4029 170079 4063
rect 173173 4029 173207 4063
rect 174645 4029 174679 4063
rect 175749 4029 175783 4063
rect 176945 4029 176979 4063
rect 177405 4029 177439 4063
rect 1593 3893 1627 3927
rect 2237 3893 2271 3927
rect 37381 3893 37415 3927
rect 47133 3893 47167 3927
rect 59369 3893 59403 3927
rect 71513 3893 71547 3927
rect 75009 3893 75043 3927
rect 76205 3893 76239 3927
rect 76849 3893 76883 3927
rect 81725 3893 81759 3927
rect 81909 3893 81943 3927
rect 84301 3893 84335 3927
rect 86233 3893 86267 3927
rect 86417 3893 86451 3927
rect 87061 3893 87095 3927
rect 91753 3893 91787 3927
rect 92581 3893 92615 3927
rect 93225 3893 93259 3927
rect 95065 3893 95099 3927
rect 96169 3893 96203 3927
rect 97273 3893 97307 3927
rect 98377 3893 98411 3927
rect 99481 3893 99515 3927
rect 101413 3893 101447 3927
rect 102057 3893 102091 3927
rect 103161 3893 103195 3927
rect 103897 3893 103931 3927
rect 104725 3893 104759 3927
rect 105001 3893 105035 3927
rect 106657 3893 106691 3927
rect 107301 3893 107335 3927
rect 111901 3893 111935 3927
rect 3157 3689 3191 3723
rect 6285 3689 6319 3723
rect 10241 3689 10275 3723
rect 11161 3689 11195 3723
rect 24685 3689 24719 3723
rect 72801 3689 72835 3723
rect 75193 3689 75227 3723
rect 79425 3689 79459 3723
rect 80621 3689 80655 3723
rect 81081 3689 81115 3723
rect 81909 3689 81943 3723
rect 85037 3689 85071 3723
rect 86233 3689 86267 3723
rect 87245 3689 87279 3723
rect 88533 3689 88567 3723
rect 91017 3689 91051 3723
rect 91661 3689 91695 3723
rect 94973 3689 95007 3723
rect 104265 3689 104299 3723
rect 105369 3689 105403 3723
rect 107577 3689 107611 3723
rect 109325 3689 109359 3723
rect 109969 3689 110003 3723
rect 1685 3621 1719 3655
rect 1961 3621 1995 3655
rect 2513 3553 2547 3587
rect 3341 3553 3375 3587
rect 4997 3553 5031 3587
rect 6469 3553 6503 3587
rect 9597 3553 9631 3587
rect 1777 3417 1811 3451
rect 4813 3417 4847 3451
rect 9781 3417 9815 3451
rect 12265 3621 12299 3655
rect 13737 3621 13771 3655
rect 14841 3621 14875 3655
rect 18889 3621 18923 3655
rect 21097 3621 21131 3655
rect 10333 3553 10367 3587
rect 10977 3553 11011 3587
rect 13369 3553 13403 3587
rect 13553 3553 13587 3587
rect 14197 3553 14231 3587
rect 15485 3553 15519 3587
rect 16681 3553 16715 3587
rect 16865 3553 16899 3587
rect 17325 3553 17359 3587
rect 18061 3553 18095 3587
rect 19993 3553 20027 3587
rect 21741 3553 21775 3587
rect 22477 3553 22511 3587
rect 23581 3553 23615 3587
rect 67189 3621 67223 3655
rect 67603 3621 67637 3655
rect 68293 3621 68327 3655
rect 68707 3621 68741 3655
rect 69811 3621 69845 3655
rect 76297 3621 76331 3655
rect 80437 3621 80471 3655
rect 87061 3621 87095 3655
rect 89545 3621 89579 3655
rect 93961 3621 93995 3655
rect 25237 3553 25271 3587
rect 25881 3553 25915 3587
rect 26893 3553 26927 3587
rect 27997 3553 28031 3587
rect 31309 3553 31343 3587
rect 32413 3553 32447 3587
rect 33517 3553 33551 3587
rect 34621 3553 34655 3587
rect 35725 3553 35759 3587
rect 37933 3553 37967 3587
rect 39773 3553 39807 3587
rect 40969 3553 41003 3587
rect 41981 3553 42015 3587
rect 43085 3553 43119 3587
rect 44189 3553 44223 3587
rect 45109 3553 45143 3587
rect 46397 3553 46431 3587
rect 47501 3553 47535 3587
rect 48605 3553 48639 3587
rect 49709 3553 49743 3587
rect 54125 3553 54159 3587
rect 55229 3553 55263 3587
rect 56701 3553 56735 3587
rect 57437 3553 57471 3587
rect 58541 3553 58575 3587
rect 59645 3553 59679 3587
rect 60657 3553 60691 3587
rect 61945 3553 61979 3587
rect 62865 3553 62899 3587
rect 63969 3553 64003 3587
rect 65073 3553 65107 3587
rect 66085 3553 66119 3587
rect 67833 3553 67867 3587
rect 69406 3553 69440 3587
rect 70501 3553 70535 3587
rect 71145 3553 71179 3587
rect 73445 3553 73479 3587
rect 74365 3553 74399 3587
rect 78321 3553 78355 3587
rect 81081 3553 81115 3587
rect 81177 3553 81211 3587
rect 81357 3553 81391 3587
rect 81449 3553 81483 3587
rect 81541 3553 81575 3587
rect 81725 3553 81759 3587
rect 82921 3553 82955 3587
rect 83105 3553 83139 3587
rect 83473 3553 83507 3587
rect 84301 3553 84335 3587
rect 84485 3553 84519 3587
rect 84853 3553 84887 3587
rect 85497 3553 85531 3587
rect 85681 3553 85715 3587
rect 86049 3553 86083 3587
rect 89177 3553 89211 3587
rect 90189 3553 90223 3587
rect 90833 3553 90867 3587
rect 91477 3553 91511 3587
rect 92121 3553 92155 3587
rect 96169 3553 96203 3587
rect 96813 3553 96847 3587
rect 97457 3553 97491 3587
rect 98653 3553 98687 3587
rect 99665 3553 99699 3587
rect 100309 3553 100343 3587
rect 102701 3553 102735 3587
rect 104081 3553 104115 3587
rect 105185 3553 105219 3587
rect 106289 3553 106323 3587
rect 107393 3553 107427 3587
rect 109141 3553 109175 3587
rect 109785 3553 109819 3587
rect 110705 3553 110739 3587
rect 111809 3553 111843 3587
rect 112913 3553 112947 3587
rect 114385 3553 114419 3587
rect 115121 3553 115155 3587
rect 116225 3553 116259 3587
rect 117329 3553 117363 3587
rect 118433 3553 118467 3587
rect 119629 3553 119663 3587
rect 120549 3553 120583 3587
rect 121653 3553 121687 3587
rect 122757 3553 122791 3587
rect 123769 3553 123803 3587
rect 124965 3553 124999 3587
rect 126069 3553 126103 3587
rect 127173 3553 127207 3587
rect 128277 3553 128311 3587
rect 129013 3553 129047 3587
rect 130117 3553 130151 3587
rect 130761 3553 130795 3587
rect 132417 3553 132451 3587
rect 133061 3553 133095 3587
rect 133797 3553 133831 3587
rect 135361 3553 135395 3587
rect 136005 3553 136039 3587
rect 137109 3553 137143 3587
rect 138213 3553 138247 3587
rect 139317 3553 139351 3587
rect 140605 3553 140639 3587
rect 141525 3553 141559 3587
rect 142629 3553 142663 3587
rect 143733 3553 143767 3587
rect 144745 3553 144779 3587
rect 145941 3553 145975 3587
rect 147045 3553 147079 3587
rect 148149 3553 148183 3587
rect 149253 3553 149287 3587
rect 149989 3553 150023 3587
rect 151093 3553 151127 3587
rect 151737 3553 151771 3587
rect 153669 3553 153703 3587
rect 154773 3553 154807 3587
rect 156337 3553 156371 3587
rect 156981 3553 157015 3587
rect 158085 3553 158119 3587
rect 159189 3553 159223 3587
rect 160293 3553 160327 3587
rect 161581 3553 161615 3587
rect 162501 3553 162535 3587
rect 163605 3553 163639 3587
rect 164249 3553 164283 3587
rect 164893 3553 164927 3587
rect 165721 3553 165755 3587
rect 166917 3553 166951 3587
rect 168021 3553 168055 3587
rect 169125 3553 169159 3587
rect 170229 3553 170263 3587
rect 170965 3553 170999 3587
rect 172069 3553 172103 3587
rect 172713 3553 172747 3587
rect 174369 3553 174403 3587
rect 175013 3553 175047 3587
rect 176393 3553 176427 3587
rect 177957 3553 177991 3587
rect 72433 3485 72467 3519
rect 75929 3485 75963 3519
rect 78505 3485 78539 3519
rect 83197 3485 83231 3519
rect 83289 3485 83323 3519
rect 84577 3485 84611 3519
rect 84669 3485 84703 3519
rect 85773 3485 85807 3519
rect 85865 3485 85899 3519
rect 24685 3417 24719 3451
rect 68845 3417 68879 3451
rect 74825 3417 74859 3451
rect 79057 3417 79091 3451
rect 79609 3417 79643 3451
rect 80069 3417 80103 3451
rect 83657 3417 83691 3451
rect 86693 3417 86727 3451
rect 88165 3417 88199 3451
rect 90373 3417 90407 3451
rect 92305 3417 92339 3451
rect 96997 3417 97031 3451
rect 99849 3417 99883 3451
rect 110889 3417 110923 3451
rect 178141 3417 178175 3451
rect 2697 3349 2731 3383
rect 10241 3349 10275 3383
rect 12357 3349 12391 3383
rect 14197 3349 14231 3383
rect 14933 3349 14967 3383
rect 18981 3349 19015 3383
rect 21189 3349 21223 3383
rect 67557 3349 67591 3383
rect 68661 3349 68695 3383
rect 69765 3349 69799 3383
rect 69949 3349 69983 3383
rect 71329 3349 71363 3383
rect 72801 3349 72835 3383
rect 72985 3349 73019 3383
rect 73629 3349 73663 3383
rect 75193 3349 75227 3383
rect 75377 3349 75411 3383
rect 76297 3349 76331 3383
rect 76481 3349 76515 3383
rect 79425 3349 79459 3383
rect 80437 3349 80471 3383
rect 87061 3349 87095 3383
rect 88533 3349 88567 3383
rect 88717 3349 88751 3383
rect 89545 3349 89579 3383
rect 89729 3349 89763 3383
rect 96353 3349 96387 3383
rect 97641 3349 97675 3383
rect 98837 3349 98871 3383
rect 100493 3349 100527 3383
rect 101137 3349 101171 3383
rect 102241 3349 102275 3383
rect 102885 3349 102919 3383
rect 106473 3349 106507 3383
rect 131957 3349 131991 3383
rect 152933 3349 152967 3383
rect 173909 3349 173943 3383
rect 16313 3145 16347 3179
rect 24501 3145 24535 3179
rect 27261 3145 27295 3179
rect 66453 3145 66487 3179
rect 67557 3145 67591 3179
rect 67741 3145 67775 3179
rect 68661 3145 68695 3179
rect 70133 3145 70167 3179
rect 71237 3145 71271 3179
rect 72341 3145 72375 3179
rect 72525 3145 72559 3179
rect 75377 3145 75411 3179
rect 76389 3145 76423 3179
rect 76573 3145 76607 3179
rect 78045 3145 78079 3179
rect 78229 3145 78263 3179
rect 79057 3145 79091 3179
rect 81265 3145 81299 3179
rect 83013 3145 83047 3179
rect 84301 3145 84335 3179
rect 87889 3145 87923 3179
rect 88809 3145 88843 3179
rect 110613 3145 110647 3179
rect 9873 3077 9907 3111
rect 17693 3077 17727 3111
rect 1685 3009 1719 3043
rect 12449 3009 12483 3043
rect 15301 3009 15335 3043
rect 17325 3009 17359 3043
rect 19257 3009 19291 3043
rect 1409 2941 1443 2975
rect 2329 2941 2363 2975
rect 3065 2941 3099 2975
rect 3709 2941 3743 2975
rect 4537 2941 4571 2975
rect 5181 2941 5215 2975
rect 6837 2941 6871 2975
rect 7941 2941 7975 2975
rect 9229 2941 9263 2975
rect 9873 2941 9907 2975
rect 12081 2941 12115 2975
rect 12633 2941 12667 2975
rect 14013 2941 14047 2975
rect 14289 2941 14323 2975
rect 15485 2941 15519 2975
rect 17509 2941 17543 2975
rect 18245 2941 18279 2975
rect 18889 2941 18923 2975
rect 19073 2941 19107 2975
rect 20177 2941 20211 2975
rect 20637 2941 20671 2975
rect 20913 2941 20947 2975
rect 22661 2941 22695 2975
rect 23397 2941 23431 2975
rect 24409 2941 24443 2975
rect 70317 3077 70351 3111
rect 76021 3077 76055 3111
rect 78689 3077 78723 3111
rect 80713 3077 80747 3111
rect 81725 3077 81759 3111
rect 86969 3077 87003 3111
rect 90925 3077 90959 3111
rect 68293 3009 68327 3043
rect 75009 3009 75043 3043
rect 85773 3009 85807 3043
rect 86518 3009 86552 3043
rect 91569 3009 91603 3043
rect 96813 3009 96847 3043
rect 101321 3009 101355 3043
rect 107761 3009 107795 3043
rect 109969 3009 110003 3043
rect 29469 2941 29503 2975
rect 30205 2941 30239 2975
rect 31033 2941 31067 2975
rect 31953 2941 31987 2975
rect 33241 2941 33275 2975
rect 34345 2941 34379 2975
rect 35449 2941 35483 2975
rect 37197 2941 37231 2975
rect 39773 2941 39807 2975
rect 40417 2941 40451 2975
rect 41245 2941 41279 2975
rect 42349 2941 42383 2975
rect 43545 2941 43579 2975
rect 44557 2941 44591 2975
rect 45661 2941 45695 2975
rect 46765 2941 46799 2975
rect 47685 2941 47719 2975
rect 48973 2941 49007 2975
rect 50077 2941 50111 2975
rect 50813 2941 50847 2975
rect 51641 2941 51675 2975
rect 52285 2941 52319 2975
rect 52929 2941 52963 2975
rect 54033 2941 54067 2975
rect 54677 2941 54711 2975
rect 55597 2941 55631 2975
rect 56701 2941 56735 2975
rect 57805 2941 57839 2975
rect 59277 2941 59311 2975
rect 60013 2941 60047 2975
rect 61025 2941 61059 2975
rect 62129 2941 62163 2975
rect 63233 2941 63267 2975
rect 64521 2941 64555 2975
rect 65441 2941 65475 2975
rect 66729 2941 66763 2975
rect 67189 2941 67223 2975
rect 69765 2941 69799 2975
rect 70869 2941 70903 2975
rect 71513 2941 71547 2975
rect 71973 2941 72007 2975
rect 73629 2941 73663 2975
rect 77217 2941 77251 2975
rect 77677 2941 77711 2975
rect 80253 2941 80287 2975
rect 80437 2941 80471 2975
rect 80529 2941 80563 2975
rect 80805 2941 80839 2975
rect 81449 2941 81483 2975
rect 81541 2941 81575 2975
rect 81817 2941 81851 2975
rect 82277 2941 82311 2975
rect 82461 2941 82495 2975
rect 82553 2941 82587 2975
rect 82645 2941 82679 2975
rect 82829 2941 82863 2975
rect 83565 2941 83599 2975
rect 83749 2941 83783 2975
rect 83841 2941 83875 2975
rect 83933 2941 83967 2975
rect 84117 2941 84151 2975
rect 86233 2941 86267 2975
rect 86405 2941 86439 2975
rect 86601 2941 86635 2975
rect 86785 2941 86819 2975
rect 87613 2941 87647 2975
rect 87705 2941 87739 2975
rect 87963 2941 87997 2975
rect 88441 2941 88475 2975
rect 89545 2941 89579 2975
rect 92305 2941 92339 2975
rect 93409 2941 93443 2975
rect 94513 2941 94547 2975
rect 96169 2941 96203 2975
rect 97825 2941 97859 2975
rect 98929 2941 98963 2975
rect 100033 2941 100067 2975
rect 103713 2941 103747 2975
rect 104449 2941 104483 2975
rect 105553 2941 105587 2975
rect 106657 2941 106691 2975
rect 108865 2941 108899 2975
rect 110429 2941 110463 2975
rect 111901 2941 111935 2975
rect 112545 2941 112579 2975
rect 113281 2941 113315 2975
rect 114385 2941 114419 2975
rect 115489 2941 115523 2975
rect 117145 2941 117179 2975
rect 117789 2941 117823 2975
rect 118801 2941 118835 2975
rect 119905 2941 119939 2975
rect 120917 2941 120951 2975
rect 122389 2941 122423 2975
rect 123125 2941 123159 2975
rect 124229 2941 124263 2975
rect 125333 2941 125367 2975
rect 126437 2941 126471 2975
rect 127633 2941 127667 2975
rect 128645 2941 128679 2975
rect 129749 2941 129783 2975
rect 130853 2941 130887 2975
rect 131313 2941 131347 2975
rect 133061 2941 133095 2975
rect 134165 2941 134199 2975
rect 135269 2941 135303 2975
rect 136373 2941 136407 2975
rect 136833 2941 136867 2975
rect 138121 2941 138155 2975
rect 138765 2941 138799 2975
rect 139685 2941 139719 2975
rect 140789 2941 140823 2975
rect 141893 2941 141927 2975
rect 143365 2941 143399 2975
rect 144101 2941 144135 2975
rect 145205 2941 145239 2975
rect 146309 2941 146343 2975
rect 147413 2941 147447 2975
rect 148609 2941 148643 2975
rect 149621 2941 149655 2975
rect 150725 2941 150759 2975
rect 151829 2941 151863 2975
rect 152565 2941 152599 2975
rect 154037 2941 154071 2975
rect 155141 2941 155175 2975
rect 156245 2941 156279 2975
rect 157349 2941 157383 2975
rect 157809 2941 157843 2975
rect 159097 2941 159131 2975
rect 159741 2941 159775 2975
rect 160661 2941 160695 2975
rect 161765 2941 161799 2975
rect 162869 2941 162903 2975
rect 164341 2941 164375 2975
rect 165077 2941 165111 2975
rect 166181 2941 166215 2975
rect 167285 2941 167319 2975
rect 168389 2941 168423 2975
rect 169585 2941 169619 2975
rect 170597 2941 170631 2975
rect 171701 2941 171735 2975
rect 172805 2941 172839 2975
rect 173265 2941 173299 2975
rect 175013 2941 175047 2975
rect 176117 2941 176151 2975
rect 176945 2941 176979 2975
rect 177957 2941 177991 2975
rect 10057 2873 10091 2907
rect 10977 2873 11011 2907
rect 13369 2873 13403 2907
rect 16221 2873 16255 2907
rect 18429 2873 18463 2907
rect 19993 2873 20027 2907
rect 25513 2873 25547 2907
rect 26617 2873 26651 2907
rect 27261 2873 27295 2907
rect 27905 2873 27939 2907
rect 28825 2873 28859 2907
rect 36553 2873 36587 2907
rect 38393 2873 38427 2907
rect 39129 2873 39163 2907
rect 66085 2873 66119 2907
rect 66499 2873 66533 2907
rect 67603 2873 67637 2907
rect 68661 2873 68695 2907
rect 70179 2873 70213 2907
rect 71283 2873 71317 2907
rect 75377 2873 75411 2907
rect 76389 2873 76423 2907
rect 78045 2873 78079 2907
rect 79057 2873 79091 2907
rect 85589 2873 85623 2907
rect 87429 2873 87463 2907
rect 178141 2873 178175 2907
rect 3157 2805 3191 2839
rect 4629 2805 4663 2839
rect 7757 2805 7791 2839
rect 10149 2805 10183 2839
rect 11069 2805 11103 2839
rect 13461 2805 13495 2839
rect 15669 2805 15703 2839
rect 22753 2805 22787 2839
rect 23489 2805 23523 2839
rect 25605 2805 25639 2839
rect 26709 2805 26743 2839
rect 27997 2805 28031 2839
rect 28917 2805 28951 2839
rect 31125 2805 31159 2839
rect 32045 2805 32079 2839
rect 33333 2805 33367 2839
rect 34437 2805 34471 2839
rect 35541 2805 35575 2839
rect 36645 2805 36679 2839
rect 38485 2805 38519 2839
rect 39221 2805 39255 2839
rect 68845 2805 68879 2839
rect 72341 2805 72375 2839
rect 73721 2805 73755 2839
rect 75561 2805 75595 2839
rect 79241 2805 79275 2839
rect 88809 2805 88843 2839
rect 88993 2805 89027 2839
rect 89637 2805 89671 2839
rect 102333 2805 102367 2839
rect 10517 2601 10551 2635
rect 37381 2601 37415 2635
rect 74549 2601 74583 2635
rect 82921 2601 82955 2635
rect 84301 2601 84335 2635
rect 85313 2601 85347 2635
rect 89821 2601 89855 2635
rect 95893 2601 95927 2635
rect 111165 2601 111199 2635
rect 5825 2533 5859 2567
rect 11161 2533 11195 2567
rect 31953 2533 31987 2567
rect 39773 2533 39807 2567
rect 40509 2533 40543 2567
rect 45109 2533 45143 2567
rect 45845 2533 45879 2567
rect 47225 2533 47259 2567
rect 50537 2533 50571 2567
rect 52377 2533 52411 2567
rect 53849 2533 53883 2567
rect 55045 2533 55079 2567
rect 61485 2533 61519 2567
rect 63049 2533 63083 2567
rect 63785 2533 63819 2567
rect 67005 2533 67039 2567
rect 68385 2533 68419 2567
rect 69213 2533 69247 2567
rect 71881 2533 71915 2567
rect 73721 2533 73755 2567
rect 74457 2533 74491 2567
rect 75193 2533 75227 2567
rect 76573 2533 76607 2567
rect 76849 2533 76883 2567
rect 79057 2533 79091 2567
rect 80069 2533 80103 2567
rect 80345 2533 80379 2567
rect 86877 2533 86911 2567
rect 87153 2533 87187 2567
rect 87889 2533 87923 2567
rect 88165 2533 88199 2567
rect 90465 2533 90499 2567
rect 92397 2533 92431 2567
rect 93133 2533 93167 2567
rect 93869 2533 93903 2567
rect 95801 2533 95835 2567
rect 96537 2533 96571 2567
rect 97733 2533 97767 2567
rect 98469 2533 98503 2567
rect 99205 2533 99239 2567
rect 100401 2533 100435 2567
rect 101137 2533 101171 2567
rect 101873 2533 101907 2567
rect 103069 2533 103103 2567
rect 103805 2533 103839 2567
rect 104541 2533 104575 2567
rect 105737 2533 105771 2567
rect 106749 2533 106783 2567
rect 109141 2533 109175 2567
rect 109877 2533 109911 2567
rect 111809 2533 111843 2567
rect 112545 2533 112579 2567
rect 113741 2533 113775 2567
rect 114477 2533 114511 2567
rect 115213 2533 115247 2567
rect 116409 2533 116443 2567
rect 117145 2533 117179 2567
rect 117881 2533 117915 2567
rect 119077 2533 119111 2567
rect 119997 2533 120031 2567
rect 121745 2533 121779 2567
rect 122481 2533 122515 2567
rect 123217 2533 123251 2567
rect 124413 2533 124447 2567
rect 125425 2533 125459 2567
rect 127081 2533 127115 2567
rect 127817 2533 127851 2567
rect 128553 2533 128587 2567
rect 129841 2533 129875 2567
rect 130945 2533 130979 2567
rect 132417 2533 132451 2567
rect 133153 2533 133187 2567
rect 135085 2533 135119 2567
rect 135821 2533 135855 2567
rect 136557 2533 136591 2567
rect 137753 2533 137787 2567
rect 138673 2533 138707 2567
rect 140421 2533 140455 2567
rect 141157 2533 141191 2567
rect 141893 2533 141927 2567
rect 143089 2533 143123 2567
rect 144193 2533 144227 2567
rect 145757 2533 145791 2567
rect 146493 2533 146527 2567
rect 147229 2533 147263 2567
rect 148609 2533 148643 2567
rect 149713 2533 149747 2567
rect 151093 2533 151127 2567
rect 151921 2533 151955 2567
rect 153761 2533 153795 2567
rect 154497 2533 154531 2567
rect 155233 2533 155267 2567
rect 156429 2533 156463 2567
rect 157441 2533 157475 2567
rect 159097 2533 159131 2567
rect 159833 2533 159867 2567
rect 160569 2533 160603 2567
rect 161857 2533 161891 2567
rect 162961 2533 162995 2567
rect 164433 2533 164467 2567
rect 165169 2533 165203 2567
rect 167101 2533 167135 2567
rect 167837 2533 167871 2567
rect 168573 2533 168607 2567
rect 169769 2533 169803 2567
rect 170689 2533 170723 2567
rect 172437 2533 172471 2567
rect 173173 2533 173207 2567
rect 173909 2533 173943 2567
rect 175105 2533 175139 2567
rect 176209 2533 176243 2567
rect 177773 2533 177807 2567
rect 1409 2465 1443 2499
rect 1685 2465 1719 2499
rect 2697 2465 2731 2499
rect 4353 2465 4387 2499
rect 5641 2465 5675 2499
rect 7113 2465 7147 2499
rect 7757 2465 7791 2499
rect 8493 2465 8527 2499
rect 9689 2465 9723 2499
rect 10425 2465 10459 2499
rect 12265 2465 12299 2499
rect 13185 2465 13219 2499
rect 15209 2465 15243 2499
rect 16313 2465 16347 2499
rect 17693 2465 17727 2499
rect 18705 2465 18739 2499
rect 21833 2465 21867 2499
rect 23029 2465 23063 2499
rect 24041 2465 24075 2499
rect 25697 2465 25731 2499
rect 26433 2465 26467 2499
rect 27169 2465 27203 2499
rect 28457 2465 28491 2499
rect 29561 2465 29595 2499
rect 31033 2465 31067 2499
rect 31769 2465 31803 2499
rect 32505 2465 32539 2499
rect 33701 2465 33735 2499
rect 34437 2465 34471 2499
rect 35173 2465 35207 2499
rect 36369 2465 36403 2499
rect 37289 2465 37323 2499
rect 39037 2465 39071 2499
rect 41705 2465 41739 2499
rect 42809 2465 42843 2499
rect 44373 2465 44407 2499
rect 48329 2465 48363 2499
rect 49709 2465 49743 2499
rect 51181 2465 51215 2499
rect 53113 2465 53147 2499
rect 56057 2465 56091 2499
rect 57713 2465 57747 2499
rect 58449 2465 58483 2499
rect 59185 2465 59219 2499
rect 60381 2465 60415 2499
rect 64521 2465 64555 2499
rect 65901 2465 65935 2499
rect 69857 2465 69891 2499
rect 72525 2465 72559 2499
rect 77769 2465 77803 2499
rect 82185 2465 82219 2499
rect 82369 2465 82403 2499
rect 82553 2465 82587 2499
rect 82737 2465 82771 2499
rect 84485 2465 84519 2499
rect 84577 2465 84611 2499
rect 84853 2465 84887 2499
rect 85497 2465 85531 2499
rect 85589 2465 85623 2499
rect 85865 2465 85899 2499
rect 88533 2465 88567 2499
rect 89729 2465 89763 2499
rect 91201 2465 91235 2499
rect 95065 2465 95099 2499
rect 108405 2465 108439 2499
rect 111073 2465 111107 2499
rect 133797 2465 133831 2499
rect 152565 2465 152599 2499
rect 165813 2465 165847 2499
rect 9873 2397 9907 2431
rect 12909 2397 12943 2431
rect 18429 2397 18463 2431
rect 20269 2397 20303 2431
rect 20545 2397 20579 2431
rect 77217 2397 77251 2431
rect 82461 2397 82495 2431
rect 87521 2397 87555 2431
rect 92581 2397 92615 2431
rect 95249 2397 95283 2431
rect 97917 2397 97951 2431
rect 99389 2397 99423 2431
rect 101321 2397 101355 2431
rect 109325 2397 109359 2431
rect 111993 2397 112027 2431
rect 4537 2329 4571 2363
rect 26617 2329 26651 2363
rect 27353 2329 27387 2363
rect 28641 2329 28675 2363
rect 29745 2329 29779 2363
rect 32689 2329 32723 2363
rect 33885 2329 33919 2363
rect 35357 2329 35391 2363
rect 59369 2329 59403 2363
rect 64705 2329 64739 2363
rect 71513 2329 71547 2363
rect 73905 2329 73939 2363
rect 75377 2329 75411 2363
rect 79241 2329 79275 2363
rect 80713 2329 80747 2363
rect 90649 2329 90683 2363
rect 94053 2329 94087 2363
rect 98653 2329 98687 2363
rect 100585 2329 100619 2363
rect 102057 2329 102091 2363
rect 110061 2329 110095 2363
rect 113925 2329 113959 2363
rect 115397 2329 115431 2363
rect 117329 2329 117363 2363
rect 125609 2329 125643 2363
rect 131129 2329 131163 2363
rect 147413 2329 147447 2363
rect 175289 2329 175323 2363
rect 2789 2261 2823 2295
rect 7205 2261 7239 2295
rect 8585 2261 8619 2295
rect 11253 2261 11287 2295
rect 15301 2261 15335 2295
rect 16405 2261 16439 2295
rect 17785 2261 17819 2295
rect 21925 2261 21959 2295
rect 23121 2261 23155 2295
rect 24133 2261 24167 2295
rect 25789 2261 25823 2295
rect 31125 2261 31159 2295
rect 34529 2261 34563 2295
rect 36461 2261 36495 2295
rect 39129 2261 39163 2295
rect 39865 2261 39899 2295
rect 40601 2261 40635 2295
rect 41797 2261 41831 2295
rect 42901 2261 42935 2295
rect 44465 2261 44499 2295
rect 45201 2261 45235 2295
rect 45937 2261 45971 2295
rect 47317 2261 47351 2295
rect 48421 2261 48455 2295
rect 49801 2261 49835 2295
rect 50629 2261 50663 2295
rect 52469 2261 52503 2295
rect 53205 2261 53239 2295
rect 53941 2261 53975 2295
rect 55137 2261 55171 2295
rect 56149 2261 56183 2295
rect 57805 2261 57839 2295
rect 58541 2261 58575 2295
rect 60473 2261 60507 2295
rect 61577 2261 61611 2295
rect 63141 2261 63175 2295
rect 63877 2261 63911 2295
rect 65993 2261 66027 2295
rect 67097 2261 67131 2295
rect 68477 2261 68511 2295
rect 69305 2261 69339 2295
rect 71881 2261 71915 2295
rect 72065 2261 72099 2295
rect 76665 2261 76699 2295
rect 76849 2261 76883 2295
rect 77861 2261 77895 2295
rect 80161 2261 80195 2295
rect 80345 2261 80379 2295
rect 84761 2261 84795 2295
rect 85773 2261 85807 2295
rect 86969 2261 87003 2295
rect 87153 2261 87187 2295
rect 87981 2261 88015 2295
rect 88165 2261 88199 2295
rect 91293 2261 91327 2295
rect 93225 2261 93259 2295
rect 96629 2261 96663 2295
rect 103161 2261 103195 2295
rect 103897 2261 103931 2295
rect 104633 2261 104667 2295
rect 105829 2261 105863 2295
rect 106841 2261 106875 2295
rect 108497 2261 108531 2295
rect 112637 2261 112671 2295
rect 114569 2261 114603 2295
rect 116501 2261 116535 2295
rect 117973 2261 118007 2295
rect 119169 2261 119203 2295
rect 120089 2261 120123 2295
rect 121837 2261 121871 2295
rect 122573 2261 122607 2295
rect 123309 2261 123343 2295
rect 124505 2261 124539 2295
rect 127173 2261 127207 2295
rect 127909 2261 127943 2295
rect 128645 2261 128679 2295
rect 129933 2261 129967 2295
rect 132509 2261 132543 2295
rect 133245 2261 133279 2295
rect 135177 2261 135211 2295
rect 135913 2261 135947 2295
rect 136649 2261 136683 2295
rect 137845 2261 137879 2295
rect 138765 2261 138799 2295
rect 140513 2261 140547 2295
rect 141249 2261 141283 2295
rect 141985 2261 142019 2295
rect 143181 2261 143215 2295
rect 144285 2261 144319 2295
rect 145849 2261 145883 2295
rect 146585 2261 146619 2295
rect 148701 2261 148735 2295
rect 149805 2261 149839 2295
rect 151185 2261 151219 2295
rect 152013 2261 152047 2295
rect 153853 2261 153887 2295
rect 154589 2261 154623 2295
rect 155325 2261 155359 2295
rect 156521 2261 156555 2295
rect 157533 2261 157567 2295
rect 159189 2261 159223 2295
rect 159925 2261 159959 2295
rect 160661 2261 160695 2295
rect 161949 2261 161983 2295
rect 163053 2261 163087 2295
rect 164525 2261 164559 2295
rect 165261 2261 165295 2295
rect 167193 2261 167227 2295
rect 167929 2261 167963 2295
rect 168665 2261 168699 2295
rect 169861 2261 169895 2295
rect 170781 2261 170815 2295
rect 172529 2261 172563 2295
rect 173265 2261 173299 2295
rect 174001 2261 174035 2295
rect 176301 2261 176335 2295
rect 177865 2261 177899 2295
rect 61209 2057 61243 2091
rect 48605 1989 48639 2023
rect 61209 1649 61243 1683
rect 77125 2057 77159 2091
rect 48605 1581 48639 1615
rect 90281 2057 90315 2091
rect 88625 1853 88659 1887
rect 87061 1649 87095 1683
rect 87061 1513 87095 1547
rect 88625 1513 88659 1547
rect 90189 1717 90223 1751
rect 90281 1717 90315 1751
rect 90189 1513 90223 1547
rect 77125 1445 77159 1479
<< metal1 >>
rect 1104 117530 178848 117552
rect 1104 117478 4246 117530
rect 4298 117478 4310 117530
rect 4362 117478 4374 117530
rect 4426 117478 4438 117530
rect 4490 117478 34966 117530
rect 35018 117478 35030 117530
rect 35082 117478 35094 117530
rect 35146 117478 35158 117530
rect 35210 117478 65686 117530
rect 65738 117478 65750 117530
rect 65802 117478 65814 117530
rect 65866 117478 65878 117530
rect 65930 117478 96406 117530
rect 96458 117478 96470 117530
rect 96522 117478 96534 117530
rect 96586 117478 96598 117530
rect 96650 117478 127126 117530
rect 127178 117478 127190 117530
rect 127242 117478 127254 117530
rect 127306 117478 127318 117530
rect 127370 117478 157846 117530
rect 157898 117478 157910 117530
rect 157962 117478 157974 117530
rect 158026 117478 158038 117530
rect 158090 117478 178848 117530
rect 1104 117456 178848 117478
rect 2314 117240 2320 117292
rect 2372 117280 2378 117292
rect 2593 117283 2651 117289
rect 2593 117280 2605 117283
rect 2372 117252 2605 117280
rect 2372 117240 2378 117252
rect 2593 117249 2605 117252
rect 2639 117249 2651 117283
rect 2593 117243 2651 117249
rect 3878 117240 3884 117292
rect 3936 117280 3942 117292
rect 4525 117283 4583 117289
rect 4525 117280 4537 117283
rect 3936 117252 4537 117280
rect 3936 117240 3942 117252
rect 4525 117249 4537 117252
rect 4571 117249 4583 117283
rect 4525 117243 4583 117249
rect 7006 117240 7012 117292
rect 7064 117280 7070 117292
rect 7285 117283 7343 117289
rect 7285 117280 7297 117283
rect 7064 117252 7297 117280
rect 7064 117240 7070 117252
rect 7285 117249 7297 117252
rect 7331 117249 7343 117283
rect 7285 117243 7343 117249
rect 8570 117240 8576 117292
rect 8628 117280 8634 117292
rect 8665 117283 8723 117289
rect 8665 117280 8677 117283
rect 8628 117252 8677 117280
rect 8628 117240 8634 117252
rect 8665 117249 8677 117252
rect 8711 117249 8723 117283
rect 8665 117243 8723 117249
rect 11698 117240 11704 117292
rect 11756 117280 11762 117292
rect 12529 117283 12587 117289
rect 12529 117280 12541 117283
rect 11756 117252 12541 117280
rect 11756 117240 11762 117252
rect 12529 117249 12541 117252
rect 12575 117249 12587 117283
rect 12529 117243 12587 117249
rect 13262 117240 13268 117292
rect 13320 117280 13326 117292
rect 13541 117283 13599 117289
rect 13541 117280 13553 117283
rect 13320 117252 13553 117280
rect 13320 117240 13326 117252
rect 13541 117249 13553 117252
rect 13587 117249 13599 117283
rect 13541 117243 13599 117249
rect 16574 117240 16580 117292
rect 16632 117280 16638 117292
rect 16669 117283 16727 117289
rect 16669 117280 16681 117283
rect 16632 117252 16681 117280
rect 16632 117240 16638 117252
rect 16669 117249 16681 117252
rect 16715 117249 16727 117283
rect 16669 117243 16727 117249
rect 17954 117240 17960 117292
rect 18012 117280 18018 117292
rect 18233 117283 18291 117289
rect 18233 117280 18245 117283
rect 18012 117252 18245 117280
rect 18012 117240 18018 117252
rect 18233 117249 18245 117252
rect 18279 117249 18291 117283
rect 18233 117243 18291 117249
rect 21082 117240 21088 117292
rect 21140 117280 21146 117292
rect 21361 117283 21419 117289
rect 21361 117280 21373 117283
rect 21140 117252 21373 117280
rect 21140 117240 21146 117252
rect 21361 117249 21373 117252
rect 21407 117249 21419 117283
rect 21361 117243 21419 117249
rect 22646 117240 22652 117292
rect 22704 117280 22710 117292
rect 23201 117283 23259 117289
rect 23201 117280 23213 117283
rect 22704 117252 23213 117280
rect 22704 117240 22710 117252
rect 23201 117249 23213 117252
rect 23247 117249 23259 117283
rect 23201 117243 23259 117249
rect 25774 117240 25780 117292
rect 25832 117280 25838 117292
rect 26053 117283 26111 117289
rect 26053 117280 26065 117283
rect 25832 117252 26065 117280
rect 25832 117240 25838 117252
rect 26053 117249 26065 117252
rect 26099 117249 26111 117283
rect 27338 117280 27344 117292
rect 27299 117252 27344 117280
rect 26053 117243 26111 117249
rect 27338 117240 27344 117252
rect 27396 117240 27402 117292
rect 30466 117240 30472 117292
rect 30524 117280 30530 117292
rect 31205 117283 31263 117289
rect 31205 117280 31217 117283
rect 30524 117252 31217 117280
rect 30524 117240 30530 117252
rect 31205 117249 31217 117252
rect 31251 117249 31263 117283
rect 31205 117243 31263 117249
rect 32030 117240 32036 117292
rect 32088 117280 32094 117292
rect 32309 117283 32367 117289
rect 32309 117280 32321 117283
rect 32088 117252 32321 117280
rect 32088 117240 32094 117252
rect 32309 117249 32321 117252
rect 32355 117249 32367 117283
rect 35342 117280 35348 117292
rect 35303 117252 35348 117280
rect 32309 117243 32367 117249
rect 35342 117240 35348 117252
rect 35400 117240 35406 117292
rect 36722 117240 36728 117292
rect 36780 117280 36786 117292
rect 37001 117283 37059 117289
rect 37001 117280 37013 117283
rect 36780 117252 37013 117280
rect 36780 117240 36786 117252
rect 37001 117249 37013 117252
rect 37047 117249 37059 117283
rect 37001 117243 37059 117249
rect 40034 117240 40040 117292
rect 40092 117280 40098 117292
rect 40129 117283 40187 117289
rect 40129 117280 40141 117283
rect 40092 117252 40141 117280
rect 40092 117240 40098 117252
rect 40129 117249 40141 117252
rect 40175 117249 40187 117283
rect 40129 117243 40187 117249
rect 41414 117240 41420 117292
rect 41472 117280 41478 117292
rect 41877 117283 41935 117289
rect 41877 117280 41889 117283
rect 41472 117252 41889 117280
rect 41472 117240 41478 117252
rect 41877 117249 41889 117252
rect 41923 117249 41935 117283
rect 41877 117243 41935 117249
rect 44542 117240 44548 117292
rect 44600 117280 44606 117292
rect 44821 117283 44879 117289
rect 44821 117280 44833 117283
rect 44600 117252 44833 117280
rect 44600 117240 44606 117252
rect 44821 117249 44833 117252
rect 44867 117249 44879 117283
rect 44821 117243 44879 117249
rect 46106 117240 46112 117292
rect 46164 117280 46170 117292
rect 47213 117283 47271 117289
rect 47213 117280 47225 117283
rect 46164 117252 47225 117280
rect 46164 117240 46170 117252
rect 47213 117249 47225 117252
rect 47259 117249 47271 117283
rect 47213 117243 47271 117249
rect 49234 117240 49240 117292
rect 49292 117280 49298 117292
rect 49881 117283 49939 117289
rect 49881 117280 49893 117283
rect 49292 117252 49893 117280
rect 49292 117240 49298 117252
rect 49881 117249 49893 117252
rect 49927 117249 49939 117283
rect 51074 117280 51080 117292
rect 51035 117252 51080 117280
rect 49881 117243 49939 117249
rect 51074 117240 51080 117252
rect 51132 117240 51138 117292
rect 53926 117240 53932 117292
rect 53984 117280 53990 117292
rect 54021 117283 54079 117289
rect 54021 117280 54033 117283
rect 53984 117252 54033 117280
rect 53984 117240 53990 117252
rect 54021 117249 54033 117252
rect 54067 117249 54079 117283
rect 54021 117243 54079 117249
rect 55490 117240 55496 117292
rect 55548 117280 55554 117292
rect 55769 117283 55827 117289
rect 55769 117280 55781 117283
rect 55548 117252 55781 117280
rect 55548 117240 55554 117252
rect 55769 117249 55781 117252
rect 55815 117249 55827 117283
rect 55769 117243 55827 117249
rect 58618 117240 58624 117292
rect 58676 117280 58682 117292
rect 58897 117283 58955 117289
rect 58897 117280 58909 117283
rect 58676 117252 58909 117280
rect 58676 117240 58682 117252
rect 58897 117249 58909 117252
rect 58943 117249 58955 117283
rect 58897 117243 58955 117249
rect 60182 117240 60188 117292
rect 60240 117280 60246 117292
rect 60553 117283 60611 117289
rect 60553 117280 60565 117283
rect 60240 117252 60565 117280
rect 60240 117240 60246 117252
rect 60553 117249 60565 117252
rect 60599 117249 60611 117283
rect 60553 117243 60611 117249
rect 63494 117240 63500 117292
rect 63552 117280 63558 117292
rect 63589 117283 63647 117289
rect 63589 117280 63601 117283
rect 63552 117252 63601 117280
rect 63552 117240 63558 117252
rect 63589 117249 63601 117252
rect 63635 117249 63647 117283
rect 63589 117243 63647 117249
rect 64874 117240 64880 117292
rect 64932 117280 64938 117292
rect 65889 117283 65947 117289
rect 65889 117280 65901 117283
rect 64932 117252 65901 117280
rect 64932 117240 64938 117252
rect 65889 117249 65901 117252
rect 65935 117249 65947 117283
rect 65889 117243 65947 117249
rect 68002 117240 68008 117292
rect 68060 117280 68066 117292
rect 68557 117283 68615 117289
rect 68557 117280 68569 117283
rect 68060 117252 68569 117280
rect 68060 117240 68066 117252
rect 68557 117249 68569 117252
rect 68603 117249 68615 117283
rect 68557 117243 68615 117249
rect 69566 117240 69572 117292
rect 69624 117280 69630 117292
rect 69845 117283 69903 117289
rect 69845 117280 69857 117283
rect 69624 117252 69857 117280
rect 69624 117240 69630 117252
rect 69845 117249 69857 117252
rect 69891 117249 69903 117283
rect 72694 117280 72700 117292
rect 72655 117252 72700 117280
rect 69845 117243 69903 117249
rect 72694 117240 72700 117252
rect 72752 117240 72758 117292
rect 74258 117240 74264 117292
rect 74316 117280 74322 117292
rect 74537 117283 74595 117289
rect 74537 117280 74549 117283
rect 74316 117252 74549 117280
rect 74316 117240 74322 117252
rect 74537 117249 74549 117252
rect 74583 117249 74595 117283
rect 74537 117243 74595 117249
rect 77386 117240 77392 117292
rect 77444 117280 77450 117292
rect 77665 117283 77723 117289
rect 77665 117280 77677 117283
rect 77444 117252 77677 117280
rect 77444 117240 77450 117252
rect 77665 117249 77677 117252
rect 77711 117249 77723 117283
rect 77665 117243 77723 117249
rect 78950 117240 78956 117292
rect 79008 117280 79014 117292
rect 79229 117283 79287 117289
rect 79229 117280 79241 117283
rect 79008 117252 79241 117280
rect 79008 117240 79014 117252
rect 79229 117249 79241 117252
rect 79275 117249 79287 117283
rect 79229 117243 79287 117249
rect 79336 117252 80652 117280
rect 750 117172 756 117224
rect 808 117212 814 117224
rect 1397 117215 1455 117221
rect 1397 117212 1409 117215
rect 808 117184 1409 117212
rect 808 117172 814 117184
rect 1397 117181 1409 117184
rect 1443 117181 1455 117215
rect 5442 117212 5448 117224
rect 5403 117184 5448 117212
rect 1397 117175 1455 117181
rect 5442 117172 5448 117184
rect 5500 117172 5506 117224
rect 10134 117212 10140 117224
rect 10095 117184 10140 117212
rect 10134 117172 10140 117184
rect 10192 117172 10198 117224
rect 14826 117172 14832 117224
rect 14884 117212 14890 117224
rect 14921 117215 14979 117221
rect 14921 117212 14933 117215
rect 14884 117184 14933 117212
rect 14884 117172 14890 117184
rect 14921 117181 14933 117184
rect 14967 117181 14979 117215
rect 14921 117175 14979 117181
rect 19518 117172 19524 117224
rect 19576 117212 19582 117224
rect 20257 117215 20315 117221
rect 20257 117212 20269 117215
rect 19576 117184 20269 117212
rect 19576 117172 19582 117184
rect 20257 117181 20269 117184
rect 20303 117181 20315 117215
rect 24210 117212 24216 117224
rect 24171 117184 24216 117212
rect 20257 117175 20315 117181
rect 24210 117172 24216 117184
rect 24268 117172 24274 117224
rect 28902 117212 28908 117224
rect 28863 117184 28908 117212
rect 28902 117172 28908 117184
rect 28960 117172 28966 117224
rect 33594 117212 33600 117224
rect 33555 117184 33600 117212
rect 33594 117172 33600 117184
rect 33652 117172 33658 117224
rect 35161 117215 35219 117221
rect 35161 117181 35173 117215
rect 35207 117212 35219 117215
rect 35250 117212 35256 117224
rect 35207 117184 35256 117212
rect 35207 117181 35219 117184
rect 35161 117175 35219 117181
rect 35250 117172 35256 117184
rect 35308 117172 35314 117224
rect 38286 117172 38292 117224
rect 38344 117212 38350 117224
rect 38933 117215 38991 117221
rect 38933 117212 38945 117215
rect 38344 117184 38945 117212
rect 38344 117172 38350 117184
rect 38933 117181 38945 117184
rect 38979 117181 38991 117215
rect 42978 117212 42984 117224
rect 42939 117184 42984 117212
rect 38933 117175 38991 117181
rect 42978 117172 42984 117184
rect 43036 117172 43042 117224
rect 47670 117212 47676 117224
rect 47631 117184 47676 117212
rect 47670 117172 47676 117184
rect 47728 117172 47734 117224
rect 52362 117212 52368 117224
rect 52323 117184 52368 117212
rect 52362 117172 52368 117184
rect 52420 117172 52426 117224
rect 57054 117172 57060 117224
rect 57112 117212 57118 117224
rect 57609 117215 57667 117221
rect 57609 117212 57621 117215
rect 57112 117184 57621 117212
rect 57112 117172 57118 117184
rect 57609 117181 57621 117184
rect 57655 117181 57667 117215
rect 61746 117212 61752 117224
rect 61707 117184 61752 117212
rect 57609 117175 57667 117181
rect 61746 117172 61752 117184
rect 61804 117172 61810 117224
rect 66438 117212 66444 117224
rect 66399 117184 66444 117212
rect 66438 117172 66444 117184
rect 66496 117172 66502 117224
rect 71130 117212 71136 117224
rect 71091 117184 71136 117212
rect 71130 117172 71136 117184
rect 71188 117172 71194 117224
rect 75822 117172 75828 117224
rect 75880 117212 75886 117224
rect 76285 117215 76343 117221
rect 76285 117212 76297 117215
rect 75880 117184 76297 117212
rect 75880 117172 75886 117184
rect 76285 117181 76297 117184
rect 76331 117181 76343 117215
rect 76285 117175 76343 117181
rect 76926 117172 76932 117224
rect 76984 117212 76990 117224
rect 79336 117212 79364 117252
rect 80514 117212 80520 117224
rect 76984 117184 79364 117212
rect 80475 117184 80520 117212
rect 76984 117172 76990 117184
rect 80514 117172 80520 117184
rect 80572 117172 80578 117224
rect 80624 117212 80652 117252
rect 82078 117240 82084 117292
rect 82136 117280 82142 117292
rect 82357 117283 82415 117289
rect 82357 117280 82369 117283
rect 82136 117252 82369 117280
rect 82136 117240 82142 117252
rect 82357 117249 82369 117252
rect 82403 117249 82415 117283
rect 82357 117243 82415 117249
rect 83642 117240 83648 117292
rect 83700 117280 83706 117292
rect 84565 117283 84623 117289
rect 84565 117280 84577 117283
rect 83700 117252 84577 117280
rect 83700 117240 83706 117252
rect 84565 117249 84577 117252
rect 84611 117249 84623 117283
rect 84565 117243 84623 117249
rect 86954 117240 86960 117292
rect 87012 117280 87018 117292
rect 87233 117283 87291 117289
rect 87233 117280 87245 117283
rect 87012 117252 87245 117280
rect 87012 117240 87018 117252
rect 87233 117249 87245 117252
rect 87279 117249 87291 117283
rect 87233 117243 87291 117249
rect 88334 117240 88340 117292
rect 88392 117280 88398 117292
rect 88613 117283 88671 117289
rect 88613 117280 88625 117283
rect 88392 117252 88625 117280
rect 88392 117240 88398 117252
rect 88613 117249 88625 117252
rect 88659 117249 88671 117283
rect 88613 117243 88671 117249
rect 91554 117240 91560 117292
rect 91612 117280 91618 117292
rect 92569 117283 92627 117289
rect 92569 117280 92581 117283
rect 91612 117252 92581 117280
rect 91612 117240 91618 117252
rect 92569 117249 92581 117252
rect 92615 117249 92627 117283
rect 92569 117243 92627 117249
rect 93118 117240 93124 117292
rect 93176 117280 93182 117292
rect 93397 117283 93455 117289
rect 93397 117280 93409 117283
rect 93176 117252 93409 117280
rect 93176 117240 93182 117252
rect 93397 117249 93409 117252
rect 93443 117249 93455 117283
rect 93397 117243 93455 117249
rect 96246 117240 96252 117292
rect 96304 117280 96310 117292
rect 96525 117283 96583 117289
rect 96525 117280 96537 117283
rect 96304 117252 96537 117280
rect 96304 117240 96310 117252
rect 96525 117249 96537 117252
rect 96571 117249 96583 117283
rect 97810 117280 97816 117292
rect 97771 117252 97816 117280
rect 96525 117243 96583 117249
rect 97810 117240 97816 117252
rect 97868 117240 97874 117292
rect 100938 117240 100944 117292
rect 100996 117280 101002 117292
rect 101217 117283 101275 117289
rect 101217 117280 101229 117283
rect 100996 117252 101229 117280
rect 100996 117240 101002 117252
rect 101217 117249 101229 117252
rect 101263 117249 101275 117283
rect 101217 117243 101275 117249
rect 102502 117240 102508 117292
rect 102560 117280 102566 117292
rect 103241 117283 103299 117289
rect 103241 117280 103253 117283
rect 102560 117252 103253 117280
rect 102560 117240 102566 117252
rect 103241 117249 103253 117252
rect 103287 117249 103299 117283
rect 103241 117243 103299 117249
rect 105630 117240 105636 117292
rect 105688 117280 105694 117292
rect 105909 117283 105967 117289
rect 105909 117280 105921 117283
rect 105688 117252 105921 117280
rect 105688 117240 105694 117252
rect 105909 117249 105921 117252
rect 105955 117249 105967 117283
rect 105909 117243 105967 117249
rect 107194 117240 107200 117292
rect 107252 117280 107258 117292
rect 107381 117283 107439 117289
rect 107381 117280 107393 117283
rect 107252 117252 107393 117280
rect 107252 117240 107258 117252
rect 107381 117249 107393 117252
rect 107427 117249 107439 117283
rect 107381 117243 107439 117249
rect 110414 117240 110420 117292
rect 110472 117280 110478 117292
rect 111245 117283 111303 117289
rect 111245 117280 111257 117283
rect 110472 117252 111257 117280
rect 110472 117240 110478 117252
rect 111245 117249 111257 117252
rect 111291 117249 111303 117283
rect 111245 117243 111303 117249
rect 111886 117240 111892 117292
rect 111944 117280 111950 117292
rect 112165 117283 112223 117289
rect 112165 117280 112177 117283
rect 111944 117252 112177 117280
rect 111944 117240 111950 117252
rect 112165 117249 112177 117252
rect 112211 117249 112223 117283
rect 112165 117243 112223 117249
rect 115014 117240 115020 117292
rect 115072 117280 115078 117292
rect 115293 117283 115351 117289
rect 115293 117280 115305 117283
rect 115072 117252 115305 117280
rect 115072 117240 115078 117252
rect 115293 117249 115305 117252
rect 115339 117249 115351 117283
rect 115293 117243 115351 117249
rect 116578 117240 116584 117292
rect 116636 117280 116642 117292
rect 116857 117283 116915 117289
rect 116857 117280 116869 117283
rect 116636 117252 116869 117280
rect 116636 117240 116642 117252
rect 116857 117249 116869 117252
rect 116903 117249 116915 117283
rect 116857 117243 116915 117249
rect 119706 117240 119712 117292
rect 119764 117280 119770 117292
rect 119985 117283 120043 117289
rect 119985 117280 119997 117283
rect 119764 117252 119997 117280
rect 119764 117240 119770 117252
rect 119985 117249 119997 117252
rect 120031 117249 120043 117283
rect 119985 117243 120043 117249
rect 121454 117240 121460 117292
rect 121512 117280 121518 117292
rect 121917 117283 121975 117289
rect 121917 117280 121929 117283
rect 121512 117252 121929 117280
rect 121512 117240 121518 117252
rect 121917 117249 121929 117252
rect 121963 117249 121975 117283
rect 121917 117243 121975 117249
rect 124398 117240 124404 117292
rect 124456 117280 124462 117292
rect 124677 117283 124735 117289
rect 124677 117280 124689 117283
rect 124456 117252 124689 117280
rect 124456 117240 124462 117252
rect 124677 117249 124689 117252
rect 124723 117249 124735 117283
rect 124677 117243 124735 117249
rect 125962 117240 125968 117292
rect 126020 117280 126026 117292
rect 126057 117283 126115 117289
rect 126057 117280 126069 117283
rect 126020 117252 126069 117280
rect 126020 117240 126026 117252
rect 126057 117249 126069 117252
rect 126103 117249 126115 117283
rect 126057 117243 126115 117249
rect 129090 117240 129096 117292
rect 129148 117280 129154 117292
rect 129921 117283 129979 117289
rect 129921 117280 129933 117283
rect 129148 117252 129933 117280
rect 129148 117240 129154 117252
rect 129921 117249 129933 117252
rect 129967 117249 129979 117283
rect 129921 117243 129979 117249
rect 130654 117240 130660 117292
rect 130712 117280 130718 117292
rect 130933 117283 130991 117289
rect 130933 117280 130945 117283
rect 130712 117252 130945 117280
rect 130712 117240 130718 117252
rect 130933 117249 130945 117252
rect 130979 117249 130991 117283
rect 130933 117243 130991 117249
rect 133874 117240 133880 117292
rect 133932 117280 133938 117292
rect 134061 117283 134119 117289
rect 134061 117280 134073 117283
rect 133932 117252 134073 117280
rect 133932 117240 133938 117252
rect 134061 117249 134073 117252
rect 134107 117249 134119 117283
rect 134061 117243 134119 117249
rect 135346 117240 135352 117292
rect 135404 117280 135410 117292
rect 135625 117283 135683 117289
rect 135625 117280 135637 117283
rect 135404 117252 135637 117280
rect 135404 117240 135410 117252
rect 135625 117249 135637 117252
rect 135671 117249 135683 117283
rect 135625 117243 135683 117249
rect 138474 117240 138480 117292
rect 138532 117280 138538 117292
rect 138753 117283 138811 117289
rect 138753 117280 138765 117283
rect 138532 117252 138765 117280
rect 138532 117240 138538 117252
rect 138753 117249 138765 117252
rect 138799 117249 138811 117283
rect 138753 117243 138811 117249
rect 140038 117240 140044 117292
rect 140096 117280 140102 117292
rect 140593 117283 140651 117289
rect 140593 117280 140605 117283
rect 140096 117252 140605 117280
rect 140096 117240 140102 117252
rect 140593 117249 140605 117252
rect 140639 117249 140651 117283
rect 140593 117243 140651 117249
rect 143166 117240 143172 117292
rect 143224 117280 143230 117292
rect 143445 117283 143503 117289
rect 143445 117280 143457 117283
rect 143224 117252 143457 117280
rect 143224 117240 143230 117252
rect 143445 117249 143457 117252
rect 143491 117249 143503 117283
rect 144730 117280 144736 117292
rect 144691 117252 144736 117280
rect 143445 117243 143503 117249
rect 144730 117240 144736 117252
rect 144788 117240 144794 117292
rect 147858 117240 147864 117292
rect 147916 117280 147922 117292
rect 148597 117283 148655 117289
rect 148597 117280 148609 117283
rect 147916 117252 148609 117280
rect 147916 117240 147922 117252
rect 148597 117249 148609 117252
rect 148643 117249 148655 117283
rect 148597 117243 148655 117249
rect 149422 117240 149428 117292
rect 149480 117280 149486 117292
rect 149701 117283 149759 117289
rect 149701 117280 149713 117283
rect 149480 117252 149713 117280
rect 149480 117240 149486 117252
rect 149701 117249 149713 117252
rect 149747 117249 149759 117283
rect 149701 117243 149759 117249
rect 152550 117240 152556 117292
rect 152608 117280 152614 117292
rect 152737 117283 152795 117289
rect 152737 117280 152749 117283
rect 152608 117252 152749 117280
rect 152608 117240 152614 117252
rect 152737 117249 152749 117252
rect 152783 117249 152795 117283
rect 152737 117243 152795 117249
rect 154114 117240 154120 117292
rect 154172 117280 154178 117292
rect 154393 117283 154451 117289
rect 154393 117280 154405 117283
rect 154172 117252 154405 117280
rect 154172 117240 154178 117252
rect 154393 117249 154405 117252
rect 154439 117249 154451 117283
rect 154393 117243 154451 117249
rect 157334 117240 157340 117292
rect 157392 117280 157398 117292
rect 157521 117283 157579 117289
rect 157521 117280 157533 117283
rect 157392 117252 157533 117280
rect 157392 117240 157398 117252
rect 157521 117249 157533 117252
rect 157567 117249 157579 117283
rect 157521 117243 157579 117249
rect 158806 117240 158812 117292
rect 158864 117280 158870 117292
rect 159269 117283 159327 117289
rect 159269 117280 159281 117283
rect 158864 117252 159281 117280
rect 158864 117240 158870 117252
rect 159269 117249 159281 117252
rect 159315 117249 159327 117283
rect 159269 117243 159327 117249
rect 161934 117240 161940 117292
rect 161992 117280 161998 117292
rect 162213 117283 162271 117289
rect 162213 117280 162225 117283
rect 161992 117252 162225 117280
rect 161992 117240 161998 117252
rect 162213 117249 162225 117252
rect 162259 117249 162271 117283
rect 162213 117243 162271 117249
rect 163498 117240 163504 117292
rect 163556 117280 163562 117292
rect 164605 117283 164663 117289
rect 164605 117280 164617 117283
rect 163556 117252 164617 117280
rect 163556 117240 163562 117252
rect 164605 117249 164617 117252
rect 164651 117249 164663 117283
rect 164605 117243 164663 117249
rect 166626 117240 166632 117292
rect 166684 117280 166690 117292
rect 167273 117283 167331 117289
rect 167273 117280 167285 117283
rect 166684 117252 167285 117280
rect 166684 117240 166690 117252
rect 167273 117249 167285 117252
rect 167319 117249 167331 117283
rect 167273 117243 167331 117249
rect 168374 117240 168380 117292
rect 168432 117280 168438 117292
rect 168469 117283 168527 117289
rect 168469 117280 168481 117283
rect 168432 117252 168481 117280
rect 168432 117240 168438 117252
rect 168469 117249 168481 117252
rect 168515 117249 168527 117283
rect 168469 117243 168527 117249
rect 171318 117240 171324 117292
rect 171376 117280 171382 117292
rect 171413 117283 171471 117289
rect 171413 117280 171425 117283
rect 171376 117252 171425 117280
rect 171376 117240 171382 117252
rect 171413 117249 171425 117252
rect 171459 117249 171471 117283
rect 171413 117243 171471 117249
rect 172882 117240 172888 117292
rect 172940 117280 172946 117292
rect 173161 117283 173219 117289
rect 173161 117280 173173 117283
rect 172940 117252 173173 117280
rect 172940 117240 172946 117252
rect 173161 117249 173173 117252
rect 173207 117249 173219 117283
rect 173161 117243 173219 117249
rect 176010 117240 176016 117292
rect 176068 117280 176074 117292
rect 176289 117283 176347 117289
rect 176289 117280 176301 117283
rect 176068 117252 176301 117280
rect 176068 117240 176074 117252
rect 176289 117249 176301 117252
rect 176335 117249 176347 117283
rect 176289 117243 176347 117249
rect 177574 117240 177580 117292
rect 177632 117280 177638 117292
rect 177945 117283 178003 117289
rect 177945 117280 177957 117283
rect 177632 117252 177957 117280
rect 177632 117240 177638 117252
rect 177945 117249 177957 117252
rect 177991 117249 178003 117283
rect 177945 117243 178003 117249
rect 84381 117215 84439 117221
rect 84381 117212 84393 117215
rect 80624 117184 84393 117212
rect 84381 117181 84393 117184
rect 84427 117181 84439 117215
rect 85206 117212 85212 117224
rect 85167 117184 85212 117212
rect 84381 117175 84439 117181
rect 85206 117172 85212 117184
rect 85264 117172 85270 117224
rect 89898 117212 89904 117224
rect 89859 117184 89904 117212
rect 89898 117172 89904 117184
rect 89956 117172 89962 117224
rect 94682 117172 94688 117224
rect 94740 117212 94746 117224
rect 94961 117215 95019 117221
rect 94961 117212 94973 117215
rect 94740 117184 94973 117212
rect 94740 117172 94746 117184
rect 94961 117181 94973 117184
rect 95007 117181 95019 117215
rect 94961 117175 95019 117181
rect 97626 117172 97632 117224
rect 97684 117212 97690 117224
rect 97997 117215 98055 117221
rect 97997 117212 98009 117215
rect 97684 117184 98009 117212
rect 97684 117172 97690 117184
rect 97997 117181 98009 117184
rect 98043 117181 98055 117215
rect 97997 117175 98055 117181
rect 99193 117215 99251 117221
rect 99193 117181 99205 117215
rect 99239 117212 99251 117215
rect 99374 117212 99380 117224
rect 99239 117184 99380 117212
rect 99239 117181 99251 117184
rect 99193 117175 99251 117181
rect 99374 117172 99380 117184
rect 99432 117172 99438 117224
rect 104066 117212 104072 117224
rect 104027 117184 104072 117212
rect 104066 117172 104072 117184
rect 104124 117172 104130 117224
rect 108758 117212 108764 117224
rect 108719 117184 108764 117212
rect 108758 117172 108764 117184
rect 108816 117172 108822 117224
rect 113450 117172 113456 117224
rect 113508 117212 113514 117224
rect 113637 117215 113695 117221
rect 113637 117212 113649 117215
rect 113508 117184 113649 117212
rect 113508 117172 113514 117184
rect 113637 117181 113649 117184
rect 113683 117181 113695 117215
rect 113637 117175 113695 117181
rect 118142 117172 118148 117224
rect 118200 117212 118206 117224
rect 118973 117215 119031 117221
rect 118973 117212 118985 117215
rect 118200 117184 118985 117212
rect 118200 117172 118206 117184
rect 118973 117181 118985 117184
rect 119019 117181 119031 117215
rect 118973 117175 119031 117181
rect 122834 117172 122840 117224
rect 122892 117212 122898 117224
rect 127526 117212 127532 117224
rect 122892 117184 122937 117212
rect 127487 117184 127532 117212
rect 122892 117172 122898 117184
rect 127526 117172 127532 117184
rect 127584 117172 127590 117224
rect 132218 117172 132224 117224
rect 132276 117212 132282 117224
rect 132313 117215 132371 117221
rect 132313 117212 132325 117215
rect 132276 117184 132325 117212
rect 132276 117172 132282 117184
rect 132313 117181 132325 117184
rect 132359 117181 132371 117215
rect 132313 117175 132371 117181
rect 136910 117172 136916 117224
rect 136968 117212 136974 117224
rect 137649 117215 137707 117221
rect 137649 117212 137661 117215
rect 136968 117184 137661 117212
rect 136968 117172 136974 117184
rect 137649 117181 137661 117184
rect 137695 117181 137707 117215
rect 141602 117212 141608 117224
rect 141563 117184 141608 117212
rect 137649 117175 137707 117181
rect 141602 117172 141608 117184
rect 141660 117172 141666 117224
rect 146294 117212 146300 117224
rect 146255 117184 146300 117212
rect 146294 117172 146300 117184
rect 146352 117172 146358 117224
rect 150986 117212 150992 117224
rect 150947 117184 150992 117212
rect 150986 117172 150992 117184
rect 151044 117172 151050 117224
rect 155678 117172 155684 117224
rect 155736 117212 155742 117224
rect 156325 117215 156383 117221
rect 156325 117212 156337 117215
rect 155736 117184 156337 117212
rect 155736 117172 155742 117184
rect 156325 117181 156337 117184
rect 156371 117181 156383 117215
rect 160370 117212 160376 117224
rect 160331 117184 160376 117212
rect 156325 117175 156383 117181
rect 160370 117172 160376 117184
rect 160428 117172 160434 117224
rect 165062 117212 165068 117224
rect 165023 117184 165068 117212
rect 165062 117172 165068 117184
rect 165120 117172 165126 117224
rect 169754 117212 169760 117224
rect 169715 117184 169760 117212
rect 169754 117172 169760 117184
rect 169812 117172 169818 117224
rect 173897 117215 173955 117221
rect 173897 117181 173909 117215
rect 173943 117212 173955 117215
rect 174446 117212 174452 117224
rect 173943 117184 174452 117212
rect 173943 117181 173955 117184
rect 173897 117175 173955 117181
rect 174446 117172 174452 117184
rect 174504 117172 174510 117224
rect 175553 117215 175611 117221
rect 175553 117181 175565 117215
rect 175599 117212 175611 117215
rect 179138 117212 179144 117224
rect 175599 117184 179144 117212
rect 175599 117181 175611 117184
rect 175553 117175 175611 117181
rect 179138 117172 179144 117184
rect 179196 117172 179202 117224
rect 2406 117144 2412 117156
rect 2367 117116 2412 117144
rect 2406 117104 2412 117116
rect 2464 117104 2470 117156
rect 4338 117144 4344 117156
rect 4299 117116 4344 117144
rect 4338 117104 4344 117116
rect 4396 117104 4402 117156
rect 7101 117147 7159 117153
rect 7101 117113 7113 117147
rect 7147 117144 7159 117147
rect 8294 117144 8300 117156
rect 7147 117116 8300 117144
rect 7147 117113 7159 117116
rect 7101 117107 7159 117113
rect 8294 117104 8300 117116
rect 8352 117104 8358 117156
rect 8478 117144 8484 117156
rect 8439 117116 8484 117144
rect 8478 117104 8484 117116
rect 8536 117104 8542 117156
rect 12342 117144 12348 117156
rect 12303 117116 12348 117144
rect 12342 117104 12348 117116
rect 12400 117104 12406 117156
rect 13354 117144 13360 117156
rect 13315 117116 13360 117144
rect 13354 117104 13360 117116
rect 13412 117104 13418 117156
rect 16482 117144 16488 117156
rect 16443 117116 16488 117144
rect 16482 117104 16488 117116
rect 16540 117104 16546 117156
rect 18046 117144 18052 117156
rect 18007 117116 18052 117144
rect 18046 117104 18052 117116
rect 18104 117104 18110 117156
rect 21177 117147 21235 117153
rect 21177 117113 21189 117147
rect 21223 117144 21235 117147
rect 22554 117144 22560 117156
rect 21223 117116 22560 117144
rect 21223 117113 21235 117116
rect 21177 117107 21235 117113
rect 22554 117104 22560 117116
rect 22612 117104 22618 117156
rect 23014 117144 23020 117156
rect 22975 117116 23020 117144
rect 23014 117104 23020 117116
rect 23072 117104 23078 117156
rect 25869 117147 25927 117153
rect 25869 117113 25881 117147
rect 25915 117144 25927 117147
rect 26510 117144 26516 117156
rect 25915 117116 26516 117144
rect 25915 117113 25927 117116
rect 25869 117107 25927 117113
rect 26510 117104 26516 117116
rect 26568 117104 26574 117156
rect 27157 117147 27215 117153
rect 27157 117113 27169 117147
rect 27203 117113 27215 117147
rect 27157 117107 27215 117113
rect 27172 117076 27200 117107
rect 30834 117104 30840 117156
rect 30892 117144 30898 117156
rect 31021 117147 31079 117153
rect 31021 117144 31033 117147
rect 30892 117116 31033 117144
rect 30892 117104 30898 117116
rect 31021 117113 31033 117116
rect 31067 117113 31079 117147
rect 32122 117144 32128 117156
rect 32083 117116 32128 117144
rect 31021 117107 31079 117113
rect 32122 117104 32128 117116
rect 32180 117104 32186 117156
rect 36814 117144 36820 117156
rect 36775 117116 36820 117144
rect 36814 117104 36820 117116
rect 36872 117104 36878 117156
rect 39758 117104 39764 117156
rect 39816 117144 39822 117156
rect 39945 117147 40003 117153
rect 39945 117144 39957 117147
rect 39816 117116 39957 117144
rect 39816 117104 39822 117116
rect 39945 117113 39957 117116
rect 39991 117113 40003 117147
rect 41690 117144 41696 117156
rect 41651 117116 41696 117144
rect 39945 117107 40003 117113
rect 41690 117104 41696 117116
rect 41748 117104 41754 117156
rect 44358 117104 44364 117156
rect 44416 117144 44422 117156
rect 44637 117147 44695 117153
rect 44637 117144 44649 117147
rect 44416 117116 44649 117144
rect 44416 117104 44422 117116
rect 44637 117113 44649 117116
rect 44683 117113 44695 117147
rect 47026 117144 47032 117156
rect 46987 117116 47032 117144
rect 44637 117107 44695 117113
rect 47026 117104 47032 117116
rect 47084 117104 47090 117156
rect 48958 117104 48964 117156
rect 49016 117144 49022 117156
rect 49697 117147 49755 117153
rect 49697 117144 49709 117147
rect 49016 117116 49709 117144
rect 49016 117104 49022 117116
rect 49697 117113 49709 117116
rect 49743 117113 49755 117147
rect 50890 117144 50896 117156
rect 50851 117116 50896 117144
rect 49697 117107 49755 117113
rect 50890 117104 50896 117116
rect 50948 117104 50954 117156
rect 53837 117147 53895 117153
rect 53837 117113 53849 117147
rect 53883 117144 53895 117147
rect 54018 117144 54024 117156
rect 53883 117116 54024 117144
rect 53883 117113 53895 117116
rect 53837 117107 53895 117113
rect 54018 117104 54024 117116
rect 54076 117104 54082 117156
rect 55582 117144 55588 117156
rect 55543 117116 55588 117144
rect 55582 117104 55588 117116
rect 55640 117104 55646 117156
rect 58250 117104 58256 117156
rect 58308 117144 58314 117156
rect 58713 117147 58771 117153
rect 58713 117144 58725 117147
rect 58308 117116 58725 117144
rect 58308 117104 58314 117116
rect 58713 117113 58725 117116
rect 58759 117113 58771 117147
rect 60366 117144 60372 117156
rect 60327 117116 60372 117144
rect 58713 117107 58771 117113
rect 60366 117104 60372 117116
rect 60424 117104 60430 117156
rect 62942 117104 62948 117156
rect 63000 117144 63006 117156
rect 63405 117147 63463 117153
rect 63405 117144 63417 117147
rect 63000 117116 63417 117144
rect 63000 117104 63006 117116
rect 63405 117113 63417 117116
rect 63451 117113 63463 117147
rect 63405 117107 63463 117113
rect 65518 117104 65524 117156
rect 65576 117144 65582 117156
rect 65705 117147 65763 117153
rect 65705 117144 65717 117147
rect 65576 117116 65717 117144
rect 65576 117104 65582 117116
rect 65705 117113 65717 117116
rect 65751 117113 65763 117147
rect 65705 117107 65763 117113
rect 67634 117104 67640 117156
rect 67692 117144 67698 117156
rect 68373 117147 68431 117153
rect 68373 117144 68385 117147
rect 67692 117116 68385 117144
rect 67692 117104 67698 117116
rect 68373 117113 68385 117116
rect 68419 117113 68431 117147
rect 69658 117144 69664 117156
rect 69619 117116 69664 117144
rect 68373 117107 68431 117113
rect 69658 117104 69664 117116
rect 69716 117104 69722 117156
rect 72418 117104 72424 117156
rect 72476 117144 72482 117156
rect 72513 117147 72571 117153
rect 72513 117144 72525 117147
rect 72476 117116 72525 117144
rect 72476 117104 72482 117116
rect 72513 117113 72525 117116
rect 72559 117113 72571 117147
rect 74353 117147 74411 117153
rect 74353 117144 74365 117147
rect 72513 117107 72571 117113
rect 72620 117116 74365 117144
rect 33410 117076 33416 117088
rect 27172 117048 33416 117076
rect 33410 117036 33416 117048
rect 33468 117036 33474 117088
rect 69566 117036 69572 117088
rect 69624 117076 69630 117088
rect 72620 117076 72648 117116
rect 74353 117113 74365 117116
rect 74399 117113 74411 117147
rect 74353 117107 74411 117113
rect 77110 117104 77116 117156
rect 77168 117144 77174 117156
rect 77481 117147 77539 117153
rect 77481 117144 77493 117147
rect 77168 117116 77493 117144
rect 77168 117104 77174 117116
rect 77481 117113 77493 117116
rect 77527 117113 77539 117147
rect 79042 117144 79048 117156
rect 79003 117116 79048 117144
rect 77481 117107 77539 117113
rect 79042 117104 79048 117116
rect 79100 117104 79106 117156
rect 81802 117104 81808 117156
rect 81860 117144 81866 117156
rect 82173 117147 82231 117153
rect 82173 117144 82185 117147
rect 81860 117116 82185 117144
rect 81860 117104 81866 117116
rect 82173 117113 82185 117116
rect 82219 117113 82231 117147
rect 82173 117107 82231 117113
rect 86586 117104 86592 117156
rect 86644 117144 86650 117156
rect 87049 117147 87107 117153
rect 87049 117144 87061 117147
rect 86644 117116 87061 117144
rect 86644 117104 86650 117116
rect 87049 117113 87061 117116
rect 87095 117113 87107 117147
rect 88426 117144 88432 117156
rect 88387 117116 88432 117144
rect 87049 117107 87107 117113
rect 88426 117104 88432 117116
rect 88484 117104 88490 117156
rect 91370 117104 91376 117156
rect 91428 117144 91434 117156
rect 92385 117147 92443 117153
rect 92385 117144 92397 117147
rect 91428 117116 92397 117144
rect 91428 117104 91434 117116
rect 92385 117113 92397 117116
rect 92431 117113 92443 117147
rect 93210 117144 93216 117156
rect 93171 117116 93216 117144
rect 92385 117107 92443 117113
rect 93210 117104 93216 117116
rect 93268 117104 93274 117156
rect 96062 117104 96068 117156
rect 96120 117144 96126 117156
rect 96341 117147 96399 117153
rect 96341 117144 96353 117147
rect 96120 117116 96353 117144
rect 96120 117104 96126 117116
rect 96341 117113 96353 117116
rect 96387 117113 96399 117147
rect 101033 117147 101091 117153
rect 96341 117107 96399 117113
rect 97552 117116 97856 117144
rect 69624 117048 72648 117076
rect 69624 117036 69630 117048
rect 73062 117036 73068 117088
rect 73120 117076 73126 117088
rect 97552 117076 97580 117116
rect 73120 117048 97580 117076
rect 73120 117036 73126 117048
rect 97626 117036 97632 117088
rect 97684 117076 97690 117088
rect 97828 117076 97856 117116
rect 101033 117113 101045 117147
rect 101079 117144 101091 117147
rect 101214 117144 101220 117156
rect 101079 117116 101220 117144
rect 101079 117113 101091 117116
rect 101033 117107 101091 117113
rect 101214 117104 101220 117116
rect 101272 117104 101278 117156
rect 103054 117144 103060 117156
rect 103015 117116 103060 117144
rect 103054 117104 103060 117116
rect 103112 117104 103118 117156
rect 105354 117104 105360 117156
rect 105412 117144 105418 117156
rect 105725 117147 105783 117153
rect 105725 117144 105737 117147
rect 105412 117116 105737 117144
rect 105412 117104 105418 117116
rect 105725 117113 105737 117116
rect 105771 117113 105783 117147
rect 107194 117144 107200 117156
rect 107155 117116 107200 117144
rect 105725 117107 105783 117113
rect 107194 117104 107200 117116
rect 107252 117104 107258 117156
rect 110230 117104 110236 117156
rect 110288 117144 110294 117156
rect 111061 117147 111119 117153
rect 111061 117144 111073 117147
rect 110288 117116 111073 117144
rect 110288 117104 110294 117116
rect 111061 117113 111073 117116
rect 111107 117113 111119 117147
rect 111061 117107 111119 117113
rect 111150 117104 111156 117156
rect 111208 117144 111214 117156
rect 111981 117147 112039 117153
rect 111981 117144 111993 117147
rect 111208 117116 111993 117144
rect 111208 117104 111214 117116
rect 111981 117113 111993 117116
rect 112027 117113 112039 117147
rect 111981 117107 112039 117113
rect 114922 117104 114928 117156
rect 114980 117144 114986 117156
rect 115109 117147 115167 117153
rect 115109 117144 115121 117147
rect 114980 117116 115121 117144
rect 114980 117104 114986 117116
rect 115109 117113 115121 117116
rect 115155 117113 115167 117147
rect 116670 117144 116676 117156
rect 116631 117116 116676 117144
rect 115109 117107 115167 117113
rect 116670 117104 116676 117116
rect 116728 117104 116734 117156
rect 119614 117104 119620 117156
rect 119672 117144 119678 117156
rect 119801 117147 119859 117153
rect 119801 117144 119813 117147
rect 119672 117116 119813 117144
rect 119672 117104 119678 117116
rect 119801 117113 119813 117116
rect 119847 117113 119859 117147
rect 121730 117144 121736 117156
rect 121691 117116 121736 117144
rect 119801 117107 119859 117113
rect 121730 117104 121736 117116
rect 121788 117104 121794 117156
rect 124306 117104 124312 117156
rect 124364 117144 124370 117156
rect 124493 117147 124551 117153
rect 124493 117144 124505 117147
rect 124364 117116 124505 117144
rect 124364 117104 124370 117116
rect 124493 117113 124505 117116
rect 124539 117113 124551 117147
rect 124493 117107 124551 117113
rect 125873 117147 125931 117153
rect 125873 117113 125885 117147
rect 125919 117113 125931 117147
rect 125873 117107 125931 117113
rect 125888 117076 125916 117107
rect 128906 117104 128912 117156
rect 128964 117144 128970 117156
rect 129737 117147 129795 117153
rect 129737 117144 129749 117147
rect 128964 117116 129749 117144
rect 128964 117104 128970 117116
rect 129737 117113 129749 117116
rect 129783 117113 129795 117147
rect 130746 117144 130752 117156
rect 130707 117116 130752 117144
rect 129737 117107 129795 117113
rect 130746 117104 130752 117116
rect 130804 117104 130810 117156
rect 133506 117104 133512 117156
rect 133564 117144 133570 117156
rect 133877 117147 133935 117153
rect 133877 117144 133889 117147
rect 133564 117116 133889 117144
rect 133564 117104 133570 117116
rect 133877 117113 133889 117116
rect 133923 117113 133935 117147
rect 135438 117144 135444 117156
rect 135399 117116 135444 117144
rect 133877 117107 133935 117113
rect 135438 117104 135444 117116
rect 135496 117104 135502 117156
rect 138014 117104 138020 117156
rect 138072 117144 138078 117156
rect 138569 117147 138627 117153
rect 138569 117144 138581 117147
rect 138072 117116 138581 117144
rect 138072 117104 138078 117116
rect 138569 117113 138581 117116
rect 138615 117113 138627 117147
rect 140406 117144 140412 117156
rect 140367 117116 140412 117144
rect 138569 117107 138627 117113
rect 140406 117104 140412 117116
rect 140464 117104 140470 117156
rect 143166 117104 143172 117156
rect 143224 117144 143230 117156
rect 143261 117147 143319 117153
rect 143261 117144 143273 117147
rect 143224 117116 143273 117144
rect 143224 117104 143230 117116
rect 143261 117113 143273 117116
rect 143307 117113 143319 117147
rect 144546 117144 144552 117156
rect 144507 117116 144552 117144
rect 143261 117107 143319 117113
rect 144546 117104 144552 117116
rect 144604 117104 144610 117156
rect 146754 117104 146760 117156
rect 146812 117144 146818 117156
rect 148413 117147 148471 117153
rect 148413 117144 148425 117147
rect 146812 117116 148425 117144
rect 146812 117104 146818 117116
rect 148413 117113 148425 117116
rect 148459 117113 148471 117147
rect 149514 117144 149520 117156
rect 149475 117116 149520 117144
rect 148413 117107 148471 117113
rect 149514 117104 149520 117116
rect 149572 117104 149578 117156
rect 150894 117104 150900 117156
rect 150952 117144 150958 117156
rect 152553 117147 152611 117153
rect 152553 117144 152565 117147
rect 150952 117116 152565 117144
rect 150952 117104 150958 117116
rect 152553 117113 152565 117116
rect 152599 117113 152611 117147
rect 152553 117107 152611 117113
rect 154114 117104 154120 117156
rect 154172 117144 154178 117156
rect 154209 117147 154267 117153
rect 154209 117144 154221 117147
rect 154172 117116 154221 117144
rect 154172 117104 154178 117116
rect 154209 117113 154221 117116
rect 154255 117113 154267 117147
rect 154209 117107 154267 117113
rect 154850 117104 154856 117156
rect 154908 117144 154914 117156
rect 157337 117147 157395 117153
rect 157337 117144 157349 117147
rect 154908 117116 157349 117144
rect 154908 117104 154914 117116
rect 157337 117113 157349 117116
rect 157383 117113 157395 117147
rect 159082 117144 159088 117156
rect 159043 117116 159088 117144
rect 157337 117107 157395 117113
rect 159082 117104 159088 117116
rect 159140 117104 159146 117156
rect 162026 117144 162032 117156
rect 161987 117116 162032 117144
rect 162026 117104 162032 117116
rect 162084 117104 162090 117156
rect 164326 117104 164332 117156
rect 164384 117144 164390 117156
rect 164421 117147 164479 117153
rect 164421 117144 164433 117147
rect 164384 117116 164433 117144
rect 164384 117104 164390 117116
rect 164421 117113 164433 117116
rect 164467 117113 164479 117147
rect 164421 117107 164479 117113
rect 167089 117147 167147 117153
rect 167089 117113 167101 117147
rect 167135 117113 167147 117147
rect 167089 117107 167147 117113
rect 97684 117048 97729 117076
rect 97828 117048 125916 117076
rect 97684 117036 97690 117048
rect 162118 117036 162124 117088
rect 162176 117076 162182 117088
rect 167104 117076 167132 117107
rect 168190 117104 168196 117156
rect 168248 117144 168254 117156
rect 168285 117147 168343 117153
rect 168285 117144 168297 117147
rect 168248 117116 168297 117144
rect 168248 117104 168254 117116
rect 168285 117113 168297 117116
rect 168331 117113 168343 117147
rect 171226 117144 171232 117156
rect 171187 117116 171232 117144
rect 168285 117107 168343 117113
rect 171226 117104 171232 117116
rect 171284 117104 171290 117156
rect 172882 117104 172888 117156
rect 172940 117144 172946 117156
rect 172977 117147 173035 117153
rect 172977 117144 172989 117147
rect 172940 117116 172989 117144
rect 172940 117104 172946 117116
rect 172977 117113 172989 117116
rect 173023 117113 173035 117147
rect 172977 117107 173035 117113
rect 175369 117147 175427 117153
rect 175369 117113 175381 117147
rect 175415 117144 175427 117147
rect 175415 117116 175964 117144
rect 175415 117113 175427 117116
rect 175369 117107 175427 117113
rect 162176 117048 167132 117076
rect 175936 117076 175964 117116
rect 176010 117104 176016 117156
rect 176068 117144 176074 117156
rect 176105 117147 176163 117153
rect 176105 117144 176117 117147
rect 176068 117116 176117 117144
rect 176068 117104 176074 117116
rect 176105 117113 176117 117116
rect 176151 117113 176163 117147
rect 176105 117107 176163 117113
rect 176930 117104 176936 117156
rect 176988 117144 176994 117156
rect 177761 117147 177819 117153
rect 177761 117144 177773 117147
rect 176988 117116 177773 117144
rect 176988 117104 176994 117116
rect 177761 117113 177773 117116
rect 177807 117113 177819 117147
rect 177761 117107 177819 117113
rect 177574 117076 177580 117088
rect 175936 117048 177580 117076
rect 162176 117036 162182 117048
rect 177574 117036 177580 117048
rect 177632 117036 177638 117088
rect 1104 116986 178848 117008
rect 1104 116934 19606 116986
rect 19658 116934 19670 116986
rect 19722 116934 19734 116986
rect 19786 116934 19798 116986
rect 19850 116934 50326 116986
rect 50378 116934 50390 116986
rect 50442 116934 50454 116986
rect 50506 116934 50518 116986
rect 50570 116934 81046 116986
rect 81098 116934 81110 116986
rect 81162 116934 81174 116986
rect 81226 116934 81238 116986
rect 81290 116934 111766 116986
rect 111818 116934 111830 116986
rect 111882 116934 111894 116986
rect 111946 116934 111958 116986
rect 112010 116934 142486 116986
rect 142538 116934 142550 116986
rect 142602 116934 142614 116986
rect 142666 116934 142678 116986
rect 142730 116934 173206 116986
rect 173258 116934 173270 116986
rect 173322 116934 173334 116986
rect 173386 116934 173398 116986
rect 173450 116934 178848 116986
rect 1104 116912 178848 116934
rect 13354 116832 13360 116884
rect 13412 116872 13418 116884
rect 29270 116872 29276 116884
rect 13412 116844 29276 116872
rect 13412 116832 13418 116844
rect 29270 116832 29276 116844
rect 29328 116832 29334 116884
rect 58250 116872 58256 116884
rect 58211 116844 58256 116872
rect 58250 116832 58256 116844
rect 58308 116832 58314 116884
rect 68462 116832 68468 116884
rect 68520 116872 68526 116884
rect 111150 116872 111156 116884
rect 68520 116844 111156 116872
rect 68520 116832 68526 116844
rect 111150 116832 111156 116844
rect 111208 116832 111214 116884
rect 158625 116875 158683 116881
rect 158625 116841 158637 116875
rect 158671 116872 158683 116875
rect 162026 116872 162032 116884
rect 158671 116844 162032 116872
rect 158671 116841 158683 116844
rect 158625 116835 158683 116841
rect 162026 116832 162032 116844
rect 162084 116832 162090 116884
rect 18046 116764 18052 116816
rect 18104 116804 18110 116816
rect 29086 116804 29092 116816
rect 18104 116776 29092 116804
rect 18104 116764 18110 116776
rect 29086 116764 29092 116776
rect 29144 116764 29150 116816
rect 67818 116764 67824 116816
rect 67876 116804 67882 116816
rect 107194 116804 107200 116816
rect 67876 116776 107200 116804
rect 67876 116764 67882 116776
rect 107194 116764 107200 116776
rect 107252 116764 107258 116816
rect 4338 116696 4344 116748
rect 4396 116736 4402 116748
rect 26418 116736 26424 116748
rect 4396 116708 26424 116736
rect 4396 116696 4402 116708
rect 26418 116696 26424 116708
rect 26476 116696 26482 116748
rect 58434 116736 58440 116748
rect 58395 116708 58440 116736
rect 58434 116696 58440 116708
rect 58492 116696 58498 116748
rect 66070 116696 66076 116748
rect 66128 116736 66134 116748
rect 103054 116736 103060 116748
rect 66128 116708 103060 116736
rect 66128 116696 66134 116708
rect 103054 116696 103060 116708
rect 103112 116696 103118 116748
rect 158806 116736 158812 116748
rect 158767 116708 158812 116736
rect 158806 116696 158812 116708
rect 158864 116696 158870 116748
rect 23014 116628 23020 116680
rect 23072 116668 23078 116680
rect 31018 116668 31024 116680
rect 23072 116640 31024 116668
rect 23072 116628 23078 116640
rect 31018 116628 31024 116640
rect 31076 116628 31082 116680
rect 65242 116628 65248 116680
rect 65300 116668 65306 116680
rect 97626 116668 97632 116680
rect 65300 116640 97632 116668
rect 65300 116628 65306 116640
rect 97626 116628 97632 116640
rect 97684 116628 97690 116680
rect 8478 116560 8484 116612
rect 8536 116600 8542 116612
rect 26602 116600 26608 116612
rect 8536 116572 26608 116600
rect 8536 116560 8542 116572
rect 26602 116560 26608 116572
rect 26660 116560 26666 116612
rect 61010 116560 61016 116612
rect 61068 116600 61074 116612
rect 93210 116600 93216 116612
rect 61068 116572 93216 116600
rect 61068 116560 61074 116572
rect 93210 116560 93216 116572
rect 93268 116560 93274 116612
rect 60182 116492 60188 116544
rect 60240 116532 60246 116544
rect 88426 116532 88432 116544
rect 60240 116504 88432 116532
rect 60240 116492 60246 116504
rect 88426 116492 88432 116504
rect 88484 116492 88490 116544
rect 1104 116442 178848 116464
rect 1104 116390 4246 116442
rect 4298 116390 4310 116442
rect 4362 116390 4374 116442
rect 4426 116390 4438 116442
rect 4490 116390 34966 116442
rect 35018 116390 35030 116442
rect 35082 116390 35094 116442
rect 35146 116390 35158 116442
rect 35210 116390 65686 116442
rect 65738 116390 65750 116442
rect 65802 116390 65814 116442
rect 65866 116390 65878 116442
rect 65930 116390 96406 116442
rect 96458 116390 96470 116442
rect 96522 116390 96534 116442
rect 96586 116390 96598 116442
rect 96650 116390 127126 116442
rect 127178 116390 127190 116442
rect 127242 116390 127254 116442
rect 127306 116390 127318 116442
rect 127370 116390 157846 116442
rect 157898 116390 157910 116442
rect 157962 116390 157974 116442
rect 158026 116390 158038 116442
rect 158090 116390 178848 116442
rect 1104 116368 178848 116390
rect 2406 116288 2412 116340
rect 2464 116328 2470 116340
rect 7929 116331 7987 116337
rect 7929 116328 7941 116331
rect 2464 116300 7941 116328
rect 2464 116288 2470 116300
rect 7929 116297 7941 116300
rect 7975 116297 7987 116331
rect 7929 116291 7987 116297
rect 8294 116288 8300 116340
rect 8352 116328 8358 116340
rect 12069 116331 12127 116337
rect 12069 116328 12081 116331
rect 8352 116300 12081 116328
rect 8352 116288 8358 116300
rect 12069 116297 12081 116300
rect 12115 116297 12127 116331
rect 12069 116291 12127 116297
rect 12342 116288 12348 116340
rect 12400 116328 12406 116340
rect 14737 116331 14795 116337
rect 14737 116328 14749 116331
rect 12400 116300 14749 116328
rect 12400 116288 12406 116300
rect 14737 116297 14749 116300
rect 14783 116297 14795 116331
rect 14737 116291 14795 116297
rect 16482 116288 16488 116340
rect 16540 116328 16546 116340
rect 18509 116331 18567 116337
rect 18509 116328 18521 116331
rect 16540 116300 18521 116328
rect 16540 116288 16546 116300
rect 18509 116297 18521 116300
rect 18555 116297 18567 116331
rect 22554 116328 22560 116340
rect 22515 116300 22560 116328
rect 18509 116291 18567 116297
rect 22554 116288 22560 116300
rect 22612 116288 22618 116340
rect 26510 116288 26516 116340
rect 26568 116328 26574 116340
rect 26605 116331 26663 116337
rect 26605 116328 26617 116331
rect 26568 116300 26617 116328
rect 26568 116288 26574 116300
rect 26605 116297 26617 116300
rect 26651 116297 26663 116331
rect 30834 116328 30840 116340
rect 30795 116300 30840 116328
rect 26605 116291 26663 116297
rect 30834 116288 30840 116300
rect 30892 116288 30898 116340
rect 35250 116328 35256 116340
rect 35211 116300 35256 116328
rect 35250 116288 35256 116300
rect 35308 116288 35314 116340
rect 39758 116328 39764 116340
rect 39719 116300 39764 116328
rect 39758 116288 39764 116300
rect 39816 116288 39822 116340
rect 44358 116328 44364 116340
rect 44319 116300 44364 116328
rect 44358 116288 44364 116300
rect 44416 116288 44422 116340
rect 48958 116328 48964 116340
rect 48919 116300 48964 116328
rect 48958 116288 48964 116300
rect 49016 116288 49022 116340
rect 54018 116328 54024 116340
rect 53979 116300 54024 116328
rect 54018 116288 54024 116300
rect 54076 116288 54082 116340
rect 62942 116328 62948 116340
rect 62903 116300 62948 116328
rect 62942 116288 62948 116300
rect 63000 116288 63006 116340
rect 76926 116328 76932 116340
rect 63052 116300 76932 116328
rect 59262 116220 59268 116272
rect 59320 116260 59326 116272
rect 63052 116260 63080 116300
rect 76926 116288 76932 116300
rect 76984 116288 76990 116340
rect 77110 116328 77116 116340
rect 77071 116300 77116 116328
rect 77110 116288 77116 116300
rect 77168 116288 77174 116340
rect 81802 116328 81808 116340
rect 81763 116300 81808 116328
rect 81802 116288 81808 116300
rect 81860 116288 81866 116340
rect 86586 116328 86592 116340
rect 86547 116300 86592 116328
rect 86586 116288 86592 116300
rect 86644 116288 86650 116340
rect 91370 116328 91376 116340
rect 91331 116300 91376 116328
rect 91370 116288 91376 116300
rect 91428 116288 91434 116340
rect 96062 116328 96068 116340
rect 96023 116300 96068 116328
rect 96062 116288 96068 116300
rect 96120 116288 96126 116340
rect 101214 116328 101220 116340
rect 101175 116300 101220 116328
rect 101214 116288 101220 116300
rect 101272 116288 101278 116340
rect 105354 116328 105360 116340
rect 105315 116300 105360 116328
rect 105354 116288 105360 116300
rect 105412 116288 105418 116340
rect 110230 116328 110236 116340
rect 110191 116300 110236 116328
rect 110230 116288 110236 116300
rect 110288 116288 110294 116340
rect 114922 116328 114928 116340
rect 114883 116300 114928 116328
rect 114922 116288 114928 116300
rect 114980 116288 114986 116340
rect 119614 116328 119620 116340
rect 119575 116300 119620 116328
rect 119614 116288 119620 116300
rect 119672 116288 119678 116340
rect 124306 116328 124312 116340
rect 124267 116300 124312 116328
rect 124306 116288 124312 116300
rect 124364 116288 124370 116340
rect 128906 116328 128912 116340
rect 128867 116300 128912 116328
rect 128906 116288 128912 116300
rect 128964 116288 128970 116340
rect 133506 116328 133512 116340
rect 133467 116300 133512 116328
rect 133506 116288 133512 116300
rect 133564 116288 133570 116340
rect 138014 116328 138020 116340
rect 137975 116300 138020 116328
rect 138014 116288 138020 116300
rect 138072 116288 138078 116340
rect 143166 116328 143172 116340
rect 143127 116300 143172 116328
rect 143166 116288 143172 116300
rect 143224 116288 143230 116340
rect 146754 116328 146760 116340
rect 146715 116300 146760 116328
rect 146754 116288 146760 116300
rect 146812 116288 146818 116340
rect 150894 116328 150900 116340
rect 150855 116300 150900 116328
rect 150894 116288 150900 116300
rect 150952 116288 150958 116340
rect 154114 116328 154120 116340
rect 154075 116300 154120 116328
rect 154114 116288 154120 116300
rect 154172 116288 154178 116340
rect 154850 116328 154856 116340
rect 154811 116300 154856 116328
rect 154850 116288 154856 116300
rect 154908 116288 154914 116340
rect 159082 116328 159088 116340
rect 159043 116300 159088 116328
rect 159082 116288 159088 116300
rect 159140 116288 159146 116340
rect 162118 116328 162124 116340
rect 162079 116300 162124 116328
rect 162118 116288 162124 116300
rect 162176 116288 162182 116340
rect 164326 116328 164332 116340
rect 164287 116300 164332 116328
rect 164326 116288 164332 116300
rect 164384 116288 164390 116340
rect 168190 116328 168196 116340
rect 168151 116300 168196 116328
rect 168190 116288 168196 116300
rect 168248 116288 168254 116340
rect 172882 116328 172888 116340
rect 172843 116300 172888 116328
rect 172882 116288 172888 116300
rect 172940 116288 172946 116340
rect 176010 116328 176016 116340
rect 175971 116300 176016 116328
rect 176010 116288 176016 116300
rect 176068 116288 176074 116340
rect 176930 116328 176936 116340
rect 176891 116300 176936 116328
rect 176930 116288 176936 116300
rect 176988 116288 176994 116340
rect 177574 116328 177580 116340
rect 177535 116300 177580 116328
rect 177574 116288 177580 116300
rect 177632 116288 177638 116340
rect 67634 116260 67640 116272
rect 59320 116232 63080 116260
rect 67595 116232 67640 116260
rect 59320 116220 59326 116232
rect 67634 116220 67640 116232
rect 67692 116220 67698 116272
rect 72418 116260 72424 116272
rect 72379 116232 72424 116260
rect 72418 116220 72424 116232
rect 72476 116220 72482 116272
rect 79042 116260 79048 116272
rect 74506 116232 79048 116260
rect 49160 116164 55214 116192
rect 8113 116127 8171 116133
rect 8113 116093 8125 116127
rect 8159 116124 8171 116127
rect 12253 116127 12311 116133
rect 12253 116124 12265 116127
rect 8159 116096 12265 116124
rect 8159 116093 8171 116096
rect 8113 116087 8171 116093
rect 12253 116093 12265 116096
rect 12299 116124 12311 116127
rect 14921 116127 14979 116133
rect 14921 116124 14933 116127
rect 12299 116096 14933 116124
rect 12299 116093 12311 116096
rect 12253 116087 12311 116093
rect 14921 116093 14933 116096
rect 14967 116124 14979 116127
rect 18693 116127 18751 116133
rect 18693 116124 18705 116127
rect 14967 116096 18705 116124
rect 14967 116093 14979 116096
rect 14921 116087 14979 116093
rect 18693 116093 18705 116096
rect 18739 116124 18751 116127
rect 22741 116127 22799 116133
rect 22741 116124 22753 116127
rect 18739 116096 22753 116124
rect 18739 116093 18751 116096
rect 18693 116087 18751 116093
rect 22741 116093 22753 116096
rect 22787 116124 22799 116127
rect 26789 116127 26847 116133
rect 26789 116124 26801 116127
rect 22787 116096 26801 116124
rect 22787 116093 22799 116096
rect 22741 116087 22799 116093
rect 26789 116093 26801 116096
rect 26835 116124 26847 116127
rect 31021 116127 31079 116133
rect 31021 116124 31033 116127
rect 26835 116096 31033 116124
rect 26835 116093 26847 116096
rect 26789 116087 26847 116093
rect 31021 116093 31033 116096
rect 31067 116124 31079 116127
rect 31754 116124 31760 116136
rect 31067 116096 31760 116124
rect 31067 116093 31079 116096
rect 31021 116087 31079 116093
rect 31754 116084 31760 116096
rect 31812 116124 31818 116136
rect 49160 116133 49188 116164
rect 35437 116127 35495 116133
rect 35437 116124 35449 116127
rect 31812 116096 35449 116124
rect 31812 116084 31818 116096
rect 35437 116093 35449 116096
rect 35483 116124 35495 116127
rect 39945 116127 40003 116133
rect 39945 116124 39957 116127
rect 35483 116096 39957 116124
rect 35483 116093 35495 116096
rect 35437 116087 35495 116093
rect 39945 116093 39957 116096
rect 39991 116124 40003 116127
rect 44545 116127 44603 116133
rect 44545 116124 44557 116127
rect 39991 116096 44557 116124
rect 39991 116093 40003 116096
rect 39945 116087 40003 116093
rect 44545 116093 44557 116096
rect 44591 116124 44603 116127
rect 49145 116127 49203 116133
rect 49145 116124 49157 116127
rect 44591 116096 49157 116124
rect 44591 116093 44603 116096
rect 44545 116087 44603 116093
rect 49145 116093 49157 116096
rect 49191 116093 49203 116127
rect 49145 116087 49203 116093
rect 54205 116127 54263 116133
rect 54205 116093 54217 116127
rect 54251 116093 54263 116127
rect 55186 116124 55214 116164
rect 57146 116152 57152 116204
rect 57204 116192 57210 116204
rect 74506 116192 74534 116232
rect 79042 116220 79048 116232
rect 79100 116220 79106 116272
rect 57204 116164 74534 116192
rect 57204 116152 57210 116164
rect 56781 116127 56839 116133
rect 56781 116124 56793 116127
rect 55186 116096 56793 116124
rect 54205 116087 54263 116093
rect 56781 116093 56793 116096
rect 56827 116093 56839 116127
rect 57977 116127 58035 116133
rect 57977 116124 57989 116127
rect 56781 116087 56839 116093
rect 57808 116096 57989 116124
rect 54220 116056 54248 116087
rect 57808 116056 57836 116096
rect 57977 116093 57989 116096
rect 58023 116124 58035 116127
rect 58434 116124 58440 116136
rect 58023 116096 58440 116124
rect 58023 116093 58035 116096
rect 57977 116087 58035 116093
rect 58434 116084 58440 116096
rect 58492 116124 58498 116136
rect 63129 116127 63187 116133
rect 63129 116124 63141 116127
rect 58492 116096 63141 116124
rect 58492 116084 58498 116096
rect 63129 116093 63141 116096
rect 63175 116124 63187 116127
rect 67821 116127 67879 116133
rect 67821 116124 67833 116127
rect 63175 116096 67833 116124
rect 63175 116093 63187 116096
rect 63129 116087 63187 116093
rect 67821 116093 67833 116096
rect 67867 116124 67879 116127
rect 72605 116127 72663 116133
rect 72605 116124 72617 116127
rect 67867 116096 72617 116124
rect 67867 116093 67879 116096
rect 67821 116087 67879 116093
rect 72605 116093 72617 116096
rect 72651 116124 72663 116127
rect 77297 116127 77355 116133
rect 77297 116124 77309 116127
rect 72651 116096 77309 116124
rect 72651 116093 72663 116096
rect 72605 116087 72663 116093
rect 77297 116093 77309 116096
rect 77343 116124 77355 116127
rect 81989 116127 82047 116133
rect 81989 116124 82001 116127
rect 77343 116096 82001 116124
rect 77343 116093 77355 116096
rect 77297 116087 77355 116093
rect 81989 116093 82001 116096
rect 82035 116124 82047 116127
rect 86773 116127 86831 116133
rect 86773 116124 86785 116127
rect 82035 116096 86785 116124
rect 82035 116093 82047 116096
rect 81989 116087 82047 116093
rect 86773 116093 86785 116096
rect 86819 116124 86831 116127
rect 91557 116127 91615 116133
rect 91557 116124 91569 116127
rect 86819 116096 91569 116124
rect 86819 116093 86831 116096
rect 86773 116087 86831 116093
rect 91557 116093 91569 116096
rect 91603 116124 91615 116127
rect 96249 116127 96307 116133
rect 96249 116124 96261 116127
rect 91603 116096 96261 116124
rect 91603 116093 91615 116096
rect 91557 116087 91615 116093
rect 96249 116093 96261 116096
rect 96295 116124 96307 116127
rect 101401 116127 101459 116133
rect 101401 116124 101413 116127
rect 96295 116096 101413 116124
rect 96295 116093 96307 116096
rect 96249 116087 96307 116093
rect 101401 116093 101413 116096
rect 101447 116124 101459 116127
rect 105541 116127 105599 116133
rect 105541 116124 105553 116127
rect 101447 116096 105553 116124
rect 101447 116093 101459 116096
rect 101401 116087 101459 116093
rect 105541 116093 105553 116096
rect 105587 116124 105599 116127
rect 110417 116127 110475 116133
rect 110417 116124 110429 116127
rect 105587 116096 110429 116124
rect 105587 116093 105599 116096
rect 105541 116087 105599 116093
rect 110417 116093 110429 116096
rect 110463 116124 110475 116127
rect 115109 116127 115167 116133
rect 115109 116124 115121 116127
rect 110463 116096 115121 116124
rect 110463 116093 110475 116096
rect 110417 116087 110475 116093
rect 115109 116093 115121 116096
rect 115155 116124 115167 116127
rect 119801 116127 119859 116133
rect 119801 116124 119813 116127
rect 115155 116096 119813 116124
rect 115155 116093 115167 116096
rect 115109 116087 115167 116093
rect 119801 116093 119813 116096
rect 119847 116124 119859 116127
rect 124493 116127 124551 116133
rect 124493 116124 124505 116127
rect 119847 116096 124505 116124
rect 119847 116093 119859 116096
rect 119801 116087 119859 116093
rect 124493 116093 124505 116096
rect 124539 116124 124551 116127
rect 129093 116127 129151 116133
rect 129093 116124 129105 116127
rect 124539 116096 129105 116124
rect 124539 116093 124551 116096
rect 124493 116087 124551 116093
rect 129093 116093 129105 116096
rect 129139 116124 129151 116127
rect 133693 116127 133751 116133
rect 133693 116124 133705 116127
rect 129139 116096 133705 116124
rect 129139 116093 129151 116096
rect 129093 116087 129151 116093
rect 133693 116093 133705 116096
rect 133739 116124 133751 116127
rect 138201 116127 138259 116133
rect 138201 116124 138213 116127
rect 133739 116096 138213 116124
rect 133739 116093 133751 116096
rect 133693 116087 133751 116093
rect 138201 116093 138213 116096
rect 138247 116124 138259 116127
rect 143353 116127 143411 116133
rect 143353 116124 143365 116127
rect 138247 116096 143365 116124
rect 138247 116093 138259 116096
rect 138201 116087 138259 116093
rect 143353 116093 143365 116096
rect 143399 116124 143411 116127
rect 146941 116127 146999 116133
rect 146941 116124 146953 116127
rect 143399 116096 146953 116124
rect 143399 116093 143411 116096
rect 143353 116087 143411 116093
rect 146941 116093 146953 116096
rect 146987 116124 146999 116127
rect 151081 116127 151139 116133
rect 151081 116124 151093 116127
rect 146987 116096 151093 116124
rect 146987 116093 146999 116096
rect 146941 116087 146999 116093
rect 151081 116093 151093 116096
rect 151127 116124 151139 116127
rect 155037 116127 155095 116133
rect 155037 116124 155049 116127
rect 151127 116096 155049 116124
rect 151127 116093 151139 116096
rect 151081 116087 151139 116093
rect 155037 116093 155049 116096
rect 155083 116124 155095 116127
rect 158806 116124 158812 116136
rect 155083 116096 158812 116124
rect 155083 116093 155095 116096
rect 155037 116087 155095 116093
rect 158806 116084 158812 116096
rect 158864 116124 158870 116136
rect 162305 116127 162363 116133
rect 162305 116124 162317 116127
rect 158864 116096 162317 116124
rect 158864 116084 158870 116096
rect 162305 116093 162317 116096
rect 162351 116124 162363 116127
rect 171226 116124 171232 116136
rect 162351 116096 171232 116124
rect 162351 116093 162363 116096
rect 162305 116087 162363 116093
rect 171226 116084 171232 116096
rect 171284 116084 171290 116136
rect 69566 116056 69572 116068
rect 54220 116028 57836 116056
rect 57900 116028 69572 116056
rect 54202 115948 54208 116000
rect 54260 115988 54266 116000
rect 57900 115988 57928 116028
rect 69566 116016 69572 116028
rect 69624 116016 69630 116068
rect 72418 116016 72424 116068
rect 72476 116056 72482 116068
rect 116670 116056 116676 116068
rect 72476 116028 116676 116056
rect 72476 116016 72482 116028
rect 116670 116016 116676 116028
rect 116728 116016 116734 116068
rect 54260 115960 57928 115988
rect 54260 115948 54266 115960
rect 1104 115898 178848 115920
rect 1104 115846 19606 115898
rect 19658 115846 19670 115898
rect 19722 115846 19734 115898
rect 19786 115846 19798 115898
rect 19850 115846 50326 115898
rect 50378 115846 50390 115898
rect 50442 115846 50454 115898
rect 50506 115846 50518 115898
rect 50570 115846 81046 115898
rect 81098 115846 81110 115898
rect 81162 115846 81174 115898
rect 81226 115846 81238 115898
rect 81290 115846 111766 115898
rect 111818 115846 111830 115898
rect 111882 115846 111894 115898
rect 111946 115846 111958 115898
rect 112010 115846 142486 115898
rect 142538 115846 142550 115898
rect 142602 115846 142614 115898
rect 142666 115846 142678 115898
rect 142730 115846 173206 115898
rect 173258 115846 173270 115898
rect 173322 115846 173334 115898
rect 173386 115846 173398 115898
rect 173450 115846 178848 115898
rect 1104 115824 178848 115846
rect 1104 115354 178848 115376
rect 1104 115302 4246 115354
rect 4298 115302 4310 115354
rect 4362 115302 4374 115354
rect 4426 115302 4438 115354
rect 4490 115302 34966 115354
rect 35018 115302 35030 115354
rect 35082 115302 35094 115354
rect 35146 115302 35158 115354
rect 35210 115302 65686 115354
rect 65738 115302 65750 115354
rect 65802 115302 65814 115354
rect 65866 115302 65878 115354
rect 65930 115302 96406 115354
rect 96458 115302 96470 115354
rect 96522 115302 96534 115354
rect 96586 115302 96598 115354
rect 96650 115302 127126 115354
rect 127178 115302 127190 115354
rect 127242 115302 127254 115354
rect 127306 115302 127318 115354
rect 127370 115302 157846 115354
rect 157898 115302 157910 115354
rect 157962 115302 157974 115354
rect 158026 115302 158038 115354
rect 158090 115302 178848 115354
rect 1104 115280 178848 115302
rect 1104 114810 178848 114832
rect 1104 114758 19606 114810
rect 19658 114758 19670 114810
rect 19722 114758 19734 114810
rect 19786 114758 19798 114810
rect 19850 114758 50326 114810
rect 50378 114758 50390 114810
rect 50442 114758 50454 114810
rect 50506 114758 50518 114810
rect 50570 114758 81046 114810
rect 81098 114758 81110 114810
rect 81162 114758 81174 114810
rect 81226 114758 81238 114810
rect 81290 114758 111766 114810
rect 111818 114758 111830 114810
rect 111882 114758 111894 114810
rect 111946 114758 111958 114810
rect 112010 114758 142486 114810
rect 142538 114758 142550 114810
rect 142602 114758 142614 114810
rect 142666 114758 142678 114810
rect 142730 114758 173206 114810
rect 173258 114758 173270 114810
rect 173322 114758 173334 114810
rect 173386 114758 173398 114810
rect 173450 114758 178848 114810
rect 1104 114736 178848 114758
rect 1104 114266 178848 114288
rect 1104 114214 4246 114266
rect 4298 114214 4310 114266
rect 4362 114214 4374 114266
rect 4426 114214 4438 114266
rect 4490 114214 34966 114266
rect 35018 114214 35030 114266
rect 35082 114214 35094 114266
rect 35146 114214 35158 114266
rect 35210 114214 65686 114266
rect 65738 114214 65750 114266
rect 65802 114214 65814 114266
rect 65866 114214 65878 114266
rect 65930 114214 96406 114266
rect 96458 114214 96470 114266
rect 96522 114214 96534 114266
rect 96586 114214 96598 114266
rect 96650 114214 127126 114266
rect 127178 114214 127190 114266
rect 127242 114214 127254 114266
rect 127306 114214 127318 114266
rect 127370 114214 157846 114266
rect 157898 114214 157910 114266
rect 157962 114214 157974 114266
rect 158026 114214 158038 114266
rect 158090 114214 178848 114266
rect 1104 114192 178848 114214
rect 1104 113722 178848 113744
rect 1104 113670 19606 113722
rect 19658 113670 19670 113722
rect 19722 113670 19734 113722
rect 19786 113670 19798 113722
rect 19850 113670 50326 113722
rect 50378 113670 50390 113722
rect 50442 113670 50454 113722
rect 50506 113670 50518 113722
rect 50570 113670 81046 113722
rect 81098 113670 81110 113722
rect 81162 113670 81174 113722
rect 81226 113670 81238 113722
rect 81290 113670 111766 113722
rect 111818 113670 111830 113722
rect 111882 113670 111894 113722
rect 111946 113670 111958 113722
rect 112010 113670 142486 113722
rect 142538 113670 142550 113722
rect 142602 113670 142614 113722
rect 142666 113670 142678 113722
rect 142730 113670 173206 113722
rect 173258 113670 173270 113722
rect 173322 113670 173334 113722
rect 173386 113670 173398 113722
rect 173450 113670 178848 113722
rect 1104 113648 178848 113670
rect 1104 113178 178848 113200
rect 1104 113126 4246 113178
rect 4298 113126 4310 113178
rect 4362 113126 4374 113178
rect 4426 113126 4438 113178
rect 4490 113126 34966 113178
rect 35018 113126 35030 113178
rect 35082 113126 35094 113178
rect 35146 113126 35158 113178
rect 35210 113126 65686 113178
rect 65738 113126 65750 113178
rect 65802 113126 65814 113178
rect 65866 113126 65878 113178
rect 65930 113126 96406 113178
rect 96458 113126 96470 113178
rect 96522 113126 96534 113178
rect 96586 113126 96598 113178
rect 96650 113126 127126 113178
rect 127178 113126 127190 113178
rect 127242 113126 127254 113178
rect 127306 113126 127318 113178
rect 127370 113126 157846 113178
rect 157898 113126 157910 113178
rect 157962 113126 157974 113178
rect 158026 113126 158038 113178
rect 158090 113126 178848 113178
rect 1104 113104 178848 113126
rect 1104 112634 178848 112656
rect 1104 112582 19606 112634
rect 19658 112582 19670 112634
rect 19722 112582 19734 112634
rect 19786 112582 19798 112634
rect 19850 112582 50326 112634
rect 50378 112582 50390 112634
rect 50442 112582 50454 112634
rect 50506 112582 50518 112634
rect 50570 112582 81046 112634
rect 81098 112582 81110 112634
rect 81162 112582 81174 112634
rect 81226 112582 81238 112634
rect 81290 112582 111766 112634
rect 111818 112582 111830 112634
rect 111882 112582 111894 112634
rect 111946 112582 111958 112634
rect 112010 112582 142486 112634
rect 142538 112582 142550 112634
rect 142602 112582 142614 112634
rect 142666 112582 142678 112634
rect 142730 112582 173206 112634
rect 173258 112582 173270 112634
rect 173322 112582 173334 112634
rect 173386 112582 173398 112634
rect 173450 112582 178848 112634
rect 1104 112560 178848 112582
rect 1104 112090 178848 112112
rect 1104 112038 4246 112090
rect 4298 112038 4310 112090
rect 4362 112038 4374 112090
rect 4426 112038 4438 112090
rect 4490 112038 34966 112090
rect 35018 112038 35030 112090
rect 35082 112038 35094 112090
rect 35146 112038 35158 112090
rect 35210 112038 65686 112090
rect 65738 112038 65750 112090
rect 65802 112038 65814 112090
rect 65866 112038 65878 112090
rect 65930 112038 96406 112090
rect 96458 112038 96470 112090
rect 96522 112038 96534 112090
rect 96586 112038 96598 112090
rect 96650 112038 127126 112090
rect 127178 112038 127190 112090
rect 127242 112038 127254 112090
rect 127306 112038 127318 112090
rect 127370 112038 157846 112090
rect 157898 112038 157910 112090
rect 157962 112038 157974 112090
rect 158026 112038 158038 112090
rect 158090 112038 178848 112090
rect 1104 112016 178848 112038
rect 1104 111546 178848 111568
rect 1104 111494 19606 111546
rect 19658 111494 19670 111546
rect 19722 111494 19734 111546
rect 19786 111494 19798 111546
rect 19850 111494 50326 111546
rect 50378 111494 50390 111546
rect 50442 111494 50454 111546
rect 50506 111494 50518 111546
rect 50570 111494 81046 111546
rect 81098 111494 81110 111546
rect 81162 111494 81174 111546
rect 81226 111494 81238 111546
rect 81290 111494 111766 111546
rect 111818 111494 111830 111546
rect 111882 111494 111894 111546
rect 111946 111494 111958 111546
rect 112010 111494 142486 111546
rect 142538 111494 142550 111546
rect 142602 111494 142614 111546
rect 142666 111494 142678 111546
rect 142730 111494 173206 111546
rect 173258 111494 173270 111546
rect 173322 111494 173334 111546
rect 173386 111494 173398 111546
rect 173450 111494 178848 111546
rect 1104 111472 178848 111494
rect 1104 111002 178848 111024
rect 1104 110950 4246 111002
rect 4298 110950 4310 111002
rect 4362 110950 4374 111002
rect 4426 110950 4438 111002
rect 4490 110950 34966 111002
rect 35018 110950 35030 111002
rect 35082 110950 35094 111002
rect 35146 110950 35158 111002
rect 35210 110950 65686 111002
rect 65738 110950 65750 111002
rect 65802 110950 65814 111002
rect 65866 110950 65878 111002
rect 65930 110950 96406 111002
rect 96458 110950 96470 111002
rect 96522 110950 96534 111002
rect 96586 110950 96598 111002
rect 96650 110950 127126 111002
rect 127178 110950 127190 111002
rect 127242 110950 127254 111002
rect 127306 110950 127318 111002
rect 127370 110950 157846 111002
rect 157898 110950 157910 111002
rect 157962 110950 157974 111002
rect 158026 110950 158038 111002
rect 158090 110950 178848 111002
rect 1104 110928 178848 110950
rect 1104 110458 178848 110480
rect 1104 110406 19606 110458
rect 19658 110406 19670 110458
rect 19722 110406 19734 110458
rect 19786 110406 19798 110458
rect 19850 110406 50326 110458
rect 50378 110406 50390 110458
rect 50442 110406 50454 110458
rect 50506 110406 50518 110458
rect 50570 110406 81046 110458
rect 81098 110406 81110 110458
rect 81162 110406 81174 110458
rect 81226 110406 81238 110458
rect 81290 110406 111766 110458
rect 111818 110406 111830 110458
rect 111882 110406 111894 110458
rect 111946 110406 111958 110458
rect 112010 110406 142486 110458
rect 142538 110406 142550 110458
rect 142602 110406 142614 110458
rect 142666 110406 142678 110458
rect 142730 110406 173206 110458
rect 173258 110406 173270 110458
rect 173322 110406 173334 110458
rect 173386 110406 173398 110458
rect 173450 110406 178848 110458
rect 1104 110384 178848 110406
rect 1104 109914 178848 109936
rect 1104 109862 4246 109914
rect 4298 109862 4310 109914
rect 4362 109862 4374 109914
rect 4426 109862 4438 109914
rect 4490 109862 34966 109914
rect 35018 109862 35030 109914
rect 35082 109862 35094 109914
rect 35146 109862 35158 109914
rect 35210 109862 65686 109914
rect 65738 109862 65750 109914
rect 65802 109862 65814 109914
rect 65866 109862 65878 109914
rect 65930 109862 96406 109914
rect 96458 109862 96470 109914
rect 96522 109862 96534 109914
rect 96586 109862 96598 109914
rect 96650 109862 127126 109914
rect 127178 109862 127190 109914
rect 127242 109862 127254 109914
rect 127306 109862 127318 109914
rect 127370 109862 157846 109914
rect 157898 109862 157910 109914
rect 157962 109862 157974 109914
rect 158026 109862 158038 109914
rect 158090 109862 178848 109914
rect 1104 109840 178848 109862
rect 1104 109370 178848 109392
rect 1104 109318 19606 109370
rect 19658 109318 19670 109370
rect 19722 109318 19734 109370
rect 19786 109318 19798 109370
rect 19850 109318 50326 109370
rect 50378 109318 50390 109370
rect 50442 109318 50454 109370
rect 50506 109318 50518 109370
rect 50570 109318 81046 109370
rect 81098 109318 81110 109370
rect 81162 109318 81174 109370
rect 81226 109318 81238 109370
rect 81290 109318 111766 109370
rect 111818 109318 111830 109370
rect 111882 109318 111894 109370
rect 111946 109318 111958 109370
rect 112010 109318 142486 109370
rect 142538 109318 142550 109370
rect 142602 109318 142614 109370
rect 142666 109318 142678 109370
rect 142730 109318 173206 109370
rect 173258 109318 173270 109370
rect 173322 109318 173334 109370
rect 173386 109318 173398 109370
rect 173450 109318 178848 109370
rect 1104 109296 178848 109318
rect 1104 108826 178848 108848
rect 1104 108774 4246 108826
rect 4298 108774 4310 108826
rect 4362 108774 4374 108826
rect 4426 108774 4438 108826
rect 4490 108774 34966 108826
rect 35018 108774 35030 108826
rect 35082 108774 35094 108826
rect 35146 108774 35158 108826
rect 35210 108774 65686 108826
rect 65738 108774 65750 108826
rect 65802 108774 65814 108826
rect 65866 108774 65878 108826
rect 65930 108774 96406 108826
rect 96458 108774 96470 108826
rect 96522 108774 96534 108826
rect 96586 108774 96598 108826
rect 96650 108774 127126 108826
rect 127178 108774 127190 108826
rect 127242 108774 127254 108826
rect 127306 108774 127318 108826
rect 127370 108774 157846 108826
rect 157898 108774 157910 108826
rect 157962 108774 157974 108826
rect 158026 108774 158038 108826
rect 158090 108774 178848 108826
rect 1104 108752 178848 108774
rect 1104 108282 178848 108304
rect 1104 108230 19606 108282
rect 19658 108230 19670 108282
rect 19722 108230 19734 108282
rect 19786 108230 19798 108282
rect 19850 108230 50326 108282
rect 50378 108230 50390 108282
rect 50442 108230 50454 108282
rect 50506 108230 50518 108282
rect 50570 108230 81046 108282
rect 81098 108230 81110 108282
rect 81162 108230 81174 108282
rect 81226 108230 81238 108282
rect 81290 108230 111766 108282
rect 111818 108230 111830 108282
rect 111882 108230 111894 108282
rect 111946 108230 111958 108282
rect 112010 108230 142486 108282
rect 142538 108230 142550 108282
rect 142602 108230 142614 108282
rect 142666 108230 142678 108282
rect 142730 108230 173206 108282
rect 173258 108230 173270 108282
rect 173322 108230 173334 108282
rect 173386 108230 173398 108282
rect 173450 108230 178848 108282
rect 1104 108208 178848 108230
rect 1104 107738 178848 107760
rect 1104 107686 4246 107738
rect 4298 107686 4310 107738
rect 4362 107686 4374 107738
rect 4426 107686 4438 107738
rect 4490 107686 34966 107738
rect 35018 107686 35030 107738
rect 35082 107686 35094 107738
rect 35146 107686 35158 107738
rect 35210 107686 65686 107738
rect 65738 107686 65750 107738
rect 65802 107686 65814 107738
rect 65866 107686 65878 107738
rect 65930 107686 96406 107738
rect 96458 107686 96470 107738
rect 96522 107686 96534 107738
rect 96586 107686 96598 107738
rect 96650 107686 127126 107738
rect 127178 107686 127190 107738
rect 127242 107686 127254 107738
rect 127306 107686 127318 107738
rect 127370 107686 157846 107738
rect 157898 107686 157910 107738
rect 157962 107686 157974 107738
rect 158026 107686 158038 107738
rect 158090 107686 178848 107738
rect 1104 107664 178848 107686
rect 1104 107194 178848 107216
rect 1104 107142 19606 107194
rect 19658 107142 19670 107194
rect 19722 107142 19734 107194
rect 19786 107142 19798 107194
rect 19850 107142 50326 107194
rect 50378 107142 50390 107194
rect 50442 107142 50454 107194
rect 50506 107142 50518 107194
rect 50570 107142 81046 107194
rect 81098 107142 81110 107194
rect 81162 107142 81174 107194
rect 81226 107142 81238 107194
rect 81290 107142 111766 107194
rect 111818 107142 111830 107194
rect 111882 107142 111894 107194
rect 111946 107142 111958 107194
rect 112010 107142 142486 107194
rect 142538 107142 142550 107194
rect 142602 107142 142614 107194
rect 142666 107142 142678 107194
rect 142730 107142 173206 107194
rect 173258 107142 173270 107194
rect 173322 107142 173334 107194
rect 173386 107142 173398 107194
rect 173450 107142 178848 107194
rect 1104 107120 178848 107142
rect 1104 106650 178848 106672
rect 1104 106598 4246 106650
rect 4298 106598 4310 106650
rect 4362 106598 4374 106650
rect 4426 106598 4438 106650
rect 4490 106598 34966 106650
rect 35018 106598 35030 106650
rect 35082 106598 35094 106650
rect 35146 106598 35158 106650
rect 35210 106598 65686 106650
rect 65738 106598 65750 106650
rect 65802 106598 65814 106650
rect 65866 106598 65878 106650
rect 65930 106598 96406 106650
rect 96458 106598 96470 106650
rect 96522 106598 96534 106650
rect 96586 106598 96598 106650
rect 96650 106598 127126 106650
rect 127178 106598 127190 106650
rect 127242 106598 127254 106650
rect 127306 106598 127318 106650
rect 127370 106598 157846 106650
rect 157898 106598 157910 106650
rect 157962 106598 157974 106650
rect 158026 106598 158038 106650
rect 158090 106598 178848 106650
rect 1104 106576 178848 106598
rect 1104 106106 178848 106128
rect 1104 106054 19606 106106
rect 19658 106054 19670 106106
rect 19722 106054 19734 106106
rect 19786 106054 19798 106106
rect 19850 106054 50326 106106
rect 50378 106054 50390 106106
rect 50442 106054 50454 106106
rect 50506 106054 50518 106106
rect 50570 106054 81046 106106
rect 81098 106054 81110 106106
rect 81162 106054 81174 106106
rect 81226 106054 81238 106106
rect 81290 106054 111766 106106
rect 111818 106054 111830 106106
rect 111882 106054 111894 106106
rect 111946 106054 111958 106106
rect 112010 106054 142486 106106
rect 142538 106054 142550 106106
rect 142602 106054 142614 106106
rect 142666 106054 142678 106106
rect 142730 106054 173206 106106
rect 173258 106054 173270 106106
rect 173322 106054 173334 106106
rect 173386 106054 173398 106106
rect 173450 106054 178848 106106
rect 1104 106032 178848 106054
rect 1104 105562 178848 105584
rect 1104 105510 4246 105562
rect 4298 105510 4310 105562
rect 4362 105510 4374 105562
rect 4426 105510 4438 105562
rect 4490 105510 34966 105562
rect 35018 105510 35030 105562
rect 35082 105510 35094 105562
rect 35146 105510 35158 105562
rect 35210 105510 65686 105562
rect 65738 105510 65750 105562
rect 65802 105510 65814 105562
rect 65866 105510 65878 105562
rect 65930 105510 96406 105562
rect 96458 105510 96470 105562
rect 96522 105510 96534 105562
rect 96586 105510 96598 105562
rect 96650 105510 127126 105562
rect 127178 105510 127190 105562
rect 127242 105510 127254 105562
rect 127306 105510 127318 105562
rect 127370 105510 157846 105562
rect 157898 105510 157910 105562
rect 157962 105510 157974 105562
rect 158026 105510 158038 105562
rect 158090 105510 178848 105562
rect 1104 105488 178848 105510
rect 1104 105018 178848 105040
rect 1104 104966 19606 105018
rect 19658 104966 19670 105018
rect 19722 104966 19734 105018
rect 19786 104966 19798 105018
rect 19850 104966 50326 105018
rect 50378 104966 50390 105018
rect 50442 104966 50454 105018
rect 50506 104966 50518 105018
rect 50570 104966 81046 105018
rect 81098 104966 81110 105018
rect 81162 104966 81174 105018
rect 81226 104966 81238 105018
rect 81290 104966 111766 105018
rect 111818 104966 111830 105018
rect 111882 104966 111894 105018
rect 111946 104966 111958 105018
rect 112010 104966 142486 105018
rect 142538 104966 142550 105018
rect 142602 104966 142614 105018
rect 142666 104966 142678 105018
rect 142730 104966 173206 105018
rect 173258 104966 173270 105018
rect 173322 104966 173334 105018
rect 173386 104966 173398 105018
rect 173450 104966 178848 105018
rect 1104 104944 178848 104966
rect 1104 104474 178848 104496
rect 1104 104422 4246 104474
rect 4298 104422 4310 104474
rect 4362 104422 4374 104474
rect 4426 104422 4438 104474
rect 4490 104422 34966 104474
rect 35018 104422 35030 104474
rect 35082 104422 35094 104474
rect 35146 104422 35158 104474
rect 35210 104422 65686 104474
rect 65738 104422 65750 104474
rect 65802 104422 65814 104474
rect 65866 104422 65878 104474
rect 65930 104422 96406 104474
rect 96458 104422 96470 104474
rect 96522 104422 96534 104474
rect 96586 104422 96598 104474
rect 96650 104422 127126 104474
rect 127178 104422 127190 104474
rect 127242 104422 127254 104474
rect 127306 104422 127318 104474
rect 127370 104422 157846 104474
rect 157898 104422 157910 104474
rect 157962 104422 157974 104474
rect 158026 104422 158038 104474
rect 158090 104422 178848 104474
rect 1104 104400 178848 104422
rect 1104 103930 178848 103952
rect 1104 103878 19606 103930
rect 19658 103878 19670 103930
rect 19722 103878 19734 103930
rect 19786 103878 19798 103930
rect 19850 103878 50326 103930
rect 50378 103878 50390 103930
rect 50442 103878 50454 103930
rect 50506 103878 50518 103930
rect 50570 103878 81046 103930
rect 81098 103878 81110 103930
rect 81162 103878 81174 103930
rect 81226 103878 81238 103930
rect 81290 103878 111766 103930
rect 111818 103878 111830 103930
rect 111882 103878 111894 103930
rect 111946 103878 111958 103930
rect 112010 103878 142486 103930
rect 142538 103878 142550 103930
rect 142602 103878 142614 103930
rect 142666 103878 142678 103930
rect 142730 103878 173206 103930
rect 173258 103878 173270 103930
rect 173322 103878 173334 103930
rect 173386 103878 173398 103930
rect 173450 103878 178848 103930
rect 1104 103856 178848 103878
rect 1104 103386 178848 103408
rect 1104 103334 4246 103386
rect 4298 103334 4310 103386
rect 4362 103334 4374 103386
rect 4426 103334 4438 103386
rect 4490 103334 34966 103386
rect 35018 103334 35030 103386
rect 35082 103334 35094 103386
rect 35146 103334 35158 103386
rect 35210 103334 65686 103386
rect 65738 103334 65750 103386
rect 65802 103334 65814 103386
rect 65866 103334 65878 103386
rect 65930 103334 96406 103386
rect 96458 103334 96470 103386
rect 96522 103334 96534 103386
rect 96586 103334 96598 103386
rect 96650 103334 127126 103386
rect 127178 103334 127190 103386
rect 127242 103334 127254 103386
rect 127306 103334 127318 103386
rect 127370 103334 157846 103386
rect 157898 103334 157910 103386
rect 157962 103334 157974 103386
rect 158026 103334 158038 103386
rect 158090 103334 178848 103386
rect 1104 103312 178848 103334
rect 1104 102842 178848 102864
rect 1104 102790 19606 102842
rect 19658 102790 19670 102842
rect 19722 102790 19734 102842
rect 19786 102790 19798 102842
rect 19850 102790 50326 102842
rect 50378 102790 50390 102842
rect 50442 102790 50454 102842
rect 50506 102790 50518 102842
rect 50570 102790 81046 102842
rect 81098 102790 81110 102842
rect 81162 102790 81174 102842
rect 81226 102790 81238 102842
rect 81290 102790 111766 102842
rect 111818 102790 111830 102842
rect 111882 102790 111894 102842
rect 111946 102790 111958 102842
rect 112010 102790 142486 102842
rect 142538 102790 142550 102842
rect 142602 102790 142614 102842
rect 142666 102790 142678 102842
rect 142730 102790 173206 102842
rect 173258 102790 173270 102842
rect 173322 102790 173334 102842
rect 173386 102790 173398 102842
rect 173450 102790 178848 102842
rect 1104 102768 178848 102790
rect 1104 102298 178848 102320
rect 1104 102246 4246 102298
rect 4298 102246 4310 102298
rect 4362 102246 4374 102298
rect 4426 102246 4438 102298
rect 4490 102246 34966 102298
rect 35018 102246 35030 102298
rect 35082 102246 35094 102298
rect 35146 102246 35158 102298
rect 35210 102246 65686 102298
rect 65738 102246 65750 102298
rect 65802 102246 65814 102298
rect 65866 102246 65878 102298
rect 65930 102246 96406 102298
rect 96458 102246 96470 102298
rect 96522 102246 96534 102298
rect 96586 102246 96598 102298
rect 96650 102246 127126 102298
rect 127178 102246 127190 102298
rect 127242 102246 127254 102298
rect 127306 102246 127318 102298
rect 127370 102246 157846 102298
rect 157898 102246 157910 102298
rect 157962 102246 157974 102298
rect 158026 102246 158038 102298
rect 158090 102246 178848 102298
rect 1104 102224 178848 102246
rect 1104 101754 178848 101776
rect 1104 101702 19606 101754
rect 19658 101702 19670 101754
rect 19722 101702 19734 101754
rect 19786 101702 19798 101754
rect 19850 101702 50326 101754
rect 50378 101702 50390 101754
rect 50442 101702 50454 101754
rect 50506 101702 50518 101754
rect 50570 101702 81046 101754
rect 81098 101702 81110 101754
rect 81162 101702 81174 101754
rect 81226 101702 81238 101754
rect 81290 101702 111766 101754
rect 111818 101702 111830 101754
rect 111882 101702 111894 101754
rect 111946 101702 111958 101754
rect 112010 101702 142486 101754
rect 142538 101702 142550 101754
rect 142602 101702 142614 101754
rect 142666 101702 142678 101754
rect 142730 101702 173206 101754
rect 173258 101702 173270 101754
rect 173322 101702 173334 101754
rect 173386 101702 173398 101754
rect 173450 101702 178848 101754
rect 1104 101680 178848 101702
rect 1104 101210 178848 101232
rect 1104 101158 4246 101210
rect 4298 101158 4310 101210
rect 4362 101158 4374 101210
rect 4426 101158 4438 101210
rect 4490 101158 34966 101210
rect 35018 101158 35030 101210
rect 35082 101158 35094 101210
rect 35146 101158 35158 101210
rect 35210 101158 65686 101210
rect 65738 101158 65750 101210
rect 65802 101158 65814 101210
rect 65866 101158 65878 101210
rect 65930 101158 96406 101210
rect 96458 101158 96470 101210
rect 96522 101158 96534 101210
rect 96586 101158 96598 101210
rect 96650 101158 127126 101210
rect 127178 101158 127190 101210
rect 127242 101158 127254 101210
rect 127306 101158 127318 101210
rect 127370 101158 157846 101210
rect 157898 101158 157910 101210
rect 157962 101158 157974 101210
rect 158026 101158 158038 101210
rect 158090 101158 178848 101210
rect 1104 101136 178848 101158
rect 1104 100666 178848 100688
rect 1104 100614 19606 100666
rect 19658 100614 19670 100666
rect 19722 100614 19734 100666
rect 19786 100614 19798 100666
rect 19850 100614 50326 100666
rect 50378 100614 50390 100666
rect 50442 100614 50454 100666
rect 50506 100614 50518 100666
rect 50570 100614 81046 100666
rect 81098 100614 81110 100666
rect 81162 100614 81174 100666
rect 81226 100614 81238 100666
rect 81290 100614 111766 100666
rect 111818 100614 111830 100666
rect 111882 100614 111894 100666
rect 111946 100614 111958 100666
rect 112010 100614 142486 100666
rect 142538 100614 142550 100666
rect 142602 100614 142614 100666
rect 142666 100614 142678 100666
rect 142730 100614 173206 100666
rect 173258 100614 173270 100666
rect 173322 100614 173334 100666
rect 173386 100614 173398 100666
rect 173450 100614 178848 100666
rect 1104 100592 178848 100614
rect 1104 100122 178848 100144
rect 1104 100070 4246 100122
rect 4298 100070 4310 100122
rect 4362 100070 4374 100122
rect 4426 100070 4438 100122
rect 4490 100070 34966 100122
rect 35018 100070 35030 100122
rect 35082 100070 35094 100122
rect 35146 100070 35158 100122
rect 35210 100070 65686 100122
rect 65738 100070 65750 100122
rect 65802 100070 65814 100122
rect 65866 100070 65878 100122
rect 65930 100070 96406 100122
rect 96458 100070 96470 100122
rect 96522 100070 96534 100122
rect 96586 100070 96598 100122
rect 96650 100070 127126 100122
rect 127178 100070 127190 100122
rect 127242 100070 127254 100122
rect 127306 100070 127318 100122
rect 127370 100070 157846 100122
rect 157898 100070 157910 100122
rect 157962 100070 157974 100122
rect 158026 100070 158038 100122
rect 158090 100070 178848 100122
rect 1104 100048 178848 100070
rect 1104 99578 178848 99600
rect 1104 99526 19606 99578
rect 19658 99526 19670 99578
rect 19722 99526 19734 99578
rect 19786 99526 19798 99578
rect 19850 99526 50326 99578
rect 50378 99526 50390 99578
rect 50442 99526 50454 99578
rect 50506 99526 50518 99578
rect 50570 99526 81046 99578
rect 81098 99526 81110 99578
rect 81162 99526 81174 99578
rect 81226 99526 81238 99578
rect 81290 99526 111766 99578
rect 111818 99526 111830 99578
rect 111882 99526 111894 99578
rect 111946 99526 111958 99578
rect 112010 99526 142486 99578
rect 142538 99526 142550 99578
rect 142602 99526 142614 99578
rect 142666 99526 142678 99578
rect 142730 99526 173206 99578
rect 173258 99526 173270 99578
rect 173322 99526 173334 99578
rect 173386 99526 173398 99578
rect 173450 99526 178848 99578
rect 1104 99504 178848 99526
rect 1104 99034 178848 99056
rect 1104 98982 4246 99034
rect 4298 98982 4310 99034
rect 4362 98982 4374 99034
rect 4426 98982 4438 99034
rect 4490 98982 34966 99034
rect 35018 98982 35030 99034
rect 35082 98982 35094 99034
rect 35146 98982 35158 99034
rect 35210 98982 65686 99034
rect 65738 98982 65750 99034
rect 65802 98982 65814 99034
rect 65866 98982 65878 99034
rect 65930 98982 96406 99034
rect 96458 98982 96470 99034
rect 96522 98982 96534 99034
rect 96586 98982 96598 99034
rect 96650 98982 127126 99034
rect 127178 98982 127190 99034
rect 127242 98982 127254 99034
rect 127306 98982 127318 99034
rect 127370 98982 157846 99034
rect 157898 98982 157910 99034
rect 157962 98982 157974 99034
rect 158026 98982 158038 99034
rect 158090 98982 178848 99034
rect 1104 98960 178848 98982
rect 1104 98490 178848 98512
rect 1104 98438 19606 98490
rect 19658 98438 19670 98490
rect 19722 98438 19734 98490
rect 19786 98438 19798 98490
rect 19850 98438 50326 98490
rect 50378 98438 50390 98490
rect 50442 98438 50454 98490
rect 50506 98438 50518 98490
rect 50570 98438 81046 98490
rect 81098 98438 81110 98490
rect 81162 98438 81174 98490
rect 81226 98438 81238 98490
rect 81290 98438 111766 98490
rect 111818 98438 111830 98490
rect 111882 98438 111894 98490
rect 111946 98438 111958 98490
rect 112010 98438 142486 98490
rect 142538 98438 142550 98490
rect 142602 98438 142614 98490
rect 142666 98438 142678 98490
rect 142730 98438 173206 98490
rect 173258 98438 173270 98490
rect 173322 98438 173334 98490
rect 173386 98438 173398 98490
rect 173450 98438 178848 98490
rect 1104 98416 178848 98438
rect 1104 97946 178848 97968
rect 1104 97894 4246 97946
rect 4298 97894 4310 97946
rect 4362 97894 4374 97946
rect 4426 97894 4438 97946
rect 4490 97894 34966 97946
rect 35018 97894 35030 97946
rect 35082 97894 35094 97946
rect 35146 97894 35158 97946
rect 35210 97894 65686 97946
rect 65738 97894 65750 97946
rect 65802 97894 65814 97946
rect 65866 97894 65878 97946
rect 65930 97894 96406 97946
rect 96458 97894 96470 97946
rect 96522 97894 96534 97946
rect 96586 97894 96598 97946
rect 96650 97894 127126 97946
rect 127178 97894 127190 97946
rect 127242 97894 127254 97946
rect 127306 97894 127318 97946
rect 127370 97894 157846 97946
rect 157898 97894 157910 97946
rect 157962 97894 157974 97946
rect 158026 97894 158038 97946
rect 158090 97894 178848 97946
rect 1104 97872 178848 97894
rect 1104 97402 178848 97424
rect 1104 97350 19606 97402
rect 19658 97350 19670 97402
rect 19722 97350 19734 97402
rect 19786 97350 19798 97402
rect 19850 97350 50326 97402
rect 50378 97350 50390 97402
rect 50442 97350 50454 97402
rect 50506 97350 50518 97402
rect 50570 97350 81046 97402
rect 81098 97350 81110 97402
rect 81162 97350 81174 97402
rect 81226 97350 81238 97402
rect 81290 97350 111766 97402
rect 111818 97350 111830 97402
rect 111882 97350 111894 97402
rect 111946 97350 111958 97402
rect 112010 97350 142486 97402
rect 142538 97350 142550 97402
rect 142602 97350 142614 97402
rect 142666 97350 142678 97402
rect 142730 97350 173206 97402
rect 173258 97350 173270 97402
rect 173322 97350 173334 97402
rect 173386 97350 173398 97402
rect 173450 97350 178848 97402
rect 1104 97328 178848 97350
rect 1104 96858 178848 96880
rect 1104 96806 4246 96858
rect 4298 96806 4310 96858
rect 4362 96806 4374 96858
rect 4426 96806 4438 96858
rect 4490 96806 34966 96858
rect 35018 96806 35030 96858
rect 35082 96806 35094 96858
rect 35146 96806 35158 96858
rect 35210 96806 65686 96858
rect 65738 96806 65750 96858
rect 65802 96806 65814 96858
rect 65866 96806 65878 96858
rect 65930 96806 96406 96858
rect 96458 96806 96470 96858
rect 96522 96806 96534 96858
rect 96586 96806 96598 96858
rect 96650 96806 127126 96858
rect 127178 96806 127190 96858
rect 127242 96806 127254 96858
rect 127306 96806 127318 96858
rect 127370 96806 157846 96858
rect 157898 96806 157910 96858
rect 157962 96806 157974 96858
rect 158026 96806 158038 96858
rect 158090 96806 178848 96858
rect 1104 96784 178848 96806
rect 1104 96314 178848 96336
rect 1104 96262 19606 96314
rect 19658 96262 19670 96314
rect 19722 96262 19734 96314
rect 19786 96262 19798 96314
rect 19850 96262 50326 96314
rect 50378 96262 50390 96314
rect 50442 96262 50454 96314
rect 50506 96262 50518 96314
rect 50570 96262 81046 96314
rect 81098 96262 81110 96314
rect 81162 96262 81174 96314
rect 81226 96262 81238 96314
rect 81290 96262 111766 96314
rect 111818 96262 111830 96314
rect 111882 96262 111894 96314
rect 111946 96262 111958 96314
rect 112010 96262 142486 96314
rect 142538 96262 142550 96314
rect 142602 96262 142614 96314
rect 142666 96262 142678 96314
rect 142730 96262 173206 96314
rect 173258 96262 173270 96314
rect 173322 96262 173334 96314
rect 173386 96262 173398 96314
rect 173450 96262 178848 96314
rect 1104 96240 178848 96262
rect 1104 95770 178848 95792
rect 1104 95718 4246 95770
rect 4298 95718 4310 95770
rect 4362 95718 4374 95770
rect 4426 95718 4438 95770
rect 4490 95718 34966 95770
rect 35018 95718 35030 95770
rect 35082 95718 35094 95770
rect 35146 95718 35158 95770
rect 35210 95718 65686 95770
rect 65738 95718 65750 95770
rect 65802 95718 65814 95770
rect 65866 95718 65878 95770
rect 65930 95718 96406 95770
rect 96458 95718 96470 95770
rect 96522 95718 96534 95770
rect 96586 95718 96598 95770
rect 96650 95718 127126 95770
rect 127178 95718 127190 95770
rect 127242 95718 127254 95770
rect 127306 95718 127318 95770
rect 127370 95718 157846 95770
rect 157898 95718 157910 95770
rect 157962 95718 157974 95770
rect 158026 95718 158038 95770
rect 158090 95718 178848 95770
rect 1104 95696 178848 95718
rect 1104 95226 178848 95248
rect 1104 95174 19606 95226
rect 19658 95174 19670 95226
rect 19722 95174 19734 95226
rect 19786 95174 19798 95226
rect 19850 95174 50326 95226
rect 50378 95174 50390 95226
rect 50442 95174 50454 95226
rect 50506 95174 50518 95226
rect 50570 95174 81046 95226
rect 81098 95174 81110 95226
rect 81162 95174 81174 95226
rect 81226 95174 81238 95226
rect 81290 95174 111766 95226
rect 111818 95174 111830 95226
rect 111882 95174 111894 95226
rect 111946 95174 111958 95226
rect 112010 95174 142486 95226
rect 142538 95174 142550 95226
rect 142602 95174 142614 95226
rect 142666 95174 142678 95226
rect 142730 95174 173206 95226
rect 173258 95174 173270 95226
rect 173322 95174 173334 95226
rect 173386 95174 173398 95226
rect 173450 95174 178848 95226
rect 1104 95152 178848 95174
rect 1104 94682 178848 94704
rect 1104 94630 4246 94682
rect 4298 94630 4310 94682
rect 4362 94630 4374 94682
rect 4426 94630 4438 94682
rect 4490 94630 34966 94682
rect 35018 94630 35030 94682
rect 35082 94630 35094 94682
rect 35146 94630 35158 94682
rect 35210 94630 65686 94682
rect 65738 94630 65750 94682
rect 65802 94630 65814 94682
rect 65866 94630 65878 94682
rect 65930 94630 96406 94682
rect 96458 94630 96470 94682
rect 96522 94630 96534 94682
rect 96586 94630 96598 94682
rect 96650 94630 127126 94682
rect 127178 94630 127190 94682
rect 127242 94630 127254 94682
rect 127306 94630 127318 94682
rect 127370 94630 157846 94682
rect 157898 94630 157910 94682
rect 157962 94630 157974 94682
rect 158026 94630 158038 94682
rect 158090 94630 178848 94682
rect 1104 94608 178848 94630
rect 1104 94138 178848 94160
rect 1104 94086 19606 94138
rect 19658 94086 19670 94138
rect 19722 94086 19734 94138
rect 19786 94086 19798 94138
rect 19850 94086 50326 94138
rect 50378 94086 50390 94138
rect 50442 94086 50454 94138
rect 50506 94086 50518 94138
rect 50570 94086 81046 94138
rect 81098 94086 81110 94138
rect 81162 94086 81174 94138
rect 81226 94086 81238 94138
rect 81290 94086 111766 94138
rect 111818 94086 111830 94138
rect 111882 94086 111894 94138
rect 111946 94086 111958 94138
rect 112010 94086 142486 94138
rect 142538 94086 142550 94138
rect 142602 94086 142614 94138
rect 142666 94086 142678 94138
rect 142730 94086 173206 94138
rect 173258 94086 173270 94138
rect 173322 94086 173334 94138
rect 173386 94086 173398 94138
rect 173450 94086 178848 94138
rect 1104 94064 178848 94086
rect 1104 93594 178848 93616
rect 1104 93542 4246 93594
rect 4298 93542 4310 93594
rect 4362 93542 4374 93594
rect 4426 93542 4438 93594
rect 4490 93542 34966 93594
rect 35018 93542 35030 93594
rect 35082 93542 35094 93594
rect 35146 93542 35158 93594
rect 35210 93542 65686 93594
rect 65738 93542 65750 93594
rect 65802 93542 65814 93594
rect 65866 93542 65878 93594
rect 65930 93542 96406 93594
rect 96458 93542 96470 93594
rect 96522 93542 96534 93594
rect 96586 93542 96598 93594
rect 96650 93542 127126 93594
rect 127178 93542 127190 93594
rect 127242 93542 127254 93594
rect 127306 93542 127318 93594
rect 127370 93542 157846 93594
rect 157898 93542 157910 93594
rect 157962 93542 157974 93594
rect 158026 93542 158038 93594
rect 158090 93542 178848 93594
rect 1104 93520 178848 93542
rect 1104 93050 178848 93072
rect 1104 92998 19606 93050
rect 19658 92998 19670 93050
rect 19722 92998 19734 93050
rect 19786 92998 19798 93050
rect 19850 92998 50326 93050
rect 50378 92998 50390 93050
rect 50442 92998 50454 93050
rect 50506 92998 50518 93050
rect 50570 92998 81046 93050
rect 81098 92998 81110 93050
rect 81162 92998 81174 93050
rect 81226 92998 81238 93050
rect 81290 92998 111766 93050
rect 111818 92998 111830 93050
rect 111882 92998 111894 93050
rect 111946 92998 111958 93050
rect 112010 92998 142486 93050
rect 142538 92998 142550 93050
rect 142602 92998 142614 93050
rect 142666 92998 142678 93050
rect 142730 92998 173206 93050
rect 173258 92998 173270 93050
rect 173322 92998 173334 93050
rect 173386 92998 173398 93050
rect 173450 92998 178848 93050
rect 1104 92976 178848 92998
rect 1104 92506 178848 92528
rect 1104 92454 4246 92506
rect 4298 92454 4310 92506
rect 4362 92454 4374 92506
rect 4426 92454 4438 92506
rect 4490 92454 34966 92506
rect 35018 92454 35030 92506
rect 35082 92454 35094 92506
rect 35146 92454 35158 92506
rect 35210 92454 65686 92506
rect 65738 92454 65750 92506
rect 65802 92454 65814 92506
rect 65866 92454 65878 92506
rect 65930 92454 96406 92506
rect 96458 92454 96470 92506
rect 96522 92454 96534 92506
rect 96586 92454 96598 92506
rect 96650 92454 127126 92506
rect 127178 92454 127190 92506
rect 127242 92454 127254 92506
rect 127306 92454 127318 92506
rect 127370 92454 157846 92506
rect 157898 92454 157910 92506
rect 157962 92454 157974 92506
rect 158026 92454 158038 92506
rect 158090 92454 178848 92506
rect 1104 92432 178848 92454
rect 1104 91962 178848 91984
rect 1104 91910 19606 91962
rect 19658 91910 19670 91962
rect 19722 91910 19734 91962
rect 19786 91910 19798 91962
rect 19850 91910 50326 91962
rect 50378 91910 50390 91962
rect 50442 91910 50454 91962
rect 50506 91910 50518 91962
rect 50570 91910 81046 91962
rect 81098 91910 81110 91962
rect 81162 91910 81174 91962
rect 81226 91910 81238 91962
rect 81290 91910 111766 91962
rect 111818 91910 111830 91962
rect 111882 91910 111894 91962
rect 111946 91910 111958 91962
rect 112010 91910 142486 91962
rect 142538 91910 142550 91962
rect 142602 91910 142614 91962
rect 142666 91910 142678 91962
rect 142730 91910 173206 91962
rect 173258 91910 173270 91962
rect 173322 91910 173334 91962
rect 173386 91910 173398 91962
rect 173450 91910 178848 91962
rect 1104 91888 178848 91910
rect 1104 91418 178848 91440
rect 1104 91366 4246 91418
rect 4298 91366 4310 91418
rect 4362 91366 4374 91418
rect 4426 91366 4438 91418
rect 4490 91366 34966 91418
rect 35018 91366 35030 91418
rect 35082 91366 35094 91418
rect 35146 91366 35158 91418
rect 35210 91366 65686 91418
rect 65738 91366 65750 91418
rect 65802 91366 65814 91418
rect 65866 91366 65878 91418
rect 65930 91366 96406 91418
rect 96458 91366 96470 91418
rect 96522 91366 96534 91418
rect 96586 91366 96598 91418
rect 96650 91366 127126 91418
rect 127178 91366 127190 91418
rect 127242 91366 127254 91418
rect 127306 91366 127318 91418
rect 127370 91366 157846 91418
rect 157898 91366 157910 91418
rect 157962 91366 157974 91418
rect 158026 91366 158038 91418
rect 158090 91366 178848 91418
rect 1104 91344 178848 91366
rect 1104 90874 178848 90896
rect 1104 90822 19606 90874
rect 19658 90822 19670 90874
rect 19722 90822 19734 90874
rect 19786 90822 19798 90874
rect 19850 90822 50326 90874
rect 50378 90822 50390 90874
rect 50442 90822 50454 90874
rect 50506 90822 50518 90874
rect 50570 90822 81046 90874
rect 81098 90822 81110 90874
rect 81162 90822 81174 90874
rect 81226 90822 81238 90874
rect 81290 90822 111766 90874
rect 111818 90822 111830 90874
rect 111882 90822 111894 90874
rect 111946 90822 111958 90874
rect 112010 90822 142486 90874
rect 142538 90822 142550 90874
rect 142602 90822 142614 90874
rect 142666 90822 142678 90874
rect 142730 90822 173206 90874
rect 173258 90822 173270 90874
rect 173322 90822 173334 90874
rect 173386 90822 173398 90874
rect 173450 90822 178848 90874
rect 1104 90800 178848 90822
rect 1104 90330 178848 90352
rect 1104 90278 4246 90330
rect 4298 90278 4310 90330
rect 4362 90278 4374 90330
rect 4426 90278 4438 90330
rect 4490 90278 34966 90330
rect 35018 90278 35030 90330
rect 35082 90278 35094 90330
rect 35146 90278 35158 90330
rect 35210 90278 65686 90330
rect 65738 90278 65750 90330
rect 65802 90278 65814 90330
rect 65866 90278 65878 90330
rect 65930 90278 96406 90330
rect 96458 90278 96470 90330
rect 96522 90278 96534 90330
rect 96586 90278 96598 90330
rect 96650 90278 127126 90330
rect 127178 90278 127190 90330
rect 127242 90278 127254 90330
rect 127306 90278 127318 90330
rect 127370 90278 157846 90330
rect 157898 90278 157910 90330
rect 157962 90278 157974 90330
rect 158026 90278 158038 90330
rect 158090 90278 178848 90330
rect 1104 90256 178848 90278
rect 1104 89786 178848 89808
rect 1104 89734 19606 89786
rect 19658 89734 19670 89786
rect 19722 89734 19734 89786
rect 19786 89734 19798 89786
rect 19850 89734 50326 89786
rect 50378 89734 50390 89786
rect 50442 89734 50454 89786
rect 50506 89734 50518 89786
rect 50570 89734 81046 89786
rect 81098 89734 81110 89786
rect 81162 89734 81174 89786
rect 81226 89734 81238 89786
rect 81290 89734 111766 89786
rect 111818 89734 111830 89786
rect 111882 89734 111894 89786
rect 111946 89734 111958 89786
rect 112010 89734 142486 89786
rect 142538 89734 142550 89786
rect 142602 89734 142614 89786
rect 142666 89734 142678 89786
rect 142730 89734 173206 89786
rect 173258 89734 173270 89786
rect 173322 89734 173334 89786
rect 173386 89734 173398 89786
rect 173450 89734 178848 89786
rect 1104 89712 178848 89734
rect 1104 89242 178848 89264
rect 1104 89190 4246 89242
rect 4298 89190 4310 89242
rect 4362 89190 4374 89242
rect 4426 89190 4438 89242
rect 4490 89190 34966 89242
rect 35018 89190 35030 89242
rect 35082 89190 35094 89242
rect 35146 89190 35158 89242
rect 35210 89190 65686 89242
rect 65738 89190 65750 89242
rect 65802 89190 65814 89242
rect 65866 89190 65878 89242
rect 65930 89190 96406 89242
rect 96458 89190 96470 89242
rect 96522 89190 96534 89242
rect 96586 89190 96598 89242
rect 96650 89190 127126 89242
rect 127178 89190 127190 89242
rect 127242 89190 127254 89242
rect 127306 89190 127318 89242
rect 127370 89190 157846 89242
rect 157898 89190 157910 89242
rect 157962 89190 157974 89242
rect 158026 89190 158038 89242
rect 158090 89190 178848 89242
rect 1104 89168 178848 89190
rect 1104 88698 178848 88720
rect 1104 88646 19606 88698
rect 19658 88646 19670 88698
rect 19722 88646 19734 88698
rect 19786 88646 19798 88698
rect 19850 88646 50326 88698
rect 50378 88646 50390 88698
rect 50442 88646 50454 88698
rect 50506 88646 50518 88698
rect 50570 88646 81046 88698
rect 81098 88646 81110 88698
rect 81162 88646 81174 88698
rect 81226 88646 81238 88698
rect 81290 88646 111766 88698
rect 111818 88646 111830 88698
rect 111882 88646 111894 88698
rect 111946 88646 111958 88698
rect 112010 88646 142486 88698
rect 142538 88646 142550 88698
rect 142602 88646 142614 88698
rect 142666 88646 142678 88698
rect 142730 88646 173206 88698
rect 173258 88646 173270 88698
rect 173322 88646 173334 88698
rect 173386 88646 173398 88698
rect 173450 88646 178848 88698
rect 1104 88624 178848 88646
rect 1104 88154 178848 88176
rect 1104 88102 4246 88154
rect 4298 88102 4310 88154
rect 4362 88102 4374 88154
rect 4426 88102 4438 88154
rect 4490 88102 34966 88154
rect 35018 88102 35030 88154
rect 35082 88102 35094 88154
rect 35146 88102 35158 88154
rect 35210 88102 65686 88154
rect 65738 88102 65750 88154
rect 65802 88102 65814 88154
rect 65866 88102 65878 88154
rect 65930 88102 96406 88154
rect 96458 88102 96470 88154
rect 96522 88102 96534 88154
rect 96586 88102 96598 88154
rect 96650 88102 127126 88154
rect 127178 88102 127190 88154
rect 127242 88102 127254 88154
rect 127306 88102 127318 88154
rect 127370 88102 157846 88154
rect 157898 88102 157910 88154
rect 157962 88102 157974 88154
rect 158026 88102 158038 88154
rect 158090 88102 178848 88154
rect 1104 88080 178848 88102
rect 1104 87610 178848 87632
rect 1104 87558 19606 87610
rect 19658 87558 19670 87610
rect 19722 87558 19734 87610
rect 19786 87558 19798 87610
rect 19850 87558 50326 87610
rect 50378 87558 50390 87610
rect 50442 87558 50454 87610
rect 50506 87558 50518 87610
rect 50570 87558 81046 87610
rect 81098 87558 81110 87610
rect 81162 87558 81174 87610
rect 81226 87558 81238 87610
rect 81290 87558 111766 87610
rect 111818 87558 111830 87610
rect 111882 87558 111894 87610
rect 111946 87558 111958 87610
rect 112010 87558 142486 87610
rect 142538 87558 142550 87610
rect 142602 87558 142614 87610
rect 142666 87558 142678 87610
rect 142730 87558 173206 87610
rect 173258 87558 173270 87610
rect 173322 87558 173334 87610
rect 173386 87558 173398 87610
rect 173450 87558 178848 87610
rect 1104 87536 178848 87558
rect 1104 87066 178848 87088
rect 1104 87014 4246 87066
rect 4298 87014 4310 87066
rect 4362 87014 4374 87066
rect 4426 87014 4438 87066
rect 4490 87014 34966 87066
rect 35018 87014 35030 87066
rect 35082 87014 35094 87066
rect 35146 87014 35158 87066
rect 35210 87014 65686 87066
rect 65738 87014 65750 87066
rect 65802 87014 65814 87066
rect 65866 87014 65878 87066
rect 65930 87014 96406 87066
rect 96458 87014 96470 87066
rect 96522 87014 96534 87066
rect 96586 87014 96598 87066
rect 96650 87014 127126 87066
rect 127178 87014 127190 87066
rect 127242 87014 127254 87066
rect 127306 87014 127318 87066
rect 127370 87014 157846 87066
rect 157898 87014 157910 87066
rect 157962 87014 157974 87066
rect 158026 87014 158038 87066
rect 158090 87014 178848 87066
rect 1104 86992 178848 87014
rect 1104 86522 178848 86544
rect 1104 86470 19606 86522
rect 19658 86470 19670 86522
rect 19722 86470 19734 86522
rect 19786 86470 19798 86522
rect 19850 86470 50326 86522
rect 50378 86470 50390 86522
rect 50442 86470 50454 86522
rect 50506 86470 50518 86522
rect 50570 86470 81046 86522
rect 81098 86470 81110 86522
rect 81162 86470 81174 86522
rect 81226 86470 81238 86522
rect 81290 86470 111766 86522
rect 111818 86470 111830 86522
rect 111882 86470 111894 86522
rect 111946 86470 111958 86522
rect 112010 86470 142486 86522
rect 142538 86470 142550 86522
rect 142602 86470 142614 86522
rect 142666 86470 142678 86522
rect 142730 86470 173206 86522
rect 173258 86470 173270 86522
rect 173322 86470 173334 86522
rect 173386 86470 173398 86522
rect 173450 86470 178848 86522
rect 1104 86448 178848 86470
rect 1104 85978 178848 86000
rect 1104 85926 4246 85978
rect 4298 85926 4310 85978
rect 4362 85926 4374 85978
rect 4426 85926 4438 85978
rect 4490 85926 34966 85978
rect 35018 85926 35030 85978
rect 35082 85926 35094 85978
rect 35146 85926 35158 85978
rect 35210 85926 65686 85978
rect 65738 85926 65750 85978
rect 65802 85926 65814 85978
rect 65866 85926 65878 85978
rect 65930 85926 96406 85978
rect 96458 85926 96470 85978
rect 96522 85926 96534 85978
rect 96586 85926 96598 85978
rect 96650 85926 127126 85978
rect 127178 85926 127190 85978
rect 127242 85926 127254 85978
rect 127306 85926 127318 85978
rect 127370 85926 157846 85978
rect 157898 85926 157910 85978
rect 157962 85926 157974 85978
rect 158026 85926 158038 85978
rect 158090 85926 178848 85978
rect 1104 85904 178848 85926
rect 1104 85434 178848 85456
rect 1104 85382 19606 85434
rect 19658 85382 19670 85434
rect 19722 85382 19734 85434
rect 19786 85382 19798 85434
rect 19850 85382 50326 85434
rect 50378 85382 50390 85434
rect 50442 85382 50454 85434
rect 50506 85382 50518 85434
rect 50570 85382 81046 85434
rect 81098 85382 81110 85434
rect 81162 85382 81174 85434
rect 81226 85382 81238 85434
rect 81290 85382 111766 85434
rect 111818 85382 111830 85434
rect 111882 85382 111894 85434
rect 111946 85382 111958 85434
rect 112010 85382 142486 85434
rect 142538 85382 142550 85434
rect 142602 85382 142614 85434
rect 142666 85382 142678 85434
rect 142730 85382 173206 85434
rect 173258 85382 173270 85434
rect 173322 85382 173334 85434
rect 173386 85382 173398 85434
rect 173450 85382 178848 85434
rect 1104 85360 178848 85382
rect 1104 84890 178848 84912
rect 1104 84838 4246 84890
rect 4298 84838 4310 84890
rect 4362 84838 4374 84890
rect 4426 84838 4438 84890
rect 4490 84838 34966 84890
rect 35018 84838 35030 84890
rect 35082 84838 35094 84890
rect 35146 84838 35158 84890
rect 35210 84838 65686 84890
rect 65738 84838 65750 84890
rect 65802 84838 65814 84890
rect 65866 84838 65878 84890
rect 65930 84838 96406 84890
rect 96458 84838 96470 84890
rect 96522 84838 96534 84890
rect 96586 84838 96598 84890
rect 96650 84838 127126 84890
rect 127178 84838 127190 84890
rect 127242 84838 127254 84890
rect 127306 84838 127318 84890
rect 127370 84838 157846 84890
rect 157898 84838 157910 84890
rect 157962 84838 157974 84890
rect 158026 84838 158038 84890
rect 158090 84838 178848 84890
rect 1104 84816 178848 84838
rect 1104 84346 178848 84368
rect 1104 84294 19606 84346
rect 19658 84294 19670 84346
rect 19722 84294 19734 84346
rect 19786 84294 19798 84346
rect 19850 84294 50326 84346
rect 50378 84294 50390 84346
rect 50442 84294 50454 84346
rect 50506 84294 50518 84346
rect 50570 84294 81046 84346
rect 81098 84294 81110 84346
rect 81162 84294 81174 84346
rect 81226 84294 81238 84346
rect 81290 84294 111766 84346
rect 111818 84294 111830 84346
rect 111882 84294 111894 84346
rect 111946 84294 111958 84346
rect 112010 84294 142486 84346
rect 142538 84294 142550 84346
rect 142602 84294 142614 84346
rect 142666 84294 142678 84346
rect 142730 84294 173206 84346
rect 173258 84294 173270 84346
rect 173322 84294 173334 84346
rect 173386 84294 173398 84346
rect 173450 84294 178848 84346
rect 1104 84272 178848 84294
rect 1104 83802 178848 83824
rect 1104 83750 4246 83802
rect 4298 83750 4310 83802
rect 4362 83750 4374 83802
rect 4426 83750 4438 83802
rect 4490 83750 34966 83802
rect 35018 83750 35030 83802
rect 35082 83750 35094 83802
rect 35146 83750 35158 83802
rect 35210 83750 65686 83802
rect 65738 83750 65750 83802
rect 65802 83750 65814 83802
rect 65866 83750 65878 83802
rect 65930 83750 96406 83802
rect 96458 83750 96470 83802
rect 96522 83750 96534 83802
rect 96586 83750 96598 83802
rect 96650 83750 127126 83802
rect 127178 83750 127190 83802
rect 127242 83750 127254 83802
rect 127306 83750 127318 83802
rect 127370 83750 157846 83802
rect 157898 83750 157910 83802
rect 157962 83750 157974 83802
rect 158026 83750 158038 83802
rect 158090 83750 178848 83802
rect 1104 83728 178848 83750
rect 1104 83258 178848 83280
rect 1104 83206 19606 83258
rect 19658 83206 19670 83258
rect 19722 83206 19734 83258
rect 19786 83206 19798 83258
rect 19850 83206 50326 83258
rect 50378 83206 50390 83258
rect 50442 83206 50454 83258
rect 50506 83206 50518 83258
rect 50570 83206 81046 83258
rect 81098 83206 81110 83258
rect 81162 83206 81174 83258
rect 81226 83206 81238 83258
rect 81290 83206 111766 83258
rect 111818 83206 111830 83258
rect 111882 83206 111894 83258
rect 111946 83206 111958 83258
rect 112010 83206 142486 83258
rect 142538 83206 142550 83258
rect 142602 83206 142614 83258
rect 142666 83206 142678 83258
rect 142730 83206 173206 83258
rect 173258 83206 173270 83258
rect 173322 83206 173334 83258
rect 173386 83206 173398 83258
rect 173450 83206 178848 83258
rect 1104 83184 178848 83206
rect 1104 82714 178848 82736
rect 1104 82662 4246 82714
rect 4298 82662 4310 82714
rect 4362 82662 4374 82714
rect 4426 82662 4438 82714
rect 4490 82662 34966 82714
rect 35018 82662 35030 82714
rect 35082 82662 35094 82714
rect 35146 82662 35158 82714
rect 35210 82662 65686 82714
rect 65738 82662 65750 82714
rect 65802 82662 65814 82714
rect 65866 82662 65878 82714
rect 65930 82662 96406 82714
rect 96458 82662 96470 82714
rect 96522 82662 96534 82714
rect 96586 82662 96598 82714
rect 96650 82662 127126 82714
rect 127178 82662 127190 82714
rect 127242 82662 127254 82714
rect 127306 82662 127318 82714
rect 127370 82662 157846 82714
rect 157898 82662 157910 82714
rect 157962 82662 157974 82714
rect 158026 82662 158038 82714
rect 158090 82662 178848 82714
rect 1104 82640 178848 82662
rect 1104 82170 178848 82192
rect 1104 82118 19606 82170
rect 19658 82118 19670 82170
rect 19722 82118 19734 82170
rect 19786 82118 19798 82170
rect 19850 82118 50326 82170
rect 50378 82118 50390 82170
rect 50442 82118 50454 82170
rect 50506 82118 50518 82170
rect 50570 82118 81046 82170
rect 81098 82118 81110 82170
rect 81162 82118 81174 82170
rect 81226 82118 81238 82170
rect 81290 82118 111766 82170
rect 111818 82118 111830 82170
rect 111882 82118 111894 82170
rect 111946 82118 111958 82170
rect 112010 82118 142486 82170
rect 142538 82118 142550 82170
rect 142602 82118 142614 82170
rect 142666 82118 142678 82170
rect 142730 82118 173206 82170
rect 173258 82118 173270 82170
rect 173322 82118 173334 82170
rect 173386 82118 173398 82170
rect 173450 82118 178848 82170
rect 1104 82096 178848 82118
rect 1104 81626 178848 81648
rect 1104 81574 4246 81626
rect 4298 81574 4310 81626
rect 4362 81574 4374 81626
rect 4426 81574 4438 81626
rect 4490 81574 34966 81626
rect 35018 81574 35030 81626
rect 35082 81574 35094 81626
rect 35146 81574 35158 81626
rect 35210 81574 65686 81626
rect 65738 81574 65750 81626
rect 65802 81574 65814 81626
rect 65866 81574 65878 81626
rect 65930 81574 96406 81626
rect 96458 81574 96470 81626
rect 96522 81574 96534 81626
rect 96586 81574 96598 81626
rect 96650 81574 127126 81626
rect 127178 81574 127190 81626
rect 127242 81574 127254 81626
rect 127306 81574 127318 81626
rect 127370 81574 157846 81626
rect 157898 81574 157910 81626
rect 157962 81574 157974 81626
rect 158026 81574 158038 81626
rect 158090 81574 178848 81626
rect 1104 81552 178848 81574
rect 1104 81082 178848 81104
rect 1104 81030 19606 81082
rect 19658 81030 19670 81082
rect 19722 81030 19734 81082
rect 19786 81030 19798 81082
rect 19850 81030 50326 81082
rect 50378 81030 50390 81082
rect 50442 81030 50454 81082
rect 50506 81030 50518 81082
rect 50570 81030 81046 81082
rect 81098 81030 81110 81082
rect 81162 81030 81174 81082
rect 81226 81030 81238 81082
rect 81290 81030 111766 81082
rect 111818 81030 111830 81082
rect 111882 81030 111894 81082
rect 111946 81030 111958 81082
rect 112010 81030 142486 81082
rect 142538 81030 142550 81082
rect 142602 81030 142614 81082
rect 142666 81030 142678 81082
rect 142730 81030 173206 81082
rect 173258 81030 173270 81082
rect 173322 81030 173334 81082
rect 173386 81030 173398 81082
rect 173450 81030 178848 81082
rect 1104 81008 178848 81030
rect 1104 80538 178848 80560
rect 1104 80486 4246 80538
rect 4298 80486 4310 80538
rect 4362 80486 4374 80538
rect 4426 80486 4438 80538
rect 4490 80486 34966 80538
rect 35018 80486 35030 80538
rect 35082 80486 35094 80538
rect 35146 80486 35158 80538
rect 35210 80486 65686 80538
rect 65738 80486 65750 80538
rect 65802 80486 65814 80538
rect 65866 80486 65878 80538
rect 65930 80486 96406 80538
rect 96458 80486 96470 80538
rect 96522 80486 96534 80538
rect 96586 80486 96598 80538
rect 96650 80486 127126 80538
rect 127178 80486 127190 80538
rect 127242 80486 127254 80538
rect 127306 80486 127318 80538
rect 127370 80486 157846 80538
rect 157898 80486 157910 80538
rect 157962 80486 157974 80538
rect 158026 80486 158038 80538
rect 158090 80486 178848 80538
rect 1104 80464 178848 80486
rect 1104 79994 178848 80016
rect 1104 79942 19606 79994
rect 19658 79942 19670 79994
rect 19722 79942 19734 79994
rect 19786 79942 19798 79994
rect 19850 79942 50326 79994
rect 50378 79942 50390 79994
rect 50442 79942 50454 79994
rect 50506 79942 50518 79994
rect 50570 79942 81046 79994
rect 81098 79942 81110 79994
rect 81162 79942 81174 79994
rect 81226 79942 81238 79994
rect 81290 79942 111766 79994
rect 111818 79942 111830 79994
rect 111882 79942 111894 79994
rect 111946 79942 111958 79994
rect 112010 79942 142486 79994
rect 142538 79942 142550 79994
rect 142602 79942 142614 79994
rect 142666 79942 142678 79994
rect 142730 79942 173206 79994
rect 173258 79942 173270 79994
rect 173322 79942 173334 79994
rect 173386 79942 173398 79994
rect 173450 79942 178848 79994
rect 1104 79920 178848 79942
rect 1104 79450 178848 79472
rect 1104 79398 4246 79450
rect 4298 79398 4310 79450
rect 4362 79398 4374 79450
rect 4426 79398 4438 79450
rect 4490 79398 34966 79450
rect 35018 79398 35030 79450
rect 35082 79398 35094 79450
rect 35146 79398 35158 79450
rect 35210 79398 65686 79450
rect 65738 79398 65750 79450
rect 65802 79398 65814 79450
rect 65866 79398 65878 79450
rect 65930 79398 96406 79450
rect 96458 79398 96470 79450
rect 96522 79398 96534 79450
rect 96586 79398 96598 79450
rect 96650 79398 127126 79450
rect 127178 79398 127190 79450
rect 127242 79398 127254 79450
rect 127306 79398 127318 79450
rect 127370 79398 157846 79450
rect 157898 79398 157910 79450
rect 157962 79398 157974 79450
rect 158026 79398 158038 79450
rect 158090 79398 178848 79450
rect 1104 79376 178848 79398
rect 1104 78906 178848 78928
rect 1104 78854 19606 78906
rect 19658 78854 19670 78906
rect 19722 78854 19734 78906
rect 19786 78854 19798 78906
rect 19850 78854 50326 78906
rect 50378 78854 50390 78906
rect 50442 78854 50454 78906
rect 50506 78854 50518 78906
rect 50570 78854 81046 78906
rect 81098 78854 81110 78906
rect 81162 78854 81174 78906
rect 81226 78854 81238 78906
rect 81290 78854 111766 78906
rect 111818 78854 111830 78906
rect 111882 78854 111894 78906
rect 111946 78854 111958 78906
rect 112010 78854 142486 78906
rect 142538 78854 142550 78906
rect 142602 78854 142614 78906
rect 142666 78854 142678 78906
rect 142730 78854 173206 78906
rect 173258 78854 173270 78906
rect 173322 78854 173334 78906
rect 173386 78854 173398 78906
rect 173450 78854 178848 78906
rect 1104 78832 178848 78854
rect 1104 78362 178848 78384
rect 1104 78310 4246 78362
rect 4298 78310 4310 78362
rect 4362 78310 4374 78362
rect 4426 78310 4438 78362
rect 4490 78310 34966 78362
rect 35018 78310 35030 78362
rect 35082 78310 35094 78362
rect 35146 78310 35158 78362
rect 35210 78310 65686 78362
rect 65738 78310 65750 78362
rect 65802 78310 65814 78362
rect 65866 78310 65878 78362
rect 65930 78310 96406 78362
rect 96458 78310 96470 78362
rect 96522 78310 96534 78362
rect 96586 78310 96598 78362
rect 96650 78310 127126 78362
rect 127178 78310 127190 78362
rect 127242 78310 127254 78362
rect 127306 78310 127318 78362
rect 127370 78310 157846 78362
rect 157898 78310 157910 78362
rect 157962 78310 157974 78362
rect 158026 78310 158038 78362
rect 158090 78310 178848 78362
rect 1104 78288 178848 78310
rect 1104 77818 178848 77840
rect 1104 77766 19606 77818
rect 19658 77766 19670 77818
rect 19722 77766 19734 77818
rect 19786 77766 19798 77818
rect 19850 77766 50326 77818
rect 50378 77766 50390 77818
rect 50442 77766 50454 77818
rect 50506 77766 50518 77818
rect 50570 77766 81046 77818
rect 81098 77766 81110 77818
rect 81162 77766 81174 77818
rect 81226 77766 81238 77818
rect 81290 77766 111766 77818
rect 111818 77766 111830 77818
rect 111882 77766 111894 77818
rect 111946 77766 111958 77818
rect 112010 77766 142486 77818
rect 142538 77766 142550 77818
rect 142602 77766 142614 77818
rect 142666 77766 142678 77818
rect 142730 77766 173206 77818
rect 173258 77766 173270 77818
rect 173322 77766 173334 77818
rect 173386 77766 173398 77818
rect 173450 77766 178848 77818
rect 1104 77744 178848 77766
rect 1104 77274 178848 77296
rect 1104 77222 4246 77274
rect 4298 77222 4310 77274
rect 4362 77222 4374 77274
rect 4426 77222 4438 77274
rect 4490 77222 34966 77274
rect 35018 77222 35030 77274
rect 35082 77222 35094 77274
rect 35146 77222 35158 77274
rect 35210 77222 65686 77274
rect 65738 77222 65750 77274
rect 65802 77222 65814 77274
rect 65866 77222 65878 77274
rect 65930 77222 96406 77274
rect 96458 77222 96470 77274
rect 96522 77222 96534 77274
rect 96586 77222 96598 77274
rect 96650 77222 127126 77274
rect 127178 77222 127190 77274
rect 127242 77222 127254 77274
rect 127306 77222 127318 77274
rect 127370 77222 157846 77274
rect 157898 77222 157910 77274
rect 157962 77222 157974 77274
rect 158026 77222 158038 77274
rect 158090 77222 178848 77274
rect 1104 77200 178848 77222
rect 1104 76730 178848 76752
rect 1104 76678 19606 76730
rect 19658 76678 19670 76730
rect 19722 76678 19734 76730
rect 19786 76678 19798 76730
rect 19850 76678 50326 76730
rect 50378 76678 50390 76730
rect 50442 76678 50454 76730
rect 50506 76678 50518 76730
rect 50570 76678 81046 76730
rect 81098 76678 81110 76730
rect 81162 76678 81174 76730
rect 81226 76678 81238 76730
rect 81290 76678 111766 76730
rect 111818 76678 111830 76730
rect 111882 76678 111894 76730
rect 111946 76678 111958 76730
rect 112010 76678 142486 76730
rect 142538 76678 142550 76730
rect 142602 76678 142614 76730
rect 142666 76678 142678 76730
rect 142730 76678 173206 76730
rect 173258 76678 173270 76730
rect 173322 76678 173334 76730
rect 173386 76678 173398 76730
rect 173450 76678 178848 76730
rect 1104 76656 178848 76678
rect 1104 76186 178848 76208
rect 1104 76134 4246 76186
rect 4298 76134 4310 76186
rect 4362 76134 4374 76186
rect 4426 76134 4438 76186
rect 4490 76134 34966 76186
rect 35018 76134 35030 76186
rect 35082 76134 35094 76186
rect 35146 76134 35158 76186
rect 35210 76134 65686 76186
rect 65738 76134 65750 76186
rect 65802 76134 65814 76186
rect 65866 76134 65878 76186
rect 65930 76134 96406 76186
rect 96458 76134 96470 76186
rect 96522 76134 96534 76186
rect 96586 76134 96598 76186
rect 96650 76134 127126 76186
rect 127178 76134 127190 76186
rect 127242 76134 127254 76186
rect 127306 76134 127318 76186
rect 127370 76134 157846 76186
rect 157898 76134 157910 76186
rect 157962 76134 157974 76186
rect 158026 76134 158038 76186
rect 158090 76134 178848 76186
rect 1104 76112 178848 76134
rect 1104 75642 178848 75664
rect 1104 75590 19606 75642
rect 19658 75590 19670 75642
rect 19722 75590 19734 75642
rect 19786 75590 19798 75642
rect 19850 75590 50326 75642
rect 50378 75590 50390 75642
rect 50442 75590 50454 75642
rect 50506 75590 50518 75642
rect 50570 75590 81046 75642
rect 81098 75590 81110 75642
rect 81162 75590 81174 75642
rect 81226 75590 81238 75642
rect 81290 75590 111766 75642
rect 111818 75590 111830 75642
rect 111882 75590 111894 75642
rect 111946 75590 111958 75642
rect 112010 75590 142486 75642
rect 142538 75590 142550 75642
rect 142602 75590 142614 75642
rect 142666 75590 142678 75642
rect 142730 75590 173206 75642
rect 173258 75590 173270 75642
rect 173322 75590 173334 75642
rect 173386 75590 173398 75642
rect 173450 75590 178848 75642
rect 1104 75568 178848 75590
rect 1104 75098 178848 75120
rect 1104 75046 4246 75098
rect 4298 75046 4310 75098
rect 4362 75046 4374 75098
rect 4426 75046 4438 75098
rect 4490 75046 34966 75098
rect 35018 75046 35030 75098
rect 35082 75046 35094 75098
rect 35146 75046 35158 75098
rect 35210 75046 65686 75098
rect 65738 75046 65750 75098
rect 65802 75046 65814 75098
rect 65866 75046 65878 75098
rect 65930 75046 96406 75098
rect 96458 75046 96470 75098
rect 96522 75046 96534 75098
rect 96586 75046 96598 75098
rect 96650 75046 127126 75098
rect 127178 75046 127190 75098
rect 127242 75046 127254 75098
rect 127306 75046 127318 75098
rect 127370 75046 157846 75098
rect 157898 75046 157910 75098
rect 157962 75046 157974 75098
rect 158026 75046 158038 75098
rect 158090 75046 178848 75098
rect 1104 75024 178848 75046
rect 1104 74554 178848 74576
rect 1104 74502 19606 74554
rect 19658 74502 19670 74554
rect 19722 74502 19734 74554
rect 19786 74502 19798 74554
rect 19850 74502 50326 74554
rect 50378 74502 50390 74554
rect 50442 74502 50454 74554
rect 50506 74502 50518 74554
rect 50570 74502 81046 74554
rect 81098 74502 81110 74554
rect 81162 74502 81174 74554
rect 81226 74502 81238 74554
rect 81290 74502 111766 74554
rect 111818 74502 111830 74554
rect 111882 74502 111894 74554
rect 111946 74502 111958 74554
rect 112010 74502 142486 74554
rect 142538 74502 142550 74554
rect 142602 74502 142614 74554
rect 142666 74502 142678 74554
rect 142730 74502 173206 74554
rect 173258 74502 173270 74554
rect 173322 74502 173334 74554
rect 173386 74502 173398 74554
rect 173450 74502 178848 74554
rect 1104 74480 178848 74502
rect 1104 74010 178848 74032
rect 1104 73958 4246 74010
rect 4298 73958 4310 74010
rect 4362 73958 4374 74010
rect 4426 73958 4438 74010
rect 4490 73958 34966 74010
rect 35018 73958 35030 74010
rect 35082 73958 35094 74010
rect 35146 73958 35158 74010
rect 35210 73958 65686 74010
rect 65738 73958 65750 74010
rect 65802 73958 65814 74010
rect 65866 73958 65878 74010
rect 65930 73958 96406 74010
rect 96458 73958 96470 74010
rect 96522 73958 96534 74010
rect 96586 73958 96598 74010
rect 96650 73958 127126 74010
rect 127178 73958 127190 74010
rect 127242 73958 127254 74010
rect 127306 73958 127318 74010
rect 127370 73958 157846 74010
rect 157898 73958 157910 74010
rect 157962 73958 157974 74010
rect 158026 73958 158038 74010
rect 158090 73958 178848 74010
rect 1104 73936 178848 73958
rect 1104 73466 178848 73488
rect 1104 73414 19606 73466
rect 19658 73414 19670 73466
rect 19722 73414 19734 73466
rect 19786 73414 19798 73466
rect 19850 73414 50326 73466
rect 50378 73414 50390 73466
rect 50442 73414 50454 73466
rect 50506 73414 50518 73466
rect 50570 73414 81046 73466
rect 81098 73414 81110 73466
rect 81162 73414 81174 73466
rect 81226 73414 81238 73466
rect 81290 73414 111766 73466
rect 111818 73414 111830 73466
rect 111882 73414 111894 73466
rect 111946 73414 111958 73466
rect 112010 73414 142486 73466
rect 142538 73414 142550 73466
rect 142602 73414 142614 73466
rect 142666 73414 142678 73466
rect 142730 73414 173206 73466
rect 173258 73414 173270 73466
rect 173322 73414 173334 73466
rect 173386 73414 173398 73466
rect 173450 73414 178848 73466
rect 1104 73392 178848 73414
rect 1104 72922 178848 72944
rect 1104 72870 4246 72922
rect 4298 72870 4310 72922
rect 4362 72870 4374 72922
rect 4426 72870 4438 72922
rect 4490 72870 34966 72922
rect 35018 72870 35030 72922
rect 35082 72870 35094 72922
rect 35146 72870 35158 72922
rect 35210 72870 65686 72922
rect 65738 72870 65750 72922
rect 65802 72870 65814 72922
rect 65866 72870 65878 72922
rect 65930 72870 96406 72922
rect 96458 72870 96470 72922
rect 96522 72870 96534 72922
rect 96586 72870 96598 72922
rect 96650 72870 127126 72922
rect 127178 72870 127190 72922
rect 127242 72870 127254 72922
rect 127306 72870 127318 72922
rect 127370 72870 157846 72922
rect 157898 72870 157910 72922
rect 157962 72870 157974 72922
rect 158026 72870 158038 72922
rect 158090 72870 178848 72922
rect 1104 72848 178848 72870
rect 1104 72378 178848 72400
rect 1104 72326 19606 72378
rect 19658 72326 19670 72378
rect 19722 72326 19734 72378
rect 19786 72326 19798 72378
rect 19850 72326 50326 72378
rect 50378 72326 50390 72378
rect 50442 72326 50454 72378
rect 50506 72326 50518 72378
rect 50570 72326 81046 72378
rect 81098 72326 81110 72378
rect 81162 72326 81174 72378
rect 81226 72326 81238 72378
rect 81290 72326 111766 72378
rect 111818 72326 111830 72378
rect 111882 72326 111894 72378
rect 111946 72326 111958 72378
rect 112010 72326 142486 72378
rect 142538 72326 142550 72378
rect 142602 72326 142614 72378
rect 142666 72326 142678 72378
rect 142730 72326 173206 72378
rect 173258 72326 173270 72378
rect 173322 72326 173334 72378
rect 173386 72326 173398 72378
rect 173450 72326 178848 72378
rect 1104 72304 178848 72326
rect 1104 71834 178848 71856
rect 1104 71782 4246 71834
rect 4298 71782 4310 71834
rect 4362 71782 4374 71834
rect 4426 71782 4438 71834
rect 4490 71782 34966 71834
rect 35018 71782 35030 71834
rect 35082 71782 35094 71834
rect 35146 71782 35158 71834
rect 35210 71782 65686 71834
rect 65738 71782 65750 71834
rect 65802 71782 65814 71834
rect 65866 71782 65878 71834
rect 65930 71782 96406 71834
rect 96458 71782 96470 71834
rect 96522 71782 96534 71834
rect 96586 71782 96598 71834
rect 96650 71782 127126 71834
rect 127178 71782 127190 71834
rect 127242 71782 127254 71834
rect 127306 71782 127318 71834
rect 127370 71782 157846 71834
rect 157898 71782 157910 71834
rect 157962 71782 157974 71834
rect 158026 71782 158038 71834
rect 158090 71782 178848 71834
rect 1104 71760 178848 71782
rect 1104 71290 178848 71312
rect 1104 71238 19606 71290
rect 19658 71238 19670 71290
rect 19722 71238 19734 71290
rect 19786 71238 19798 71290
rect 19850 71238 50326 71290
rect 50378 71238 50390 71290
rect 50442 71238 50454 71290
rect 50506 71238 50518 71290
rect 50570 71238 81046 71290
rect 81098 71238 81110 71290
rect 81162 71238 81174 71290
rect 81226 71238 81238 71290
rect 81290 71238 111766 71290
rect 111818 71238 111830 71290
rect 111882 71238 111894 71290
rect 111946 71238 111958 71290
rect 112010 71238 142486 71290
rect 142538 71238 142550 71290
rect 142602 71238 142614 71290
rect 142666 71238 142678 71290
rect 142730 71238 173206 71290
rect 173258 71238 173270 71290
rect 173322 71238 173334 71290
rect 173386 71238 173398 71290
rect 173450 71238 178848 71290
rect 1104 71216 178848 71238
rect 1104 70746 178848 70768
rect 1104 70694 4246 70746
rect 4298 70694 4310 70746
rect 4362 70694 4374 70746
rect 4426 70694 4438 70746
rect 4490 70694 34966 70746
rect 35018 70694 35030 70746
rect 35082 70694 35094 70746
rect 35146 70694 35158 70746
rect 35210 70694 65686 70746
rect 65738 70694 65750 70746
rect 65802 70694 65814 70746
rect 65866 70694 65878 70746
rect 65930 70694 96406 70746
rect 96458 70694 96470 70746
rect 96522 70694 96534 70746
rect 96586 70694 96598 70746
rect 96650 70694 127126 70746
rect 127178 70694 127190 70746
rect 127242 70694 127254 70746
rect 127306 70694 127318 70746
rect 127370 70694 157846 70746
rect 157898 70694 157910 70746
rect 157962 70694 157974 70746
rect 158026 70694 158038 70746
rect 158090 70694 178848 70746
rect 1104 70672 178848 70694
rect 1104 70202 178848 70224
rect 1104 70150 19606 70202
rect 19658 70150 19670 70202
rect 19722 70150 19734 70202
rect 19786 70150 19798 70202
rect 19850 70150 50326 70202
rect 50378 70150 50390 70202
rect 50442 70150 50454 70202
rect 50506 70150 50518 70202
rect 50570 70150 81046 70202
rect 81098 70150 81110 70202
rect 81162 70150 81174 70202
rect 81226 70150 81238 70202
rect 81290 70150 111766 70202
rect 111818 70150 111830 70202
rect 111882 70150 111894 70202
rect 111946 70150 111958 70202
rect 112010 70150 142486 70202
rect 142538 70150 142550 70202
rect 142602 70150 142614 70202
rect 142666 70150 142678 70202
rect 142730 70150 173206 70202
rect 173258 70150 173270 70202
rect 173322 70150 173334 70202
rect 173386 70150 173398 70202
rect 173450 70150 178848 70202
rect 1104 70128 178848 70150
rect 1104 69658 178848 69680
rect 1104 69606 4246 69658
rect 4298 69606 4310 69658
rect 4362 69606 4374 69658
rect 4426 69606 4438 69658
rect 4490 69606 34966 69658
rect 35018 69606 35030 69658
rect 35082 69606 35094 69658
rect 35146 69606 35158 69658
rect 35210 69606 65686 69658
rect 65738 69606 65750 69658
rect 65802 69606 65814 69658
rect 65866 69606 65878 69658
rect 65930 69606 96406 69658
rect 96458 69606 96470 69658
rect 96522 69606 96534 69658
rect 96586 69606 96598 69658
rect 96650 69606 127126 69658
rect 127178 69606 127190 69658
rect 127242 69606 127254 69658
rect 127306 69606 127318 69658
rect 127370 69606 157846 69658
rect 157898 69606 157910 69658
rect 157962 69606 157974 69658
rect 158026 69606 158038 69658
rect 158090 69606 178848 69658
rect 1104 69584 178848 69606
rect 1104 69114 178848 69136
rect 1104 69062 19606 69114
rect 19658 69062 19670 69114
rect 19722 69062 19734 69114
rect 19786 69062 19798 69114
rect 19850 69062 50326 69114
rect 50378 69062 50390 69114
rect 50442 69062 50454 69114
rect 50506 69062 50518 69114
rect 50570 69062 81046 69114
rect 81098 69062 81110 69114
rect 81162 69062 81174 69114
rect 81226 69062 81238 69114
rect 81290 69062 111766 69114
rect 111818 69062 111830 69114
rect 111882 69062 111894 69114
rect 111946 69062 111958 69114
rect 112010 69062 142486 69114
rect 142538 69062 142550 69114
rect 142602 69062 142614 69114
rect 142666 69062 142678 69114
rect 142730 69062 173206 69114
rect 173258 69062 173270 69114
rect 173322 69062 173334 69114
rect 173386 69062 173398 69114
rect 173450 69062 178848 69114
rect 1104 69040 178848 69062
rect 1104 68570 178848 68592
rect 1104 68518 4246 68570
rect 4298 68518 4310 68570
rect 4362 68518 4374 68570
rect 4426 68518 4438 68570
rect 4490 68518 34966 68570
rect 35018 68518 35030 68570
rect 35082 68518 35094 68570
rect 35146 68518 35158 68570
rect 35210 68518 65686 68570
rect 65738 68518 65750 68570
rect 65802 68518 65814 68570
rect 65866 68518 65878 68570
rect 65930 68518 96406 68570
rect 96458 68518 96470 68570
rect 96522 68518 96534 68570
rect 96586 68518 96598 68570
rect 96650 68518 127126 68570
rect 127178 68518 127190 68570
rect 127242 68518 127254 68570
rect 127306 68518 127318 68570
rect 127370 68518 157846 68570
rect 157898 68518 157910 68570
rect 157962 68518 157974 68570
rect 158026 68518 158038 68570
rect 158090 68518 178848 68570
rect 1104 68496 178848 68518
rect 1104 68026 178848 68048
rect 1104 67974 19606 68026
rect 19658 67974 19670 68026
rect 19722 67974 19734 68026
rect 19786 67974 19798 68026
rect 19850 67974 50326 68026
rect 50378 67974 50390 68026
rect 50442 67974 50454 68026
rect 50506 67974 50518 68026
rect 50570 67974 81046 68026
rect 81098 67974 81110 68026
rect 81162 67974 81174 68026
rect 81226 67974 81238 68026
rect 81290 67974 111766 68026
rect 111818 67974 111830 68026
rect 111882 67974 111894 68026
rect 111946 67974 111958 68026
rect 112010 67974 142486 68026
rect 142538 67974 142550 68026
rect 142602 67974 142614 68026
rect 142666 67974 142678 68026
rect 142730 67974 173206 68026
rect 173258 67974 173270 68026
rect 173322 67974 173334 68026
rect 173386 67974 173398 68026
rect 173450 67974 178848 68026
rect 1104 67952 178848 67974
rect 1104 67482 178848 67504
rect 1104 67430 4246 67482
rect 4298 67430 4310 67482
rect 4362 67430 4374 67482
rect 4426 67430 4438 67482
rect 4490 67430 34966 67482
rect 35018 67430 35030 67482
rect 35082 67430 35094 67482
rect 35146 67430 35158 67482
rect 35210 67430 65686 67482
rect 65738 67430 65750 67482
rect 65802 67430 65814 67482
rect 65866 67430 65878 67482
rect 65930 67430 96406 67482
rect 96458 67430 96470 67482
rect 96522 67430 96534 67482
rect 96586 67430 96598 67482
rect 96650 67430 127126 67482
rect 127178 67430 127190 67482
rect 127242 67430 127254 67482
rect 127306 67430 127318 67482
rect 127370 67430 157846 67482
rect 157898 67430 157910 67482
rect 157962 67430 157974 67482
rect 158026 67430 158038 67482
rect 158090 67430 178848 67482
rect 1104 67408 178848 67430
rect 1104 66938 178848 66960
rect 1104 66886 19606 66938
rect 19658 66886 19670 66938
rect 19722 66886 19734 66938
rect 19786 66886 19798 66938
rect 19850 66886 50326 66938
rect 50378 66886 50390 66938
rect 50442 66886 50454 66938
rect 50506 66886 50518 66938
rect 50570 66886 81046 66938
rect 81098 66886 81110 66938
rect 81162 66886 81174 66938
rect 81226 66886 81238 66938
rect 81290 66886 111766 66938
rect 111818 66886 111830 66938
rect 111882 66886 111894 66938
rect 111946 66886 111958 66938
rect 112010 66886 142486 66938
rect 142538 66886 142550 66938
rect 142602 66886 142614 66938
rect 142666 66886 142678 66938
rect 142730 66886 173206 66938
rect 173258 66886 173270 66938
rect 173322 66886 173334 66938
rect 173386 66886 173398 66938
rect 173450 66886 178848 66938
rect 1104 66864 178848 66886
rect 1104 66394 178848 66416
rect 1104 66342 4246 66394
rect 4298 66342 4310 66394
rect 4362 66342 4374 66394
rect 4426 66342 4438 66394
rect 4490 66342 34966 66394
rect 35018 66342 35030 66394
rect 35082 66342 35094 66394
rect 35146 66342 35158 66394
rect 35210 66342 65686 66394
rect 65738 66342 65750 66394
rect 65802 66342 65814 66394
rect 65866 66342 65878 66394
rect 65930 66342 96406 66394
rect 96458 66342 96470 66394
rect 96522 66342 96534 66394
rect 96586 66342 96598 66394
rect 96650 66342 127126 66394
rect 127178 66342 127190 66394
rect 127242 66342 127254 66394
rect 127306 66342 127318 66394
rect 127370 66342 157846 66394
rect 157898 66342 157910 66394
rect 157962 66342 157974 66394
rect 158026 66342 158038 66394
rect 158090 66342 178848 66394
rect 1104 66320 178848 66342
rect 1104 65850 178848 65872
rect 1104 65798 19606 65850
rect 19658 65798 19670 65850
rect 19722 65798 19734 65850
rect 19786 65798 19798 65850
rect 19850 65798 50326 65850
rect 50378 65798 50390 65850
rect 50442 65798 50454 65850
rect 50506 65798 50518 65850
rect 50570 65798 81046 65850
rect 81098 65798 81110 65850
rect 81162 65798 81174 65850
rect 81226 65798 81238 65850
rect 81290 65798 111766 65850
rect 111818 65798 111830 65850
rect 111882 65798 111894 65850
rect 111946 65798 111958 65850
rect 112010 65798 142486 65850
rect 142538 65798 142550 65850
rect 142602 65798 142614 65850
rect 142666 65798 142678 65850
rect 142730 65798 173206 65850
rect 173258 65798 173270 65850
rect 173322 65798 173334 65850
rect 173386 65798 173398 65850
rect 173450 65798 178848 65850
rect 1104 65776 178848 65798
rect 1104 65306 178848 65328
rect 1104 65254 4246 65306
rect 4298 65254 4310 65306
rect 4362 65254 4374 65306
rect 4426 65254 4438 65306
rect 4490 65254 34966 65306
rect 35018 65254 35030 65306
rect 35082 65254 35094 65306
rect 35146 65254 35158 65306
rect 35210 65254 65686 65306
rect 65738 65254 65750 65306
rect 65802 65254 65814 65306
rect 65866 65254 65878 65306
rect 65930 65254 96406 65306
rect 96458 65254 96470 65306
rect 96522 65254 96534 65306
rect 96586 65254 96598 65306
rect 96650 65254 127126 65306
rect 127178 65254 127190 65306
rect 127242 65254 127254 65306
rect 127306 65254 127318 65306
rect 127370 65254 157846 65306
rect 157898 65254 157910 65306
rect 157962 65254 157974 65306
rect 158026 65254 158038 65306
rect 158090 65254 178848 65306
rect 1104 65232 178848 65254
rect 1104 64762 178848 64784
rect 1104 64710 19606 64762
rect 19658 64710 19670 64762
rect 19722 64710 19734 64762
rect 19786 64710 19798 64762
rect 19850 64710 50326 64762
rect 50378 64710 50390 64762
rect 50442 64710 50454 64762
rect 50506 64710 50518 64762
rect 50570 64710 81046 64762
rect 81098 64710 81110 64762
rect 81162 64710 81174 64762
rect 81226 64710 81238 64762
rect 81290 64710 111766 64762
rect 111818 64710 111830 64762
rect 111882 64710 111894 64762
rect 111946 64710 111958 64762
rect 112010 64710 142486 64762
rect 142538 64710 142550 64762
rect 142602 64710 142614 64762
rect 142666 64710 142678 64762
rect 142730 64710 173206 64762
rect 173258 64710 173270 64762
rect 173322 64710 173334 64762
rect 173386 64710 173398 64762
rect 173450 64710 178848 64762
rect 1104 64688 178848 64710
rect 1104 64218 178848 64240
rect 1104 64166 4246 64218
rect 4298 64166 4310 64218
rect 4362 64166 4374 64218
rect 4426 64166 4438 64218
rect 4490 64166 34966 64218
rect 35018 64166 35030 64218
rect 35082 64166 35094 64218
rect 35146 64166 35158 64218
rect 35210 64166 65686 64218
rect 65738 64166 65750 64218
rect 65802 64166 65814 64218
rect 65866 64166 65878 64218
rect 65930 64166 96406 64218
rect 96458 64166 96470 64218
rect 96522 64166 96534 64218
rect 96586 64166 96598 64218
rect 96650 64166 127126 64218
rect 127178 64166 127190 64218
rect 127242 64166 127254 64218
rect 127306 64166 127318 64218
rect 127370 64166 157846 64218
rect 157898 64166 157910 64218
rect 157962 64166 157974 64218
rect 158026 64166 158038 64218
rect 158090 64166 178848 64218
rect 1104 64144 178848 64166
rect 1104 63674 178848 63696
rect 1104 63622 19606 63674
rect 19658 63622 19670 63674
rect 19722 63622 19734 63674
rect 19786 63622 19798 63674
rect 19850 63622 50326 63674
rect 50378 63622 50390 63674
rect 50442 63622 50454 63674
rect 50506 63622 50518 63674
rect 50570 63622 81046 63674
rect 81098 63622 81110 63674
rect 81162 63622 81174 63674
rect 81226 63622 81238 63674
rect 81290 63622 111766 63674
rect 111818 63622 111830 63674
rect 111882 63622 111894 63674
rect 111946 63622 111958 63674
rect 112010 63622 142486 63674
rect 142538 63622 142550 63674
rect 142602 63622 142614 63674
rect 142666 63622 142678 63674
rect 142730 63622 173206 63674
rect 173258 63622 173270 63674
rect 173322 63622 173334 63674
rect 173386 63622 173398 63674
rect 173450 63622 178848 63674
rect 1104 63600 178848 63622
rect 1104 63130 178848 63152
rect 1104 63078 4246 63130
rect 4298 63078 4310 63130
rect 4362 63078 4374 63130
rect 4426 63078 4438 63130
rect 4490 63078 34966 63130
rect 35018 63078 35030 63130
rect 35082 63078 35094 63130
rect 35146 63078 35158 63130
rect 35210 63078 65686 63130
rect 65738 63078 65750 63130
rect 65802 63078 65814 63130
rect 65866 63078 65878 63130
rect 65930 63078 96406 63130
rect 96458 63078 96470 63130
rect 96522 63078 96534 63130
rect 96586 63078 96598 63130
rect 96650 63078 127126 63130
rect 127178 63078 127190 63130
rect 127242 63078 127254 63130
rect 127306 63078 127318 63130
rect 127370 63078 157846 63130
rect 157898 63078 157910 63130
rect 157962 63078 157974 63130
rect 158026 63078 158038 63130
rect 158090 63078 178848 63130
rect 1104 63056 178848 63078
rect 1104 62586 178848 62608
rect 1104 62534 19606 62586
rect 19658 62534 19670 62586
rect 19722 62534 19734 62586
rect 19786 62534 19798 62586
rect 19850 62534 50326 62586
rect 50378 62534 50390 62586
rect 50442 62534 50454 62586
rect 50506 62534 50518 62586
rect 50570 62534 81046 62586
rect 81098 62534 81110 62586
rect 81162 62534 81174 62586
rect 81226 62534 81238 62586
rect 81290 62534 111766 62586
rect 111818 62534 111830 62586
rect 111882 62534 111894 62586
rect 111946 62534 111958 62586
rect 112010 62534 142486 62586
rect 142538 62534 142550 62586
rect 142602 62534 142614 62586
rect 142666 62534 142678 62586
rect 142730 62534 173206 62586
rect 173258 62534 173270 62586
rect 173322 62534 173334 62586
rect 173386 62534 173398 62586
rect 173450 62534 178848 62586
rect 1104 62512 178848 62534
rect 1104 62042 178848 62064
rect 1104 61990 4246 62042
rect 4298 61990 4310 62042
rect 4362 61990 4374 62042
rect 4426 61990 4438 62042
rect 4490 61990 34966 62042
rect 35018 61990 35030 62042
rect 35082 61990 35094 62042
rect 35146 61990 35158 62042
rect 35210 61990 65686 62042
rect 65738 61990 65750 62042
rect 65802 61990 65814 62042
rect 65866 61990 65878 62042
rect 65930 61990 96406 62042
rect 96458 61990 96470 62042
rect 96522 61990 96534 62042
rect 96586 61990 96598 62042
rect 96650 61990 127126 62042
rect 127178 61990 127190 62042
rect 127242 61990 127254 62042
rect 127306 61990 127318 62042
rect 127370 61990 157846 62042
rect 157898 61990 157910 62042
rect 157962 61990 157974 62042
rect 158026 61990 158038 62042
rect 158090 61990 178848 62042
rect 1104 61968 178848 61990
rect 1104 61498 178848 61520
rect 1104 61446 19606 61498
rect 19658 61446 19670 61498
rect 19722 61446 19734 61498
rect 19786 61446 19798 61498
rect 19850 61446 50326 61498
rect 50378 61446 50390 61498
rect 50442 61446 50454 61498
rect 50506 61446 50518 61498
rect 50570 61446 81046 61498
rect 81098 61446 81110 61498
rect 81162 61446 81174 61498
rect 81226 61446 81238 61498
rect 81290 61446 111766 61498
rect 111818 61446 111830 61498
rect 111882 61446 111894 61498
rect 111946 61446 111958 61498
rect 112010 61446 142486 61498
rect 142538 61446 142550 61498
rect 142602 61446 142614 61498
rect 142666 61446 142678 61498
rect 142730 61446 173206 61498
rect 173258 61446 173270 61498
rect 173322 61446 173334 61498
rect 173386 61446 173398 61498
rect 173450 61446 178848 61498
rect 1104 61424 178848 61446
rect 1104 60954 178848 60976
rect 1104 60902 4246 60954
rect 4298 60902 4310 60954
rect 4362 60902 4374 60954
rect 4426 60902 4438 60954
rect 4490 60902 34966 60954
rect 35018 60902 35030 60954
rect 35082 60902 35094 60954
rect 35146 60902 35158 60954
rect 35210 60902 65686 60954
rect 65738 60902 65750 60954
rect 65802 60902 65814 60954
rect 65866 60902 65878 60954
rect 65930 60902 96406 60954
rect 96458 60902 96470 60954
rect 96522 60902 96534 60954
rect 96586 60902 96598 60954
rect 96650 60902 127126 60954
rect 127178 60902 127190 60954
rect 127242 60902 127254 60954
rect 127306 60902 127318 60954
rect 127370 60902 157846 60954
rect 157898 60902 157910 60954
rect 157962 60902 157974 60954
rect 158026 60902 158038 60954
rect 158090 60902 178848 60954
rect 1104 60880 178848 60902
rect 1104 60410 178848 60432
rect 1104 60358 19606 60410
rect 19658 60358 19670 60410
rect 19722 60358 19734 60410
rect 19786 60358 19798 60410
rect 19850 60358 50326 60410
rect 50378 60358 50390 60410
rect 50442 60358 50454 60410
rect 50506 60358 50518 60410
rect 50570 60358 81046 60410
rect 81098 60358 81110 60410
rect 81162 60358 81174 60410
rect 81226 60358 81238 60410
rect 81290 60358 111766 60410
rect 111818 60358 111830 60410
rect 111882 60358 111894 60410
rect 111946 60358 111958 60410
rect 112010 60358 142486 60410
rect 142538 60358 142550 60410
rect 142602 60358 142614 60410
rect 142666 60358 142678 60410
rect 142730 60358 173206 60410
rect 173258 60358 173270 60410
rect 173322 60358 173334 60410
rect 173386 60358 173398 60410
rect 173450 60358 178848 60410
rect 1104 60336 178848 60358
rect 1857 60163 1915 60169
rect 1857 60129 1869 60163
rect 1903 60160 1915 60163
rect 3050 60160 3056 60172
rect 1903 60132 3056 60160
rect 1903 60129 1915 60132
rect 1857 60123 1915 60129
rect 3050 60120 3056 60132
rect 3108 60120 3114 60172
rect 176930 60120 176936 60172
rect 176988 60160 176994 60172
rect 177945 60163 178003 60169
rect 177945 60160 177957 60163
rect 176988 60132 177957 60160
rect 176988 60120 176994 60132
rect 177945 60129 177957 60132
rect 177991 60129 178003 60163
rect 177945 60123 178003 60129
rect 2038 60024 2044 60036
rect 1999 59996 2044 60024
rect 2038 59984 2044 59996
rect 2096 59984 2102 60036
rect 178126 60024 178132 60036
rect 178087 59996 178132 60024
rect 178126 59984 178132 59996
rect 178184 59984 178190 60036
rect 1104 59866 178848 59888
rect 1104 59814 4246 59866
rect 4298 59814 4310 59866
rect 4362 59814 4374 59866
rect 4426 59814 4438 59866
rect 4490 59814 34966 59866
rect 35018 59814 35030 59866
rect 35082 59814 35094 59866
rect 35146 59814 35158 59866
rect 35210 59814 65686 59866
rect 65738 59814 65750 59866
rect 65802 59814 65814 59866
rect 65866 59814 65878 59866
rect 65930 59814 96406 59866
rect 96458 59814 96470 59866
rect 96522 59814 96534 59866
rect 96586 59814 96598 59866
rect 96650 59814 127126 59866
rect 127178 59814 127190 59866
rect 127242 59814 127254 59866
rect 127306 59814 127318 59866
rect 127370 59814 157846 59866
rect 157898 59814 157910 59866
rect 157962 59814 157974 59866
rect 158026 59814 158038 59866
rect 158090 59814 178848 59866
rect 1104 59792 178848 59814
rect 3050 59752 3056 59764
rect 3011 59724 3056 59752
rect 3050 59712 3056 59724
rect 3108 59712 3114 59764
rect 176930 59752 176936 59764
rect 176891 59724 176936 59752
rect 176930 59712 176936 59724
rect 176988 59712 176994 59764
rect 1104 59322 178848 59344
rect 1104 59270 19606 59322
rect 19658 59270 19670 59322
rect 19722 59270 19734 59322
rect 19786 59270 19798 59322
rect 19850 59270 50326 59322
rect 50378 59270 50390 59322
rect 50442 59270 50454 59322
rect 50506 59270 50518 59322
rect 50570 59270 81046 59322
rect 81098 59270 81110 59322
rect 81162 59270 81174 59322
rect 81226 59270 81238 59322
rect 81290 59270 111766 59322
rect 111818 59270 111830 59322
rect 111882 59270 111894 59322
rect 111946 59270 111958 59322
rect 112010 59270 142486 59322
rect 142538 59270 142550 59322
rect 142602 59270 142614 59322
rect 142666 59270 142678 59322
rect 142730 59270 173206 59322
rect 173258 59270 173270 59322
rect 173322 59270 173334 59322
rect 173386 59270 173398 59322
rect 173450 59270 178848 59322
rect 1104 59248 178848 59270
rect 1104 58778 178848 58800
rect 1104 58726 4246 58778
rect 4298 58726 4310 58778
rect 4362 58726 4374 58778
rect 4426 58726 4438 58778
rect 4490 58726 34966 58778
rect 35018 58726 35030 58778
rect 35082 58726 35094 58778
rect 35146 58726 35158 58778
rect 35210 58726 65686 58778
rect 65738 58726 65750 58778
rect 65802 58726 65814 58778
rect 65866 58726 65878 58778
rect 65930 58726 96406 58778
rect 96458 58726 96470 58778
rect 96522 58726 96534 58778
rect 96586 58726 96598 58778
rect 96650 58726 127126 58778
rect 127178 58726 127190 58778
rect 127242 58726 127254 58778
rect 127306 58726 127318 58778
rect 127370 58726 157846 58778
rect 157898 58726 157910 58778
rect 157962 58726 157974 58778
rect 158026 58726 158038 58778
rect 158090 58726 178848 58778
rect 1104 58704 178848 58726
rect 1104 58234 178848 58256
rect 1104 58182 19606 58234
rect 19658 58182 19670 58234
rect 19722 58182 19734 58234
rect 19786 58182 19798 58234
rect 19850 58182 50326 58234
rect 50378 58182 50390 58234
rect 50442 58182 50454 58234
rect 50506 58182 50518 58234
rect 50570 58182 81046 58234
rect 81098 58182 81110 58234
rect 81162 58182 81174 58234
rect 81226 58182 81238 58234
rect 81290 58182 111766 58234
rect 111818 58182 111830 58234
rect 111882 58182 111894 58234
rect 111946 58182 111958 58234
rect 112010 58182 142486 58234
rect 142538 58182 142550 58234
rect 142602 58182 142614 58234
rect 142666 58182 142678 58234
rect 142730 58182 173206 58234
rect 173258 58182 173270 58234
rect 173322 58182 173334 58234
rect 173386 58182 173398 58234
rect 173450 58182 178848 58234
rect 1104 58160 178848 58182
rect 1104 57690 178848 57712
rect 1104 57638 4246 57690
rect 4298 57638 4310 57690
rect 4362 57638 4374 57690
rect 4426 57638 4438 57690
rect 4490 57638 34966 57690
rect 35018 57638 35030 57690
rect 35082 57638 35094 57690
rect 35146 57638 35158 57690
rect 35210 57638 65686 57690
rect 65738 57638 65750 57690
rect 65802 57638 65814 57690
rect 65866 57638 65878 57690
rect 65930 57638 96406 57690
rect 96458 57638 96470 57690
rect 96522 57638 96534 57690
rect 96586 57638 96598 57690
rect 96650 57638 127126 57690
rect 127178 57638 127190 57690
rect 127242 57638 127254 57690
rect 127306 57638 127318 57690
rect 127370 57638 157846 57690
rect 157898 57638 157910 57690
rect 157962 57638 157974 57690
rect 158026 57638 158038 57690
rect 158090 57638 178848 57690
rect 1104 57616 178848 57638
rect 1104 57146 178848 57168
rect 1104 57094 19606 57146
rect 19658 57094 19670 57146
rect 19722 57094 19734 57146
rect 19786 57094 19798 57146
rect 19850 57094 50326 57146
rect 50378 57094 50390 57146
rect 50442 57094 50454 57146
rect 50506 57094 50518 57146
rect 50570 57094 81046 57146
rect 81098 57094 81110 57146
rect 81162 57094 81174 57146
rect 81226 57094 81238 57146
rect 81290 57094 111766 57146
rect 111818 57094 111830 57146
rect 111882 57094 111894 57146
rect 111946 57094 111958 57146
rect 112010 57094 142486 57146
rect 142538 57094 142550 57146
rect 142602 57094 142614 57146
rect 142666 57094 142678 57146
rect 142730 57094 173206 57146
rect 173258 57094 173270 57146
rect 173322 57094 173334 57146
rect 173386 57094 173398 57146
rect 173450 57094 178848 57146
rect 1104 57072 178848 57094
rect 1104 56602 178848 56624
rect 1104 56550 4246 56602
rect 4298 56550 4310 56602
rect 4362 56550 4374 56602
rect 4426 56550 4438 56602
rect 4490 56550 34966 56602
rect 35018 56550 35030 56602
rect 35082 56550 35094 56602
rect 35146 56550 35158 56602
rect 35210 56550 65686 56602
rect 65738 56550 65750 56602
rect 65802 56550 65814 56602
rect 65866 56550 65878 56602
rect 65930 56550 96406 56602
rect 96458 56550 96470 56602
rect 96522 56550 96534 56602
rect 96586 56550 96598 56602
rect 96650 56550 127126 56602
rect 127178 56550 127190 56602
rect 127242 56550 127254 56602
rect 127306 56550 127318 56602
rect 127370 56550 157846 56602
rect 157898 56550 157910 56602
rect 157962 56550 157974 56602
rect 158026 56550 158038 56602
rect 158090 56550 178848 56602
rect 1104 56528 178848 56550
rect 1104 56058 178848 56080
rect 1104 56006 19606 56058
rect 19658 56006 19670 56058
rect 19722 56006 19734 56058
rect 19786 56006 19798 56058
rect 19850 56006 50326 56058
rect 50378 56006 50390 56058
rect 50442 56006 50454 56058
rect 50506 56006 50518 56058
rect 50570 56006 81046 56058
rect 81098 56006 81110 56058
rect 81162 56006 81174 56058
rect 81226 56006 81238 56058
rect 81290 56006 111766 56058
rect 111818 56006 111830 56058
rect 111882 56006 111894 56058
rect 111946 56006 111958 56058
rect 112010 56006 142486 56058
rect 142538 56006 142550 56058
rect 142602 56006 142614 56058
rect 142666 56006 142678 56058
rect 142730 56006 173206 56058
rect 173258 56006 173270 56058
rect 173322 56006 173334 56058
rect 173386 56006 173398 56058
rect 173450 56006 178848 56058
rect 1104 55984 178848 56006
rect 1104 55514 178848 55536
rect 1104 55462 4246 55514
rect 4298 55462 4310 55514
rect 4362 55462 4374 55514
rect 4426 55462 4438 55514
rect 4490 55462 34966 55514
rect 35018 55462 35030 55514
rect 35082 55462 35094 55514
rect 35146 55462 35158 55514
rect 35210 55462 65686 55514
rect 65738 55462 65750 55514
rect 65802 55462 65814 55514
rect 65866 55462 65878 55514
rect 65930 55462 96406 55514
rect 96458 55462 96470 55514
rect 96522 55462 96534 55514
rect 96586 55462 96598 55514
rect 96650 55462 127126 55514
rect 127178 55462 127190 55514
rect 127242 55462 127254 55514
rect 127306 55462 127318 55514
rect 127370 55462 157846 55514
rect 157898 55462 157910 55514
rect 157962 55462 157974 55514
rect 158026 55462 158038 55514
rect 158090 55462 178848 55514
rect 1104 55440 178848 55462
rect 1104 54970 178848 54992
rect 1104 54918 19606 54970
rect 19658 54918 19670 54970
rect 19722 54918 19734 54970
rect 19786 54918 19798 54970
rect 19850 54918 50326 54970
rect 50378 54918 50390 54970
rect 50442 54918 50454 54970
rect 50506 54918 50518 54970
rect 50570 54918 81046 54970
rect 81098 54918 81110 54970
rect 81162 54918 81174 54970
rect 81226 54918 81238 54970
rect 81290 54918 111766 54970
rect 111818 54918 111830 54970
rect 111882 54918 111894 54970
rect 111946 54918 111958 54970
rect 112010 54918 142486 54970
rect 142538 54918 142550 54970
rect 142602 54918 142614 54970
rect 142666 54918 142678 54970
rect 142730 54918 173206 54970
rect 173258 54918 173270 54970
rect 173322 54918 173334 54970
rect 173386 54918 173398 54970
rect 173450 54918 178848 54970
rect 1104 54896 178848 54918
rect 1104 54426 178848 54448
rect 1104 54374 4246 54426
rect 4298 54374 4310 54426
rect 4362 54374 4374 54426
rect 4426 54374 4438 54426
rect 4490 54374 34966 54426
rect 35018 54374 35030 54426
rect 35082 54374 35094 54426
rect 35146 54374 35158 54426
rect 35210 54374 65686 54426
rect 65738 54374 65750 54426
rect 65802 54374 65814 54426
rect 65866 54374 65878 54426
rect 65930 54374 96406 54426
rect 96458 54374 96470 54426
rect 96522 54374 96534 54426
rect 96586 54374 96598 54426
rect 96650 54374 127126 54426
rect 127178 54374 127190 54426
rect 127242 54374 127254 54426
rect 127306 54374 127318 54426
rect 127370 54374 157846 54426
rect 157898 54374 157910 54426
rect 157962 54374 157974 54426
rect 158026 54374 158038 54426
rect 158090 54374 178848 54426
rect 1104 54352 178848 54374
rect 1104 53882 178848 53904
rect 1104 53830 19606 53882
rect 19658 53830 19670 53882
rect 19722 53830 19734 53882
rect 19786 53830 19798 53882
rect 19850 53830 50326 53882
rect 50378 53830 50390 53882
rect 50442 53830 50454 53882
rect 50506 53830 50518 53882
rect 50570 53830 81046 53882
rect 81098 53830 81110 53882
rect 81162 53830 81174 53882
rect 81226 53830 81238 53882
rect 81290 53830 111766 53882
rect 111818 53830 111830 53882
rect 111882 53830 111894 53882
rect 111946 53830 111958 53882
rect 112010 53830 142486 53882
rect 142538 53830 142550 53882
rect 142602 53830 142614 53882
rect 142666 53830 142678 53882
rect 142730 53830 173206 53882
rect 173258 53830 173270 53882
rect 173322 53830 173334 53882
rect 173386 53830 173398 53882
rect 173450 53830 178848 53882
rect 1104 53808 178848 53830
rect 1104 53338 178848 53360
rect 1104 53286 4246 53338
rect 4298 53286 4310 53338
rect 4362 53286 4374 53338
rect 4426 53286 4438 53338
rect 4490 53286 34966 53338
rect 35018 53286 35030 53338
rect 35082 53286 35094 53338
rect 35146 53286 35158 53338
rect 35210 53286 65686 53338
rect 65738 53286 65750 53338
rect 65802 53286 65814 53338
rect 65866 53286 65878 53338
rect 65930 53286 96406 53338
rect 96458 53286 96470 53338
rect 96522 53286 96534 53338
rect 96586 53286 96598 53338
rect 96650 53286 127126 53338
rect 127178 53286 127190 53338
rect 127242 53286 127254 53338
rect 127306 53286 127318 53338
rect 127370 53286 157846 53338
rect 157898 53286 157910 53338
rect 157962 53286 157974 53338
rect 158026 53286 158038 53338
rect 158090 53286 178848 53338
rect 1104 53264 178848 53286
rect 1104 52794 178848 52816
rect 1104 52742 19606 52794
rect 19658 52742 19670 52794
rect 19722 52742 19734 52794
rect 19786 52742 19798 52794
rect 19850 52742 50326 52794
rect 50378 52742 50390 52794
rect 50442 52742 50454 52794
rect 50506 52742 50518 52794
rect 50570 52742 81046 52794
rect 81098 52742 81110 52794
rect 81162 52742 81174 52794
rect 81226 52742 81238 52794
rect 81290 52742 111766 52794
rect 111818 52742 111830 52794
rect 111882 52742 111894 52794
rect 111946 52742 111958 52794
rect 112010 52742 142486 52794
rect 142538 52742 142550 52794
rect 142602 52742 142614 52794
rect 142666 52742 142678 52794
rect 142730 52742 173206 52794
rect 173258 52742 173270 52794
rect 173322 52742 173334 52794
rect 173386 52742 173398 52794
rect 173450 52742 178848 52794
rect 1104 52720 178848 52742
rect 1104 52250 178848 52272
rect 1104 52198 4246 52250
rect 4298 52198 4310 52250
rect 4362 52198 4374 52250
rect 4426 52198 4438 52250
rect 4490 52198 34966 52250
rect 35018 52198 35030 52250
rect 35082 52198 35094 52250
rect 35146 52198 35158 52250
rect 35210 52198 65686 52250
rect 65738 52198 65750 52250
rect 65802 52198 65814 52250
rect 65866 52198 65878 52250
rect 65930 52198 96406 52250
rect 96458 52198 96470 52250
rect 96522 52198 96534 52250
rect 96586 52198 96598 52250
rect 96650 52198 127126 52250
rect 127178 52198 127190 52250
rect 127242 52198 127254 52250
rect 127306 52198 127318 52250
rect 127370 52198 157846 52250
rect 157898 52198 157910 52250
rect 157962 52198 157974 52250
rect 158026 52198 158038 52250
rect 158090 52198 178848 52250
rect 1104 52176 178848 52198
rect 1104 51706 178848 51728
rect 1104 51654 19606 51706
rect 19658 51654 19670 51706
rect 19722 51654 19734 51706
rect 19786 51654 19798 51706
rect 19850 51654 50326 51706
rect 50378 51654 50390 51706
rect 50442 51654 50454 51706
rect 50506 51654 50518 51706
rect 50570 51654 81046 51706
rect 81098 51654 81110 51706
rect 81162 51654 81174 51706
rect 81226 51654 81238 51706
rect 81290 51654 111766 51706
rect 111818 51654 111830 51706
rect 111882 51654 111894 51706
rect 111946 51654 111958 51706
rect 112010 51654 142486 51706
rect 142538 51654 142550 51706
rect 142602 51654 142614 51706
rect 142666 51654 142678 51706
rect 142730 51654 173206 51706
rect 173258 51654 173270 51706
rect 173322 51654 173334 51706
rect 173386 51654 173398 51706
rect 173450 51654 178848 51706
rect 1104 51632 178848 51654
rect 1104 51162 178848 51184
rect 1104 51110 4246 51162
rect 4298 51110 4310 51162
rect 4362 51110 4374 51162
rect 4426 51110 4438 51162
rect 4490 51110 34966 51162
rect 35018 51110 35030 51162
rect 35082 51110 35094 51162
rect 35146 51110 35158 51162
rect 35210 51110 65686 51162
rect 65738 51110 65750 51162
rect 65802 51110 65814 51162
rect 65866 51110 65878 51162
rect 65930 51110 96406 51162
rect 96458 51110 96470 51162
rect 96522 51110 96534 51162
rect 96586 51110 96598 51162
rect 96650 51110 127126 51162
rect 127178 51110 127190 51162
rect 127242 51110 127254 51162
rect 127306 51110 127318 51162
rect 127370 51110 157846 51162
rect 157898 51110 157910 51162
rect 157962 51110 157974 51162
rect 158026 51110 158038 51162
rect 158090 51110 178848 51162
rect 1104 51088 178848 51110
rect 1104 50618 178848 50640
rect 1104 50566 19606 50618
rect 19658 50566 19670 50618
rect 19722 50566 19734 50618
rect 19786 50566 19798 50618
rect 19850 50566 50326 50618
rect 50378 50566 50390 50618
rect 50442 50566 50454 50618
rect 50506 50566 50518 50618
rect 50570 50566 81046 50618
rect 81098 50566 81110 50618
rect 81162 50566 81174 50618
rect 81226 50566 81238 50618
rect 81290 50566 111766 50618
rect 111818 50566 111830 50618
rect 111882 50566 111894 50618
rect 111946 50566 111958 50618
rect 112010 50566 142486 50618
rect 142538 50566 142550 50618
rect 142602 50566 142614 50618
rect 142666 50566 142678 50618
rect 142730 50566 173206 50618
rect 173258 50566 173270 50618
rect 173322 50566 173334 50618
rect 173386 50566 173398 50618
rect 173450 50566 178848 50618
rect 1104 50544 178848 50566
rect 1104 50074 178848 50096
rect 1104 50022 4246 50074
rect 4298 50022 4310 50074
rect 4362 50022 4374 50074
rect 4426 50022 4438 50074
rect 4490 50022 34966 50074
rect 35018 50022 35030 50074
rect 35082 50022 35094 50074
rect 35146 50022 35158 50074
rect 35210 50022 65686 50074
rect 65738 50022 65750 50074
rect 65802 50022 65814 50074
rect 65866 50022 65878 50074
rect 65930 50022 96406 50074
rect 96458 50022 96470 50074
rect 96522 50022 96534 50074
rect 96586 50022 96598 50074
rect 96650 50022 127126 50074
rect 127178 50022 127190 50074
rect 127242 50022 127254 50074
rect 127306 50022 127318 50074
rect 127370 50022 157846 50074
rect 157898 50022 157910 50074
rect 157962 50022 157974 50074
rect 158026 50022 158038 50074
rect 158090 50022 178848 50074
rect 1104 50000 178848 50022
rect 1104 49530 178848 49552
rect 1104 49478 19606 49530
rect 19658 49478 19670 49530
rect 19722 49478 19734 49530
rect 19786 49478 19798 49530
rect 19850 49478 50326 49530
rect 50378 49478 50390 49530
rect 50442 49478 50454 49530
rect 50506 49478 50518 49530
rect 50570 49478 81046 49530
rect 81098 49478 81110 49530
rect 81162 49478 81174 49530
rect 81226 49478 81238 49530
rect 81290 49478 111766 49530
rect 111818 49478 111830 49530
rect 111882 49478 111894 49530
rect 111946 49478 111958 49530
rect 112010 49478 142486 49530
rect 142538 49478 142550 49530
rect 142602 49478 142614 49530
rect 142666 49478 142678 49530
rect 142730 49478 173206 49530
rect 173258 49478 173270 49530
rect 173322 49478 173334 49530
rect 173386 49478 173398 49530
rect 173450 49478 178848 49530
rect 1104 49456 178848 49478
rect 1104 48986 178848 49008
rect 1104 48934 4246 48986
rect 4298 48934 4310 48986
rect 4362 48934 4374 48986
rect 4426 48934 4438 48986
rect 4490 48934 34966 48986
rect 35018 48934 35030 48986
rect 35082 48934 35094 48986
rect 35146 48934 35158 48986
rect 35210 48934 65686 48986
rect 65738 48934 65750 48986
rect 65802 48934 65814 48986
rect 65866 48934 65878 48986
rect 65930 48934 96406 48986
rect 96458 48934 96470 48986
rect 96522 48934 96534 48986
rect 96586 48934 96598 48986
rect 96650 48934 127126 48986
rect 127178 48934 127190 48986
rect 127242 48934 127254 48986
rect 127306 48934 127318 48986
rect 127370 48934 157846 48986
rect 157898 48934 157910 48986
rect 157962 48934 157974 48986
rect 158026 48934 158038 48986
rect 158090 48934 178848 48986
rect 1104 48912 178848 48934
rect 1104 48442 178848 48464
rect 1104 48390 19606 48442
rect 19658 48390 19670 48442
rect 19722 48390 19734 48442
rect 19786 48390 19798 48442
rect 19850 48390 50326 48442
rect 50378 48390 50390 48442
rect 50442 48390 50454 48442
rect 50506 48390 50518 48442
rect 50570 48390 81046 48442
rect 81098 48390 81110 48442
rect 81162 48390 81174 48442
rect 81226 48390 81238 48442
rect 81290 48390 111766 48442
rect 111818 48390 111830 48442
rect 111882 48390 111894 48442
rect 111946 48390 111958 48442
rect 112010 48390 142486 48442
rect 142538 48390 142550 48442
rect 142602 48390 142614 48442
rect 142666 48390 142678 48442
rect 142730 48390 173206 48442
rect 173258 48390 173270 48442
rect 173322 48390 173334 48442
rect 173386 48390 173398 48442
rect 173450 48390 178848 48442
rect 1104 48368 178848 48390
rect 1104 47898 178848 47920
rect 1104 47846 4246 47898
rect 4298 47846 4310 47898
rect 4362 47846 4374 47898
rect 4426 47846 4438 47898
rect 4490 47846 34966 47898
rect 35018 47846 35030 47898
rect 35082 47846 35094 47898
rect 35146 47846 35158 47898
rect 35210 47846 65686 47898
rect 65738 47846 65750 47898
rect 65802 47846 65814 47898
rect 65866 47846 65878 47898
rect 65930 47846 96406 47898
rect 96458 47846 96470 47898
rect 96522 47846 96534 47898
rect 96586 47846 96598 47898
rect 96650 47846 127126 47898
rect 127178 47846 127190 47898
rect 127242 47846 127254 47898
rect 127306 47846 127318 47898
rect 127370 47846 157846 47898
rect 157898 47846 157910 47898
rect 157962 47846 157974 47898
rect 158026 47846 158038 47898
rect 158090 47846 178848 47898
rect 1104 47824 178848 47846
rect 1104 47354 178848 47376
rect 1104 47302 19606 47354
rect 19658 47302 19670 47354
rect 19722 47302 19734 47354
rect 19786 47302 19798 47354
rect 19850 47302 50326 47354
rect 50378 47302 50390 47354
rect 50442 47302 50454 47354
rect 50506 47302 50518 47354
rect 50570 47302 81046 47354
rect 81098 47302 81110 47354
rect 81162 47302 81174 47354
rect 81226 47302 81238 47354
rect 81290 47302 111766 47354
rect 111818 47302 111830 47354
rect 111882 47302 111894 47354
rect 111946 47302 111958 47354
rect 112010 47302 142486 47354
rect 142538 47302 142550 47354
rect 142602 47302 142614 47354
rect 142666 47302 142678 47354
rect 142730 47302 173206 47354
rect 173258 47302 173270 47354
rect 173322 47302 173334 47354
rect 173386 47302 173398 47354
rect 173450 47302 178848 47354
rect 1104 47280 178848 47302
rect 1104 46810 178848 46832
rect 1104 46758 4246 46810
rect 4298 46758 4310 46810
rect 4362 46758 4374 46810
rect 4426 46758 4438 46810
rect 4490 46758 34966 46810
rect 35018 46758 35030 46810
rect 35082 46758 35094 46810
rect 35146 46758 35158 46810
rect 35210 46758 65686 46810
rect 65738 46758 65750 46810
rect 65802 46758 65814 46810
rect 65866 46758 65878 46810
rect 65930 46758 96406 46810
rect 96458 46758 96470 46810
rect 96522 46758 96534 46810
rect 96586 46758 96598 46810
rect 96650 46758 127126 46810
rect 127178 46758 127190 46810
rect 127242 46758 127254 46810
rect 127306 46758 127318 46810
rect 127370 46758 157846 46810
rect 157898 46758 157910 46810
rect 157962 46758 157974 46810
rect 158026 46758 158038 46810
rect 158090 46758 178848 46810
rect 1104 46736 178848 46758
rect 1104 46266 178848 46288
rect 1104 46214 19606 46266
rect 19658 46214 19670 46266
rect 19722 46214 19734 46266
rect 19786 46214 19798 46266
rect 19850 46214 50326 46266
rect 50378 46214 50390 46266
rect 50442 46214 50454 46266
rect 50506 46214 50518 46266
rect 50570 46214 81046 46266
rect 81098 46214 81110 46266
rect 81162 46214 81174 46266
rect 81226 46214 81238 46266
rect 81290 46214 111766 46266
rect 111818 46214 111830 46266
rect 111882 46214 111894 46266
rect 111946 46214 111958 46266
rect 112010 46214 142486 46266
rect 142538 46214 142550 46266
rect 142602 46214 142614 46266
rect 142666 46214 142678 46266
rect 142730 46214 173206 46266
rect 173258 46214 173270 46266
rect 173322 46214 173334 46266
rect 173386 46214 173398 46266
rect 173450 46214 178848 46266
rect 1104 46192 178848 46214
rect 1104 45722 178848 45744
rect 1104 45670 4246 45722
rect 4298 45670 4310 45722
rect 4362 45670 4374 45722
rect 4426 45670 4438 45722
rect 4490 45670 34966 45722
rect 35018 45670 35030 45722
rect 35082 45670 35094 45722
rect 35146 45670 35158 45722
rect 35210 45670 65686 45722
rect 65738 45670 65750 45722
rect 65802 45670 65814 45722
rect 65866 45670 65878 45722
rect 65930 45670 96406 45722
rect 96458 45670 96470 45722
rect 96522 45670 96534 45722
rect 96586 45670 96598 45722
rect 96650 45670 127126 45722
rect 127178 45670 127190 45722
rect 127242 45670 127254 45722
rect 127306 45670 127318 45722
rect 127370 45670 157846 45722
rect 157898 45670 157910 45722
rect 157962 45670 157974 45722
rect 158026 45670 158038 45722
rect 158090 45670 178848 45722
rect 1104 45648 178848 45670
rect 1104 45178 178848 45200
rect 1104 45126 19606 45178
rect 19658 45126 19670 45178
rect 19722 45126 19734 45178
rect 19786 45126 19798 45178
rect 19850 45126 50326 45178
rect 50378 45126 50390 45178
rect 50442 45126 50454 45178
rect 50506 45126 50518 45178
rect 50570 45126 81046 45178
rect 81098 45126 81110 45178
rect 81162 45126 81174 45178
rect 81226 45126 81238 45178
rect 81290 45126 111766 45178
rect 111818 45126 111830 45178
rect 111882 45126 111894 45178
rect 111946 45126 111958 45178
rect 112010 45126 142486 45178
rect 142538 45126 142550 45178
rect 142602 45126 142614 45178
rect 142666 45126 142678 45178
rect 142730 45126 173206 45178
rect 173258 45126 173270 45178
rect 173322 45126 173334 45178
rect 173386 45126 173398 45178
rect 173450 45126 178848 45178
rect 1104 45104 178848 45126
rect 1104 44634 178848 44656
rect 1104 44582 4246 44634
rect 4298 44582 4310 44634
rect 4362 44582 4374 44634
rect 4426 44582 4438 44634
rect 4490 44582 34966 44634
rect 35018 44582 35030 44634
rect 35082 44582 35094 44634
rect 35146 44582 35158 44634
rect 35210 44582 65686 44634
rect 65738 44582 65750 44634
rect 65802 44582 65814 44634
rect 65866 44582 65878 44634
rect 65930 44582 96406 44634
rect 96458 44582 96470 44634
rect 96522 44582 96534 44634
rect 96586 44582 96598 44634
rect 96650 44582 127126 44634
rect 127178 44582 127190 44634
rect 127242 44582 127254 44634
rect 127306 44582 127318 44634
rect 127370 44582 157846 44634
rect 157898 44582 157910 44634
rect 157962 44582 157974 44634
rect 158026 44582 158038 44634
rect 158090 44582 178848 44634
rect 1104 44560 178848 44582
rect 1104 44090 178848 44112
rect 1104 44038 19606 44090
rect 19658 44038 19670 44090
rect 19722 44038 19734 44090
rect 19786 44038 19798 44090
rect 19850 44038 50326 44090
rect 50378 44038 50390 44090
rect 50442 44038 50454 44090
rect 50506 44038 50518 44090
rect 50570 44038 81046 44090
rect 81098 44038 81110 44090
rect 81162 44038 81174 44090
rect 81226 44038 81238 44090
rect 81290 44038 111766 44090
rect 111818 44038 111830 44090
rect 111882 44038 111894 44090
rect 111946 44038 111958 44090
rect 112010 44038 142486 44090
rect 142538 44038 142550 44090
rect 142602 44038 142614 44090
rect 142666 44038 142678 44090
rect 142730 44038 173206 44090
rect 173258 44038 173270 44090
rect 173322 44038 173334 44090
rect 173386 44038 173398 44090
rect 173450 44038 178848 44090
rect 1104 44016 178848 44038
rect 1104 43546 178848 43568
rect 1104 43494 4246 43546
rect 4298 43494 4310 43546
rect 4362 43494 4374 43546
rect 4426 43494 4438 43546
rect 4490 43494 34966 43546
rect 35018 43494 35030 43546
rect 35082 43494 35094 43546
rect 35146 43494 35158 43546
rect 35210 43494 65686 43546
rect 65738 43494 65750 43546
rect 65802 43494 65814 43546
rect 65866 43494 65878 43546
rect 65930 43494 96406 43546
rect 96458 43494 96470 43546
rect 96522 43494 96534 43546
rect 96586 43494 96598 43546
rect 96650 43494 127126 43546
rect 127178 43494 127190 43546
rect 127242 43494 127254 43546
rect 127306 43494 127318 43546
rect 127370 43494 157846 43546
rect 157898 43494 157910 43546
rect 157962 43494 157974 43546
rect 158026 43494 158038 43546
rect 158090 43494 178848 43546
rect 1104 43472 178848 43494
rect 1104 43002 178848 43024
rect 1104 42950 19606 43002
rect 19658 42950 19670 43002
rect 19722 42950 19734 43002
rect 19786 42950 19798 43002
rect 19850 42950 50326 43002
rect 50378 42950 50390 43002
rect 50442 42950 50454 43002
rect 50506 42950 50518 43002
rect 50570 42950 81046 43002
rect 81098 42950 81110 43002
rect 81162 42950 81174 43002
rect 81226 42950 81238 43002
rect 81290 42950 111766 43002
rect 111818 42950 111830 43002
rect 111882 42950 111894 43002
rect 111946 42950 111958 43002
rect 112010 42950 142486 43002
rect 142538 42950 142550 43002
rect 142602 42950 142614 43002
rect 142666 42950 142678 43002
rect 142730 42950 173206 43002
rect 173258 42950 173270 43002
rect 173322 42950 173334 43002
rect 173386 42950 173398 43002
rect 173450 42950 178848 43002
rect 1104 42928 178848 42950
rect 1104 42458 178848 42480
rect 1104 42406 4246 42458
rect 4298 42406 4310 42458
rect 4362 42406 4374 42458
rect 4426 42406 4438 42458
rect 4490 42406 34966 42458
rect 35018 42406 35030 42458
rect 35082 42406 35094 42458
rect 35146 42406 35158 42458
rect 35210 42406 65686 42458
rect 65738 42406 65750 42458
rect 65802 42406 65814 42458
rect 65866 42406 65878 42458
rect 65930 42406 96406 42458
rect 96458 42406 96470 42458
rect 96522 42406 96534 42458
rect 96586 42406 96598 42458
rect 96650 42406 127126 42458
rect 127178 42406 127190 42458
rect 127242 42406 127254 42458
rect 127306 42406 127318 42458
rect 127370 42406 157846 42458
rect 157898 42406 157910 42458
rect 157962 42406 157974 42458
rect 158026 42406 158038 42458
rect 158090 42406 178848 42458
rect 1104 42384 178848 42406
rect 1104 41914 178848 41936
rect 1104 41862 19606 41914
rect 19658 41862 19670 41914
rect 19722 41862 19734 41914
rect 19786 41862 19798 41914
rect 19850 41862 50326 41914
rect 50378 41862 50390 41914
rect 50442 41862 50454 41914
rect 50506 41862 50518 41914
rect 50570 41862 81046 41914
rect 81098 41862 81110 41914
rect 81162 41862 81174 41914
rect 81226 41862 81238 41914
rect 81290 41862 111766 41914
rect 111818 41862 111830 41914
rect 111882 41862 111894 41914
rect 111946 41862 111958 41914
rect 112010 41862 142486 41914
rect 142538 41862 142550 41914
rect 142602 41862 142614 41914
rect 142666 41862 142678 41914
rect 142730 41862 173206 41914
rect 173258 41862 173270 41914
rect 173322 41862 173334 41914
rect 173386 41862 173398 41914
rect 173450 41862 178848 41914
rect 1104 41840 178848 41862
rect 1104 41370 178848 41392
rect 1104 41318 4246 41370
rect 4298 41318 4310 41370
rect 4362 41318 4374 41370
rect 4426 41318 4438 41370
rect 4490 41318 34966 41370
rect 35018 41318 35030 41370
rect 35082 41318 35094 41370
rect 35146 41318 35158 41370
rect 35210 41318 65686 41370
rect 65738 41318 65750 41370
rect 65802 41318 65814 41370
rect 65866 41318 65878 41370
rect 65930 41318 96406 41370
rect 96458 41318 96470 41370
rect 96522 41318 96534 41370
rect 96586 41318 96598 41370
rect 96650 41318 127126 41370
rect 127178 41318 127190 41370
rect 127242 41318 127254 41370
rect 127306 41318 127318 41370
rect 127370 41318 157846 41370
rect 157898 41318 157910 41370
rect 157962 41318 157974 41370
rect 158026 41318 158038 41370
rect 158090 41318 178848 41370
rect 1104 41296 178848 41318
rect 1104 40826 178848 40848
rect 1104 40774 19606 40826
rect 19658 40774 19670 40826
rect 19722 40774 19734 40826
rect 19786 40774 19798 40826
rect 19850 40774 50326 40826
rect 50378 40774 50390 40826
rect 50442 40774 50454 40826
rect 50506 40774 50518 40826
rect 50570 40774 81046 40826
rect 81098 40774 81110 40826
rect 81162 40774 81174 40826
rect 81226 40774 81238 40826
rect 81290 40774 111766 40826
rect 111818 40774 111830 40826
rect 111882 40774 111894 40826
rect 111946 40774 111958 40826
rect 112010 40774 142486 40826
rect 142538 40774 142550 40826
rect 142602 40774 142614 40826
rect 142666 40774 142678 40826
rect 142730 40774 173206 40826
rect 173258 40774 173270 40826
rect 173322 40774 173334 40826
rect 173386 40774 173398 40826
rect 173450 40774 178848 40826
rect 1104 40752 178848 40774
rect 1104 40282 178848 40304
rect 1104 40230 4246 40282
rect 4298 40230 4310 40282
rect 4362 40230 4374 40282
rect 4426 40230 4438 40282
rect 4490 40230 34966 40282
rect 35018 40230 35030 40282
rect 35082 40230 35094 40282
rect 35146 40230 35158 40282
rect 35210 40230 65686 40282
rect 65738 40230 65750 40282
rect 65802 40230 65814 40282
rect 65866 40230 65878 40282
rect 65930 40230 96406 40282
rect 96458 40230 96470 40282
rect 96522 40230 96534 40282
rect 96586 40230 96598 40282
rect 96650 40230 127126 40282
rect 127178 40230 127190 40282
rect 127242 40230 127254 40282
rect 127306 40230 127318 40282
rect 127370 40230 157846 40282
rect 157898 40230 157910 40282
rect 157962 40230 157974 40282
rect 158026 40230 158038 40282
rect 158090 40230 178848 40282
rect 1104 40208 178848 40230
rect 1104 39738 178848 39760
rect 1104 39686 19606 39738
rect 19658 39686 19670 39738
rect 19722 39686 19734 39738
rect 19786 39686 19798 39738
rect 19850 39686 50326 39738
rect 50378 39686 50390 39738
rect 50442 39686 50454 39738
rect 50506 39686 50518 39738
rect 50570 39686 81046 39738
rect 81098 39686 81110 39738
rect 81162 39686 81174 39738
rect 81226 39686 81238 39738
rect 81290 39686 111766 39738
rect 111818 39686 111830 39738
rect 111882 39686 111894 39738
rect 111946 39686 111958 39738
rect 112010 39686 142486 39738
rect 142538 39686 142550 39738
rect 142602 39686 142614 39738
rect 142666 39686 142678 39738
rect 142730 39686 173206 39738
rect 173258 39686 173270 39738
rect 173322 39686 173334 39738
rect 173386 39686 173398 39738
rect 173450 39686 178848 39738
rect 1104 39664 178848 39686
rect 1104 39194 178848 39216
rect 1104 39142 4246 39194
rect 4298 39142 4310 39194
rect 4362 39142 4374 39194
rect 4426 39142 4438 39194
rect 4490 39142 34966 39194
rect 35018 39142 35030 39194
rect 35082 39142 35094 39194
rect 35146 39142 35158 39194
rect 35210 39142 65686 39194
rect 65738 39142 65750 39194
rect 65802 39142 65814 39194
rect 65866 39142 65878 39194
rect 65930 39142 96406 39194
rect 96458 39142 96470 39194
rect 96522 39142 96534 39194
rect 96586 39142 96598 39194
rect 96650 39142 127126 39194
rect 127178 39142 127190 39194
rect 127242 39142 127254 39194
rect 127306 39142 127318 39194
rect 127370 39142 157846 39194
rect 157898 39142 157910 39194
rect 157962 39142 157974 39194
rect 158026 39142 158038 39194
rect 158090 39142 178848 39194
rect 1104 39120 178848 39142
rect 1104 38650 178848 38672
rect 1104 38598 19606 38650
rect 19658 38598 19670 38650
rect 19722 38598 19734 38650
rect 19786 38598 19798 38650
rect 19850 38598 50326 38650
rect 50378 38598 50390 38650
rect 50442 38598 50454 38650
rect 50506 38598 50518 38650
rect 50570 38598 81046 38650
rect 81098 38598 81110 38650
rect 81162 38598 81174 38650
rect 81226 38598 81238 38650
rect 81290 38598 111766 38650
rect 111818 38598 111830 38650
rect 111882 38598 111894 38650
rect 111946 38598 111958 38650
rect 112010 38598 142486 38650
rect 142538 38598 142550 38650
rect 142602 38598 142614 38650
rect 142666 38598 142678 38650
rect 142730 38598 173206 38650
rect 173258 38598 173270 38650
rect 173322 38598 173334 38650
rect 173386 38598 173398 38650
rect 173450 38598 178848 38650
rect 1104 38576 178848 38598
rect 1104 38106 178848 38128
rect 1104 38054 4246 38106
rect 4298 38054 4310 38106
rect 4362 38054 4374 38106
rect 4426 38054 4438 38106
rect 4490 38054 34966 38106
rect 35018 38054 35030 38106
rect 35082 38054 35094 38106
rect 35146 38054 35158 38106
rect 35210 38054 65686 38106
rect 65738 38054 65750 38106
rect 65802 38054 65814 38106
rect 65866 38054 65878 38106
rect 65930 38054 96406 38106
rect 96458 38054 96470 38106
rect 96522 38054 96534 38106
rect 96586 38054 96598 38106
rect 96650 38054 127126 38106
rect 127178 38054 127190 38106
rect 127242 38054 127254 38106
rect 127306 38054 127318 38106
rect 127370 38054 157846 38106
rect 157898 38054 157910 38106
rect 157962 38054 157974 38106
rect 158026 38054 158038 38106
rect 158090 38054 178848 38106
rect 1104 38032 178848 38054
rect 1104 37562 178848 37584
rect 1104 37510 19606 37562
rect 19658 37510 19670 37562
rect 19722 37510 19734 37562
rect 19786 37510 19798 37562
rect 19850 37510 50326 37562
rect 50378 37510 50390 37562
rect 50442 37510 50454 37562
rect 50506 37510 50518 37562
rect 50570 37510 81046 37562
rect 81098 37510 81110 37562
rect 81162 37510 81174 37562
rect 81226 37510 81238 37562
rect 81290 37510 111766 37562
rect 111818 37510 111830 37562
rect 111882 37510 111894 37562
rect 111946 37510 111958 37562
rect 112010 37510 142486 37562
rect 142538 37510 142550 37562
rect 142602 37510 142614 37562
rect 142666 37510 142678 37562
rect 142730 37510 173206 37562
rect 173258 37510 173270 37562
rect 173322 37510 173334 37562
rect 173386 37510 173398 37562
rect 173450 37510 178848 37562
rect 1104 37488 178848 37510
rect 1104 37018 178848 37040
rect 1104 36966 4246 37018
rect 4298 36966 4310 37018
rect 4362 36966 4374 37018
rect 4426 36966 4438 37018
rect 4490 36966 34966 37018
rect 35018 36966 35030 37018
rect 35082 36966 35094 37018
rect 35146 36966 35158 37018
rect 35210 36966 65686 37018
rect 65738 36966 65750 37018
rect 65802 36966 65814 37018
rect 65866 36966 65878 37018
rect 65930 36966 96406 37018
rect 96458 36966 96470 37018
rect 96522 36966 96534 37018
rect 96586 36966 96598 37018
rect 96650 36966 127126 37018
rect 127178 36966 127190 37018
rect 127242 36966 127254 37018
rect 127306 36966 127318 37018
rect 127370 36966 157846 37018
rect 157898 36966 157910 37018
rect 157962 36966 157974 37018
rect 158026 36966 158038 37018
rect 158090 36966 178848 37018
rect 1104 36944 178848 36966
rect 1104 36474 178848 36496
rect 1104 36422 19606 36474
rect 19658 36422 19670 36474
rect 19722 36422 19734 36474
rect 19786 36422 19798 36474
rect 19850 36422 50326 36474
rect 50378 36422 50390 36474
rect 50442 36422 50454 36474
rect 50506 36422 50518 36474
rect 50570 36422 81046 36474
rect 81098 36422 81110 36474
rect 81162 36422 81174 36474
rect 81226 36422 81238 36474
rect 81290 36422 111766 36474
rect 111818 36422 111830 36474
rect 111882 36422 111894 36474
rect 111946 36422 111958 36474
rect 112010 36422 142486 36474
rect 142538 36422 142550 36474
rect 142602 36422 142614 36474
rect 142666 36422 142678 36474
rect 142730 36422 173206 36474
rect 173258 36422 173270 36474
rect 173322 36422 173334 36474
rect 173386 36422 173398 36474
rect 173450 36422 178848 36474
rect 1104 36400 178848 36422
rect 1104 35930 178848 35952
rect 1104 35878 4246 35930
rect 4298 35878 4310 35930
rect 4362 35878 4374 35930
rect 4426 35878 4438 35930
rect 4490 35878 34966 35930
rect 35018 35878 35030 35930
rect 35082 35878 35094 35930
rect 35146 35878 35158 35930
rect 35210 35878 65686 35930
rect 65738 35878 65750 35930
rect 65802 35878 65814 35930
rect 65866 35878 65878 35930
rect 65930 35878 96406 35930
rect 96458 35878 96470 35930
rect 96522 35878 96534 35930
rect 96586 35878 96598 35930
rect 96650 35878 127126 35930
rect 127178 35878 127190 35930
rect 127242 35878 127254 35930
rect 127306 35878 127318 35930
rect 127370 35878 157846 35930
rect 157898 35878 157910 35930
rect 157962 35878 157974 35930
rect 158026 35878 158038 35930
rect 158090 35878 178848 35930
rect 1104 35856 178848 35878
rect 1104 35386 178848 35408
rect 1104 35334 19606 35386
rect 19658 35334 19670 35386
rect 19722 35334 19734 35386
rect 19786 35334 19798 35386
rect 19850 35334 50326 35386
rect 50378 35334 50390 35386
rect 50442 35334 50454 35386
rect 50506 35334 50518 35386
rect 50570 35334 81046 35386
rect 81098 35334 81110 35386
rect 81162 35334 81174 35386
rect 81226 35334 81238 35386
rect 81290 35334 111766 35386
rect 111818 35334 111830 35386
rect 111882 35334 111894 35386
rect 111946 35334 111958 35386
rect 112010 35334 142486 35386
rect 142538 35334 142550 35386
rect 142602 35334 142614 35386
rect 142666 35334 142678 35386
rect 142730 35334 173206 35386
rect 173258 35334 173270 35386
rect 173322 35334 173334 35386
rect 173386 35334 173398 35386
rect 173450 35334 178848 35386
rect 1104 35312 178848 35334
rect 1104 34842 178848 34864
rect 1104 34790 4246 34842
rect 4298 34790 4310 34842
rect 4362 34790 4374 34842
rect 4426 34790 4438 34842
rect 4490 34790 34966 34842
rect 35018 34790 35030 34842
rect 35082 34790 35094 34842
rect 35146 34790 35158 34842
rect 35210 34790 65686 34842
rect 65738 34790 65750 34842
rect 65802 34790 65814 34842
rect 65866 34790 65878 34842
rect 65930 34790 96406 34842
rect 96458 34790 96470 34842
rect 96522 34790 96534 34842
rect 96586 34790 96598 34842
rect 96650 34790 127126 34842
rect 127178 34790 127190 34842
rect 127242 34790 127254 34842
rect 127306 34790 127318 34842
rect 127370 34790 157846 34842
rect 157898 34790 157910 34842
rect 157962 34790 157974 34842
rect 158026 34790 158038 34842
rect 158090 34790 178848 34842
rect 1104 34768 178848 34790
rect 1104 34298 178848 34320
rect 1104 34246 19606 34298
rect 19658 34246 19670 34298
rect 19722 34246 19734 34298
rect 19786 34246 19798 34298
rect 19850 34246 50326 34298
rect 50378 34246 50390 34298
rect 50442 34246 50454 34298
rect 50506 34246 50518 34298
rect 50570 34246 81046 34298
rect 81098 34246 81110 34298
rect 81162 34246 81174 34298
rect 81226 34246 81238 34298
rect 81290 34246 111766 34298
rect 111818 34246 111830 34298
rect 111882 34246 111894 34298
rect 111946 34246 111958 34298
rect 112010 34246 142486 34298
rect 142538 34246 142550 34298
rect 142602 34246 142614 34298
rect 142666 34246 142678 34298
rect 142730 34246 173206 34298
rect 173258 34246 173270 34298
rect 173322 34246 173334 34298
rect 173386 34246 173398 34298
rect 173450 34246 178848 34298
rect 1104 34224 178848 34246
rect 1104 33754 178848 33776
rect 1104 33702 4246 33754
rect 4298 33702 4310 33754
rect 4362 33702 4374 33754
rect 4426 33702 4438 33754
rect 4490 33702 34966 33754
rect 35018 33702 35030 33754
rect 35082 33702 35094 33754
rect 35146 33702 35158 33754
rect 35210 33702 65686 33754
rect 65738 33702 65750 33754
rect 65802 33702 65814 33754
rect 65866 33702 65878 33754
rect 65930 33702 96406 33754
rect 96458 33702 96470 33754
rect 96522 33702 96534 33754
rect 96586 33702 96598 33754
rect 96650 33702 127126 33754
rect 127178 33702 127190 33754
rect 127242 33702 127254 33754
rect 127306 33702 127318 33754
rect 127370 33702 157846 33754
rect 157898 33702 157910 33754
rect 157962 33702 157974 33754
rect 158026 33702 158038 33754
rect 158090 33702 178848 33754
rect 1104 33680 178848 33702
rect 1104 33210 178848 33232
rect 1104 33158 19606 33210
rect 19658 33158 19670 33210
rect 19722 33158 19734 33210
rect 19786 33158 19798 33210
rect 19850 33158 50326 33210
rect 50378 33158 50390 33210
rect 50442 33158 50454 33210
rect 50506 33158 50518 33210
rect 50570 33158 81046 33210
rect 81098 33158 81110 33210
rect 81162 33158 81174 33210
rect 81226 33158 81238 33210
rect 81290 33158 111766 33210
rect 111818 33158 111830 33210
rect 111882 33158 111894 33210
rect 111946 33158 111958 33210
rect 112010 33158 142486 33210
rect 142538 33158 142550 33210
rect 142602 33158 142614 33210
rect 142666 33158 142678 33210
rect 142730 33158 173206 33210
rect 173258 33158 173270 33210
rect 173322 33158 173334 33210
rect 173386 33158 173398 33210
rect 173450 33158 178848 33210
rect 1104 33136 178848 33158
rect 1104 32666 178848 32688
rect 1104 32614 4246 32666
rect 4298 32614 4310 32666
rect 4362 32614 4374 32666
rect 4426 32614 4438 32666
rect 4490 32614 34966 32666
rect 35018 32614 35030 32666
rect 35082 32614 35094 32666
rect 35146 32614 35158 32666
rect 35210 32614 65686 32666
rect 65738 32614 65750 32666
rect 65802 32614 65814 32666
rect 65866 32614 65878 32666
rect 65930 32614 96406 32666
rect 96458 32614 96470 32666
rect 96522 32614 96534 32666
rect 96586 32614 96598 32666
rect 96650 32614 127126 32666
rect 127178 32614 127190 32666
rect 127242 32614 127254 32666
rect 127306 32614 127318 32666
rect 127370 32614 157846 32666
rect 157898 32614 157910 32666
rect 157962 32614 157974 32666
rect 158026 32614 158038 32666
rect 158090 32614 178848 32666
rect 1104 32592 178848 32614
rect 1104 32122 178848 32144
rect 1104 32070 19606 32122
rect 19658 32070 19670 32122
rect 19722 32070 19734 32122
rect 19786 32070 19798 32122
rect 19850 32070 50326 32122
rect 50378 32070 50390 32122
rect 50442 32070 50454 32122
rect 50506 32070 50518 32122
rect 50570 32070 81046 32122
rect 81098 32070 81110 32122
rect 81162 32070 81174 32122
rect 81226 32070 81238 32122
rect 81290 32070 111766 32122
rect 111818 32070 111830 32122
rect 111882 32070 111894 32122
rect 111946 32070 111958 32122
rect 112010 32070 142486 32122
rect 142538 32070 142550 32122
rect 142602 32070 142614 32122
rect 142666 32070 142678 32122
rect 142730 32070 173206 32122
rect 173258 32070 173270 32122
rect 173322 32070 173334 32122
rect 173386 32070 173398 32122
rect 173450 32070 178848 32122
rect 1104 32048 178848 32070
rect 1104 31578 178848 31600
rect 1104 31526 4246 31578
rect 4298 31526 4310 31578
rect 4362 31526 4374 31578
rect 4426 31526 4438 31578
rect 4490 31526 34966 31578
rect 35018 31526 35030 31578
rect 35082 31526 35094 31578
rect 35146 31526 35158 31578
rect 35210 31526 65686 31578
rect 65738 31526 65750 31578
rect 65802 31526 65814 31578
rect 65866 31526 65878 31578
rect 65930 31526 96406 31578
rect 96458 31526 96470 31578
rect 96522 31526 96534 31578
rect 96586 31526 96598 31578
rect 96650 31526 127126 31578
rect 127178 31526 127190 31578
rect 127242 31526 127254 31578
rect 127306 31526 127318 31578
rect 127370 31526 157846 31578
rect 157898 31526 157910 31578
rect 157962 31526 157974 31578
rect 158026 31526 158038 31578
rect 158090 31526 178848 31578
rect 1104 31504 178848 31526
rect 1104 31034 178848 31056
rect 1104 30982 19606 31034
rect 19658 30982 19670 31034
rect 19722 30982 19734 31034
rect 19786 30982 19798 31034
rect 19850 30982 50326 31034
rect 50378 30982 50390 31034
rect 50442 30982 50454 31034
rect 50506 30982 50518 31034
rect 50570 30982 81046 31034
rect 81098 30982 81110 31034
rect 81162 30982 81174 31034
rect 81226 30982 81238 31034
rect 81290 30982 111766 31034
rect 111818 30982 111830 31034
rect 111882 30982 111894 31034
rect 111946 30982 111958 31034
rect 112010 30982 142486 31034
rect 142538 30982 142550 31034
rect 142602 30982 142614 31034
rect 142666 30982 142678 31034
rect 142730 30982 173206 31034
rect 173258 30982 173270 31034
rect 173322 30982 173334 31034
rect 173386 30982 173398 31034
rect 173450 30982 178848 31034
rect 1104 30960 178848 30982
rect 1104 30490 178848 30512
rect 1104 30438 4246 30490
rect 4298 30438 4310 30490
rect 4362 30438 4374 30490
rect 4426 30438 4438 30490
rect 4490 30438 34966 30490
rect 35018 30438 35030 30490
rect 35082 30438 35094 30490
rect 35146 30438 35158 30490
rect 35210 30438 65686 30490
rect 65738 30438 65750 30490
rect 65802 30438 65814 30490
rect 65866 30438 65878 30490
rect 65930 30438 96406 30490
rect 96458 30438 96470 30490
rect 96522 30438 96534 30490
rect 96586 30438 96598 30490
rect 96650 30438 127126 30490
rect 127178 30438 127190 30490
rect 127242 30438 127254 30490
rect 127306 30438 127318 30490
rect 127370 30438 157846 30490
rect 157898 30438 157910 30490
rect 157962 30438 157974 30490
rect 158026 30438 158038 30490
rect 158090 30438 178848 30490
rect 1104 30416 178848 30438
rect 1104 29946 178848 29968
rect 1104 29894 19606 29946
rect 19658 29894 19670 29946
rect 19722 29894 19734 29946
rect 19786 29894 19798 29946
rect 19850 29894 50326 29946
rect 50378 29894 50390 29946
rect 50442 29894 50454 29946
rect 50506 29894 50518 29946
rect 50570 29894 81046 29946
rect 81098 29894 81110 29946
rect 81162 29894 81174 29946
rect 81226 29894 81238 29946
rect 81290 29894 111766 29946
rect 111818 29894 111830 29946
rect 111882 29894 111894 29946
rect 111946 29894 111958 29946
rect 112010 29894 142486 29946
rect 142538 29894 142550 29946
rect 142602 29894 142614 29946
rect 142666 29894 142678 29946
rect 142730 29894 173206 29946
rect 173258 29894 173270 29946
rect 173322 29894 173334 29946
rect 173386 29894 173398 29946
rect 173450 29894 178848 29946
rect 1104 29872 178848 29894
rect 1104 29402 178848 29424
rect 1104 29350 4246 29402
rect 4298 29350 4310 29402
rect 4362 29350 4374 29402
rect 4426 29350 4438 29402
rect 4490 29350 34966 29402
rect 35018 29350 35030 29402
rect 35082 29350 35094 29402
rect 35146 29350 35158 29402
rect 35210 29350 65686 29402
rect 65738 29350 65750 29402
rect 65802 29350 65814 29402
rect 65866 29350 65878 29402
rect 65930 29350 96406 29402
rect 96458 29350 96470 29402
rect 96522 29350 96534 29402
rect 96586 29350 96598 29402
rect 96650 29350 127126 29402
rect 127178 29350 127190 29402
rect 127242 29350 127254 29402
rect 127306 29350 127318 29402
rect 127370 29350 157846 29402
rect 157898 29350 157910 29402
rect 157962 29350 157974 29402
rect 158026 29350 158038 29402
rect 158090 29350 178848 29402
rect 1104 29328 178848 29350
rect 1104 28858 178848 28880
rect 1104 28806 19606 28858
rect 19658 28806 19670 28858
rect 19722 28806 19734 28858
rect 19786 28806 19798 28858
rect 19850 28806 50326 28858
rect 50378 28806 50390 28858
rect 50442 28806 50454 28858
rect 50506 28806 50518 28858
rect 50570 28806 81046 28858
rect 81098 28806 81110 28858
rect 81162 28806 81174 28858
rect 81226 28806 81238 28858
rect 81290 28806 111766 28858
rect 111818 28806 111830 28858
rect 111882 28806 111894 28858
rect 111946 28806 111958 28858
rect 112010 28806 142486 28858
rect 142538 28806 142550 28858
rect 142602 28806 142614 28858
rect 142666 28806 142678 28858
rect 142730 28806 173206 28858
rect 173258 28806 173270 28858
rect 173322 28806 173334 28858
rect 173386 28806 173398 28858
rect 173450 28806 178848 28858
rect 1104 28784 178848 28806
rect 1104 28314 178848 28336
rect 1104 28262 4246 28314
rect 4298 28262 4310 28314
rect 4362 28262 4374 28314
rect 4426 28262 4438 28314
rect 4490 28262 34966 28314
rect 35018 28262 35030 28314
rect 35082 28262 35094 28314
rect 35146 28262 35158 28314
rect 35210 28262 65686 28314
rect 65738 28262 65750 28314
rect 65802 28262 65814 28314
rect 65866 28262 65878 28314
rect 65930 28262 96406 28314
rect 96458 28262 96470 28314
rect 96522 28262 96534 28314
rect 96586 28262 96598 28314
rect 96650 28262 127126 28314
rect 127178 28262 127190 28314
rect 127242 28262 127254 28314
rect 127306 28262 127318 28314
rect 127370 28262 157846 28314
rect 157898 28262 157910 28314
rect 157962 28262 157974 28314
rect 158026 28262 158038 28314
rect 158090 28262 178848 28314
rect 1104 28240 178848 28262
rect 1104 27770 178848 27792
rect 1104 27718 19606 27770
rect 19658 27718 19670 27770
rect 19722 27718 19734 27770
rect 19786 27718 19798 27770
rect 19850 27718 50326 27770
rect 50378 27718 50390 27770
rect 50442 27718 50454 27770
rect 50506 27718 50518 27770
rect 50570 27718 81046 27770
rect 81098 27718 81110 27770
rect 81162 27718 81174 27770
rect 81226 27718 81238 27770
rect 81290 27718 111766 27770
rect 111818 27718 111830 27770
rect 111882 27718 111894 27770
rect 111946 27718 111958 27770
rect 112010 27718 142486 27770
rect 142538 27718 142550 27770
rect 142602 27718 142614 27770
rect 142666 27718 142678 27770
rect 142730 27718 173206 27770
rect 173258 27718 173270 27770
rect 173322 27718 173334 27770
rect 173386 27718 173398 27770
rect 173450 27718 178848 27770
rect 1104 27696 178848 27718
rect 1104 27226 178848 27248
rect 1104 27174 4246 27226
rect 4298 27174 4310 27226
rect 4362 27174 4374 27226
rect 4426 27174 4438 27226
rect 4490 27174 34966 27226
rect 35018 27174 35030 27226
rect 35082 27174 35094 27226
rect 35146 27174 35158 27226
rect 35210 27174 65686 27226
rect 65738 27174 65750 27226
rect 65802 27174 65814 27226
rect 65866 27174 65878 27226
rect 65930 27174 96406 27226
rect 96458 27174 96470 27226
rect 96522 27174 96534 27226
rect 96586 27174 96598 27226
rect 96650 27174 127126 27226
rect 127178 27174 127190 27226
rect 127242 27174 127254 27226
rect 127306 27174 127318 27226
rect 127370 27174 157846 27226
rect 157898 27174 157910 27226
rect 157962 27174 157974 27226
rect 158026 27174 158038 27226
rect 158090 27174 178848 27226
rect 1104 27152 178848 27174
rect 1104 26682 178848 26704
rect 1104 26630 19606 26682
rect 19658 26630 19670 26682
rect 19722 26630 19734 26682
rect 19786 26630 19798 26682
rect 19850 26630 50326 26682
rect 50378 26630 50390 26682
rect 50442 26630 50454 26682
rect 50506 26630 50518 26682
rect 50570 26630 81046 26682
rect 81098 26630 81110 26682
rect 81162 26630 81174 26682
rect 81226 26630 81238 26682
rect 81290 26630 111766 26682
rect 111818 26630 111830 26682
rect 111882 26630 111894 26682
rect 111946 26630 111958 26682
rect 112010 26630 142486 26682
rect 142538 26630 142550 26682
rect 142602 26630 142614 26682
rect 142666 26630 142678 26682
rect 142730 26630 173206 26682
rect 173258 26630 173270 26682
rect 173322 26630 173334 26682
rect 173386 26630 173398 26682
rect 173450 26630 178848 26682
rect 1104 26608 178848 26630
rect 1104 26138 178848 26160
rect 1104 26086 4246 26138
rect 4298 26086 4310 26138
rect 4362 26086 4374 26138
rect 4426 26086 4438 26138
rect 4490 26086 34966 26138
rect 35018 26086 35030 26138
rect 35082 26086 35094 26138
rect 35146 26086 35158 26138
rect 35210 26086 65686 26138
rect 65738 26086 65750 26138
rect 65802 26086 65814 26138
rect 65866 26086 65878 26138
rect 65930 26086 96406 26138
rect 96458 26086 96470 26138
rect 96522 26086 96534 26138
rect 96586 26086 96598 26138
rect 96650 26086 127126 26138
rect 127178 26086 127190 26138
rect 127242 26086 127254 26138
rect 127306 26086 127318 26138
rect 127370 26086 157846 26138
rect 157898 26086 157910 26138
rect 157962 26086 157974 26138
rect 158026 26086 158038 26138
rect 158090 26086 178848 26138
rect 1104 26064 178848 26086
rect 1104 25594 178848 25616
rect 1104 25542 19606 25594
rect 19658 25542 19670 25594
rect 19722 25542 19734 25594
rect 19786 25542 19798 25594
rect 19850 25542 50326 25594
rect 50378 25542 50390 25594
rect 50442 25542 50454 25594
rect 50506 25542 50518 25594
rect 50570 25542 81046 25594
rect 81098 25542 81110 25594
rect 81162 25542 81174 25594
rect 81226 25542 81238 25594
rect 81290 25542 111766 25594
rect 111818 25542 111830 25594
rect 111882 25542 111894 25594
rect 111946 25542 111958 25594
rect 112010 25542 142486 25594
rect 142538 25542 142550 25594
rect 142602 25542 142614 25594
rect 142666 25542 142678 25594
rect 142730 25542 173206 25594
rect 173258 25542 173270 25594
rect 173322 25542 173334 25594
rect 173386 25542 173398 25594
rect 173450 25542 178848 25594
rect 1104 25520 178848 25542
rect 1104 25050 178848 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 34966 25050
rect 35018 24998 35030 25050
rect 35082 24998 35094 25050
rect 35146 24998 35158 25050
rect 35210 24998 65686 25050
rect 65738 24998 65750 25050
rect 65802 24998 65814 25050
rect 65866 24998 65878 25050
rect 65930 24998 96406 25050
rect 96458 24998 96470 25050
rect 96522 24998 96534 25050
rect 96586 24998 96598 25050
rect 96650 24998 127126 25050
rect 127178 24998 127190 25050
rect 127242 24998 127254 25050
rect 127306 24998 127318 25050
rect 127370 24998 157846 25050
rect 157898 24998 157910 25050
rect 157962 24998 157974 25050
rect 158026 24998 158038 25050
rect 158090 24998 178848 25050
rect 1104 24976 178848 24998
rect 1104 24506 178848 24528
rect 1104 24454 19606 24506
rect 19658 24454 19670 24506
rect 19722 24454 19734 24506
rect 19786 24454 19798 24506
rect 19850 24454 50326 24506
rect 50378 24454 50390 24506
rect 50442 24454 50454 24506
rect 50506 24454 50518 24506
rect 50570 24454 81046 24506
rect 81098 24454 81110 24506
rect 81162 24454 81174 24506
rect 81226 24454 81238 24506
rect 81290 24454 111766 24506
rect 111818 24454 111830 24506
rect 111882 24454 111894 24506
rect 111946 24454 111958 24506
rect 112010 24454 142486 24506
rect 142538 24454 142550 24506
rect 142602 24454 142614 24506
rect 142666 24454 142678 24506
rect 142730 24454 173206 24506
rect 173258 24454 173270 24506
rect 173322 24454 173334 24506
rect 173386 24454 173398 24506
rect 173450 24454 178848 24506
rect 1104 24432 178848 24454
rect 31018 24216 31024 24268
rect 31076 24256 31082 24268
rect 31386 24256 31392 24268
rect 31076 24228 31392 24256
rect 31076 24216 31082 24228
rect 31386 24216 31392 24228
rect 31444 24256 31450 24268
rect 32769 24259 32827 24265
rect 32769 24256 32781 24259
rect 31444 24228 32781 24256
rect 31444 24216 31450 24228
rect 32769 24225 32781 24228
rect 32815 24225 32827 24259
rect 32769 24219 32827 24225
rect 32953 24259 33011 24265
rect 32953 24225 32965 24259
rect 32999 24256 33011 24259
rect 35894 24256 35900 24268
rect 32999 24228 35900 24256
rect 32999 24225 33011 24228
rect 32953 24219 33011 24225
rect 35894 24216 35900 24228
rect 35952 24256 35958 24268
rect 36814 24256 36820 24268
rect 35952 24228 36820 24256
rect 35952 24216 35958 24228
rect 36814 24216 36820 24228
rect 36872 24216 36878 24268
rect 32861 24055 32919 24061
rect 32861 24021 32873 24055
rect 32907 24052 32919 24055
rect 33134 24052 33140 24064
rect 32907 24024 33140 24052
rect 32907 24021 32919 24024
rect 32861 24015 32919 24021
rect 33134 24012 33140 24024
rect 33192 24012 33198 24064
rect 1104 23962 178848 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 34966 23962
rect 35018 23910 35030 23962
rect 35082 23910 35094 23962
rect 35146 23910 35158 23962
rect 35210 23910 65686 23962
rect 65738 23910 65750 23962
rect 65802 23910 65814 23962
rect 65866 23910 65878 23962
rect 65930 23910 96406 23962
rect 96458 23910 96470 23962
rect 96522 23910 96534 23962
rect 96586 23910 96598 23962
rect 96650 23910 127126 23962
rect 127178 23910 127190 23962
rect 127242 23910 127254 23962
rect 127306 23910 127318 23962
rect 127370 23910 157846 23962
rect 157898 23910 157910 23962
rect 157962 23910 157974 23962
rect 158026 23910 158038 23962
rect 158090 23910 178848 23962
rect 1104 23888 178848 23910
rect 1104 23418 178848 23440
rect 1104 23366 19606 23418
rect 19658 23366 19670 23418
rect 19722 23366 19734 23418
rect 19786 23366 19798 23418
rect 19850 23366 50326 23418
rect 50378 23366 50390 23418
rect 50442 23366 50454 23418
rect 50506 23366 50518 23418
rect 50570 23366 81046 23418
rect 81098 23366 81110 23418
rect 81162 23366 81174 23418
rect 81226 23366 81238 23418
rect 81290 23366 111766 23418
rect 111818 23366 111830 23418
rect 111882 23366 111894 23418
rect 111946 23366 111958 23418
rect 112010 23366 142486 23418
rect 142538 23366 142550 23418
rect 142602 23366 142614 23418
rect 142666 23366 142678 23418
rect 142730 23366 173206 23418
rect 173258 23366 173270 23418
rect 173322 23366 173334 23418
rect 173386 23366 173398 23418
rect 173450 23366 178848 23418
rect 1104 23344 178848 23366
rect 26418 23168 26424 23180
rect 26331 23140 26424 23168
rect 26418 23128 26424 23140
rect 26476 23128 26482 23180
rect 26602 23168 26608 23180
rect 26515 23140 26608 23168
rect 26602 23128 26608 23140
rect 26660 23168 26666 23180
rect 28258 23168 28264 23180
rect 26660 23140 28264 23168
rect 26660 23128 26666 23140
rect 28258 23128 28264 23140
rect 28316 23128 28322 23180
rect 26436 23100 26464 23128
rect 28166 23100 28172 23112
rect 26436 23072 28172 23100
rect 28166 23060 28172 23072
rect 28224 23060 28230 23112
rect 26513 22967 26571 22973
rect 26513 22933 26525 22967
rect 26559 22964 26571 22967
rect 27982 22964 27988 22976
rect 26559 22936 27988 22964
rect 26559 22933 26571 22936
rect 26513 22927 26571 22933
rect 27982 22924 27988 22936
rect 28040 22924 28046 22976
rect 1104 22874 178848 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 34966 22874
rect 35018 22822 35030 22874
rect 35082 22822 35094 22874
rect 35146 22822 35158 22874
rect 35210 22822 65686 22874
rect 65738 22822 65750 22874
rect 65802 22822 65814 22874
rect 65866 22822 65878 22874
rect 65930 22822 96406 22874
rect 96458 22822 96470 22874
rect 96522 22822 96534 22874
rect 96586 22822 96598 22874
rect 96650 22822 127126 22874
rect 127178 22822 127190 22874
rect 127242 22822 127254 22874
rect 127306 22822 127318 22874
rect 127370 22822 157846 22874
rect 157898 22822 157910 22874
rect 157962 22822 157974 22874
rect 158026 22822 158038 22874
rect 158090 22822 178848 22874
rect 1104 22800 178848 22822
rect 33134 22624 33140 22636
rect 33095 22596 33140 22624
rect 33134 22584 33140 22596
rect 33192 22584 33198 22636
rect 32122 22516 32128 22568
rect 32180 22556 32186 22568
rect 33505 22559 33563 22565
rect 33505 22556 33517 22559
rect 32180 22528 33517 22556
rect 32180 22516 32186 22528
rect 33505 22525 33517 22528
rect 33551 22525 33563 22559
rect 33505 22519 33563 22525
rect 30374 22448 30380 22500
rect 30432 22488 30438 22500
rect 33622 22491 33680 22497
rect 33622 22488 33634 22491
rect 30432 22460 33634 22488
rect 30432 22448 30438 22460
rect 33622 22457 33634 22460
rect 33668 22457 33680 22491
rect 33622 22451 33680 22457
rect 33410 22420 33416 22432
rect 33371 22392 33416 22420
rect 33410 22380 33416 22392
rect 33468 22380 33474 22432
rect 33781 22423 33839 22429
rect 33781 22389 33793 22423
rect 33827 22420 33839 22423
rect 35250 22420 35256 22432
rect 33827 22392 35256 22420
rect 33827 22389 33839 22392
rect 33781 22383 33839 22389
rect 35250 22380 35256 22392
rect 35308 22380 35314 22432
rect 1104 22330 178848 22352
rect 1104 22278 19606 22330
rect 19658 22278 19670 22330
rect 19722 22278 19734 22330
rect 19786 22278 19798 22330
rect 19850 22278 50326 22330
rect 50378 22278 50390 22330
rect 50442 22278 50454 22330
rect 50506 22278 50518 22330
rect 50570 22278 81046 22330
rect 81098 22278 81110 22330
rect 81162 22278 81174 22330
rect 81226 22278 81238 22330
rect 81290 22278 111766 22330
rect 111818 22278 111830 22330
rect 111882 22278 111894 22330
rect 111946 22278 111958 22330
rect 112010 22278 142486 22330
rect 142538 22278 142550 22330
rect 142602 22278 142614 22330
rect 142666 22278 142678 22330
rect 142730 22278 173206 22330
rect 173258 22278 173270 22330
rect 173322 22278 173334 22330
rect 173386 22278 173398 22330
rect 173450 22278 178848 22330
rect 1104 22256 178848 22278
rect 29086 22148 29092 22160
rect 29047 22120 29092 22148
rect 29086 22108 29092 22120
rect 29144 22108 29150 22160
rect 29270 22108 29276 22160
rect 29328 22157 29334 22160
rect 29328 22151 29352 22157
rect 29340 22117 29352 22151
rect 29328 22111 29352 22117
rect 29328 22108 29334 22111
rect 29457 21947 29515 21953
rect 29457 21913 29469 21947
rect 29503 21944 29515 21947
rect 30374 21944 30380 21956
rect 29503 21916 30380 21944
rect 29503 21913 29515 21916
rect 29457 21907 29515 21913
rect 30374 21904 30380 21916
rect 30432 21904 30438 21956
rect 29178 21836 29184 21888
rect 29236 21876 29242 21888
rect 29273 21879 29331 21885
rect 29273 21876 29285 21879
rect 29236 21848 29285 21876
rect 29236 21836 29242 21848
rect 29273 21845 29285 21848
rect 29319 21845 29331 21879
rect 29273 21839 29331 21845
rect 1104 21786 178848 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 34966 21786
rect 35018 21734 35030 21786
rect 35082 21734 35094 21786
rect 35146 21734 35158 21786
rect 35210 21734 65686 21786
rect 65738 21734 65750 21786
rect 65802 21734 65814 21786
rect 65866 21734 65878 21786
rect 65930 21734 96406 21786
rect 96458 21734 96470 21786
rect 96522 21734 96534 21786
rect 96586 21734 96598 21786
rect 96650 21734 127126 21786
rect 127178 21734 127190 21786
rect 127242 21734 127254 21786
rect 127306 21734 127318 21786
rect 127370 21734 157846 21786
rect 157898 21734 157910 21786
rect 157962 21734 157974 21786
rect 158026 21734 158038 21786
rect 158090 21734 178848 21786
rect 1104 21712 178848 21734
rect 27982 21468 27988 21480
rect 27943 21440 27988 21468
rect 27982 21428 27988 21440
rect 28040 21428 28046 21480
rect 28077 21335 28135 21341
rect 28077 21301 28089 21335
rect 28123 21332 28135 21335
rect 29270 21332 29276 21344
rect 28123 21304 29276 21332
rect 28123 21301 28135 21304
rect 28077 21295 28135 21301
rect 29270 21292 29276 21304
rect 29328 21292 29334 21344
rect 1104 21242 178848 21264
rect 1104 21190 19606 21242
rect 19658 21190 19670 21242
rect 19722 21190 19734 21242
rect 19786 21190 19798 21242
rect 19850 21190 50326 21242
rect 50378 21190 50390 21242
rect 50442 21190 50454 21242
rect 50506 21190 50518 21242
rect 50570 21190 81046 21242
rect 81098 21190 81110 21242
rect 81162 21190 81174 21242
rect 81226 21190 81238 21242
rect 81290 21190 111766 21242
rect 111818 21190 111830 21242
rect 111882 21190 111894 21242
rect 111946 21190 111958 21242
rect 112010 21190 142486 21242
rect 142538 21190 142550 21242
rect 142602 21190 142614 21242
rect 142666 21190 142678 21242
rect 142730 21190 173206 21242
rect 173258 21190 173270 21242
rect 173322 21190 173334 21242
rect 173386 21190 173398 21242
rect 173450 21190 178848 21242
rect 1104 21168 178848 21190
rect 28997 21063 29055 21069
rect 28997 21029 29009 21063
rect 29043 21060 29055 21063
rect 29086 21060 29092 21072
rect 29043 21032 29092 21060
rect 29043 21029 29055 21032
rect 28997 21023 29055 21029
rect 29086 21020 29092 21032
rect 29144 21060 29150 21072
rect 32030 21060 32036 21072
rect 29144 21032 32036 21060
rect 29144 21020 29150 21032
rect 32030 21020 32036 21032
rect 32088 21020 32094 21072
rect 29178 20992 29184 21004
rect 29139 20964 29184 20992
rect 29178 20952 29184 20964
rect 29236 20952 29242 21004
rect 29270 20952 29276 21004
rect 29328 20992 29334 21004
rect 29328 20964 29373 20992
rect 29328 20952 29334 20964
rect 28997 20791 29055 20797
rect 28997 20757 29009 20791
rect 29043 20788 29055 20791
rect 30650 20788 30656 20800
rect 29043 20760 30656 20788
rect 29043 20757 29055 20760
rect 28997 20751 29055 20757
rect 30650 20748 30656 20760
rect 30708 20748 30714 20800
rect 1104 20698 178848 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 34966 20698
rect 35018 20646 35030 20698
rect 35082 20646 35094 20698
rect 35146 20646 35158 20698
rect 35210 20646 65686 20698
rect 65738 20646 65750 20698
rect 65802 20646 65814 20698
rect 65866 20646 65878 20698
rect 65930 20646 96406 20698
rect 96458 20646 96470 20698
rect 96522 20646 96534 20698
rect 96586 20646 96598 20698
rect 96650 20646 127126 20698
rect 127178 20646 127190 20698
rect 127242 20646 127254 20698
rect 127306 20646 127318 20698
rect 127370 20646 157846 20698
rect 157898 20646 157910 20698
rect 157962 20646 157974 20698
rect 158026 20646 158038 20698
rect 158090 20646 178848 20698
rect 1104 20624 178848 20646
rect 28166 20448 28172 20460
rect 28079 20420 28172 20448
rect 28166 20408 28172 20420
rect 28224 20448 28230 20460
rect 33226 20448 33232 20460
rect 28224 20420 33232 20448
rect 28224 20408 28230 20420
rect 33226 20408 33232 20420
rect 33284 20408 33290 20460
rect 27982 20380 27988 20392
rect 27943 20352 27988 20380
rect 27982 20340 27988 20352
rect 28040 20340 28046 20392
rect 28258 20340 28264 20392
rect 28316 20380 28322 20392
rect 29086 20380 29092 20392
rect 28316 20352 29092 20380
rect 28316 20340 28322 20352
rect 29086 20340 29092 20352
rect 29144 20340 29150 20392
rect 76101 20383 76159 20389
rect 76101 20380 76113 20383
rect 75748 20352 76113 20380
rect 27801 20247 27859 20253
rect 27801 20213 27813 20247
rect 27847 20244 27859 20247
rect 28994 20244 29000 20256
rect 27847 20216 29000 20244
rect 27847 20213 27859 20216
rect 27801 20207 27859 20213
rect 28994 20204 29000 20216
rect 29052 20204 29058 20256
rect 74534 20204 74540 20256
rect 74592 20244 74598 20256
rect 75748 20253 75776 20352
rect 76101 20349 76113 20352
rect 76147 20380 76159 20383
rect 149514 20380 149520 20392
rect 76147 20352 149520 20380
rect 76147 20349 76159 20352
rect 76101 20343 76159 20349
rect 149514 20340 149520 20352
rect 149572 20340 149578 20392
rect 75733 20247 75791 20253
rect 75733 20244 75745 20247
rect 74592 20216 75745 20244
rect 74592 20204 74598 20216
rect 75733 20213 75745 20216
rect 75779 20213 75791 20247
rect 75733 20207 75791 20213
rect 75822 20204 75828 20256
rect 75880 20244 75886 20256
rect 76009 20247 76067 20253
rect 76009 20244 76021 20247
rect 75880 20216 76021 20244
rect 75880 20204 75886 20216
rect 76009 20213 76021 20216
rect 76055 20213 76067 20247
rect 76009 20207 76067 20213
rect 1104 20154 178848 20176
rect 1104 20102 19606 20154
rect 19658 20102 19670 20154
rect 19722 20102 19734 20154
rect 19786 20102 19798 20154
rect 19850 20102 50326 20154
rect 50378 20102 50390 20154
rect 50442 20102 50454 20154
rect 50506 20102 50518 20154
rect 50570 20102 81046 20154
rect 81098 20102 81110 20154
rect 81162 20102 81174 20154
rect 81226 20102 81238 20154
rect 81290 20102 111766 20154
rect 111818 20102 111830 20154
rect 111882 20102 111894 20154
rect 111946 20102 111958 20154
rect 112010 20102 142486 20154
rect 142538 20102 142550 20154
rect 142602 20102 142614 20154
rect 142666 20102 142678 20154
rect 142730 20102 173206 20154
rect 173258 20102 173270 20154
rect 173322 20102 173334 20154
rect 173386 20102 173398 20154
rect 173450 20102 178848 20154
rect 1104 20080 178848 20102
rect 29089 20043 29147 20049
rect 29089 20009 29101 20043
rect 29135 20040 29147 20043
rect 29270 20040 29276 20052
rect 29135 20012 29276 20040
rect 29135 20009 29147 20012
rect 29089 20003 29147 20009
rect 29270 20000 29276 20012
rect 29328 20040 29334 20052
rect 29328 20012 29500 20040
rect 29328 20000 29334 20012
rect 29086 19907 29144 19913
rect 29086 19873 29098 19907
rect 29132 19904 29144 19907
rect 29178 19904 29184 19916
rect 29132 19876 29184 19904
rect 29132 19873 29144 19876
rect 29086 19867 29144 19873
rect 29178 19864 29184 19876
rect 29236 19904 29242 19916
rect 29472 19913 29500 20012
rect 72142 20000 72148 20052
rect 72200 20040 72206 20052
rect 121730 20040 121736 20052
rect 72200 20012 121736 20040
rect 72200 20000 72206 20012
rect 121730 20000 121736 20012
rect 121788 20000 121794 20052
rect 73246 19932 73252 19984
rect 73304 19972 73310 19984
rect 130746 19972 130752 19984
rect 73304 19944 130752 19972
rect 73304 19932 73310 19944
rect 130746 19932 130752 19944
rect 130804 19932 130810 19984
rect 29457 19907 29515 19913
rect 29236 19876 29408 19904
rect 29236 19864 29242 19876
rect 29380 19836 29408 19876
rect 29457 19873 29469 19907
rect 29503 19873 29515 19907
rect 29457 19867 29515 19873
rect 30374 19864 30380 19916
rect 30432 19904 30438 19916
rect 31202 19904 31208 19916
rect 30432 19876 31208 19904
rect 30432 19864 30438 19876
rect 31202 19864 31208 19876
rect 31260 19864 31266 19916
rect 31386 19904 31392 19916
rect 31347 19876 31392 19904
rect 31386 19864 31392 19876
rect 31444 19904 31450 19916
rect 31938 19904 31944 19916
rect 31444 19876 31944 19904
rect 31444 19864 31450 19876
rect 31938 19864 31944 19876
rect 31996 19864 32002 19916
rect 29549 19839 29607 19845
rect 29549 19836 29561 19839
rect 29380 19808 29561 19836
rect 29549 19805 29561 19808
rect 29595 19836 29607 19839
rect 31018 19836 31024 19848
rect 29595 19808 31024 19836
rect 29595 19805 29607 19808
rect 29549 19799 29607 19805
rect 31018 19796 31024 19808
rect 31076 19796 31082 19848
rect 28902 19700 28908 19712
rect 28863 19672 28908 19700
rect 28902 19660 28908 19672
rect 28960 19660 28966 19712
rect 31294 19700 31300 19712
rect 31255 19672 31300 19700
rect 31294 19660 31300 19672
rect 31352 19660 31358 19712
rect 1104 19610 178848 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 34966 19610
rect 35018 19558 35030 19610
rect 35082 19558 35094 19610
rect 35146 19558 35158 19610
rect 35210 19558 65686 19610
rect 65738 19558 65750 19610
rect 65802 19558 65814 19610
rect 65866 19558 65878 19610
rect 65930 19558 96406 19610
rect 96458 19558 96470 19610
rect 96522 19558 96534 19610
rect 96586 19558 96598 19610
rect 96650 19558 127126 19610
rect 127178 19558 127190 19610
rect 127242 19558 127254 19610
rect 127306 19558 127318 19610
rect 127370 19558 157846 19610
rect 157898 19558 157910 19610
rect 157962 19558 157974 19610
rect 158026 19558 158038 19610
rect 158090 19558 178848 19610
rect 1104 19536 178848 19558
rect 74721 19499 74779 19505
rect 74721 19465 74733 19499
rect 74767 19496 74779 19499
rect 75181 19499 75239 19505
rect 75181 19496 75193 19499
rect 74767 19468 75193 19496
rect 74767 19465 74779 19468
rect 74721 19459 74779 19465
rect 75181 19465 75193 19468
rect 75227 19496 75239 19499
rect 135438 19496 135444 19508
rect 75227 19468 135444 19496
rect 75227 19465 75239 19468
rect 75181 19459 75239 19465
rect 135438 19456 135444 19468
rect 135496 19456 135502 19508
rect 35250 19252 35256 19304
rect 35308 19292 35314 19304
rect 35802 19292 35808 19304
rect 35308 19264 35808 19292
rect 35308 19252 35314 19264
rect 35802 19252 35808 19264
rect 35860 19292 35866 19304
rect 37001 19295 37059 19301
rect 37001 19292 37013 19295
rect 35860 19264 37013 19292
rect 35860 19252 35866 19264
rect 37001 19261 37013 19264
rect 37047 19261 37059 19295
rect 37001 19255 37059 19261
rect 37185 19295 37243 19301
rect 37185 19261 37197 19295
rect 37231 19292 37243 19295
rect 37734 19292 37740 19304
rect 37231 19264 37740 19292
rect 37231 19261 37243 19264
rect 37185 19255 37243 19261
rect 37734 19252 37740 19264
rect 37792 19292 37798 19304
rect 41690 19292 41696 19304
rect 37792 19264 41696 19292
rect 37792 19252 37798 19264
rect 41690 19252 41696 19264
rect 41748 19252 41754 19304
rect 57146 19292 57152 19304
rect 57107 19264 57152 19292
rect 57146 19252 57152 19264
rect 57204 19252 57210 19304
rect 58066 19252 58072 19304
rect 58124 19292 58130 19304
rect 59262 19292 59268 19304
rect 58124 19264 59268 19292
rect 58124 19252 58130 19264
rect 59262 19252 59268 19264
rect 59320 19252 59326 19304
rect 60182 19292 60188 19304
rect 60143 19264 60188 19292
rect 60182 19252 60188 19264
rect 60240 19252 60246 19304
rect 61010 19292 61016 19304
rect 60971 19264 61016 19292
rect 61010 19252 61016 19264
rect 61068 19252 61074 19304
rect 65242 19292 65248 19304
rect 65203 19264 65248 19292
rect 65242 19252 65248 19264
rect 65300 19252 65306 19304
rect 72878 19252 72884 19304
rect 72936 19292 72942 19304
rect 73246 19292 73252 19304
rect 72936 19264 73252 19292
rect 72936 19252 72942 19264
rect 73246 19252 73252 19264
rect 73304 19292 73310 19304
rect 73433 19295 73491 19301
rect 73433 19292 73445 19295
rect 73304 19264 73445 19292
rect 73304 19252 73310 19264
rect 73433 19261 73445 19264
rect 73479 19261 73491 19295
rect 73433 19255 73491 19261
rect 75288 19264 75592 19292
rect 75288 19236 75316 19264
rect 71314 19184 71320 19236
rect 71372 19224 71378 19236
rect 73341 19227 73399 19233
rect 73341 19224 73353 19227
rect 71372 19196 73353 19224
rect 71372 19184 71378 19196
rect 73341 19193 73353 19196
rect 73387 19193 73399 19227
rect 75149 19227 75207 19233
rect 75149 19224 75161 19227
rect 73341 19187 73399 19193
rect 73448 19196 75161 19224
rect 37185 19159 37243 19165
rect 37185 19125 37197 19159
rect 37231 19156 37243 19159
rect 37458 19156 37464 19168
rect 37231 19128 37464 19156
rect 37231 19125 37243 19128
rect 37185 19119 37243 19125
rect 37458 19116 37464 19128
rect 37516 19116 37522 19168
rect 42794 19116 42800 19168
rect 42852 19156 42858 19168
rect 43438 19156 43444 19168
rect 42852 19128 43444 19156
rect 42852 19116 42858 19128
rect 43438 19116 43444 19128
rect 43496 19156 43502 19168
rect 50890 19156 50896 19168
rect 43496 19128 50896 19156
rect 43496 19116 43502 19128
rect 50890 19116 50896 19128
rect 50948 19116 50954 19168
rect 57238 19156 57244 19168
rect 57199 19128 57244 19156
rect 57238 19116 57244 19128
rect 57296 19116 57302 19168
rect 59354 19156 59360 19168
rect 59315 19128 59360 19156
rect 59354 19116 59360 19128
rect 59412 19116 59418 19168
rect 60182 19116 60188 19168
rect 60240 19156 60246 19168
rect 60277 19159 60335 19165
rect 60277 19156 60289 19159
rect 60240 19128 60289 19156
rect 60240 19116 60246 19128
rect 60277 19125 60289 19128
rect 60323 19125 60335 19159
rect 61102 19156 61108 19168
rect 61063 19128 61108 19156
rect 60277 19119 60335 19125
rect 61102 19116 61108 19128
rect 61160 19116 61166 19168
rect 65337 19159 65395 19165
rect 65337 19125 65349 19159
rect 65383 19156 65395 19159
rect 65978 19156 65984 19168
rect 65383 19128 65984 19156
rect 65383 19125 65395 19128
rect 65337 19119 65395 19125
rect 65978 19116 65984 19128
rect 66036 19116 66042 19168
rect 68646 19116 68652 19168
rect 68704 19156 68710 19168
rect 72878 19156 72884 19168
rect 68704 19128 72884 19156
rect 68704 19116 68710 19128
rect 72878 19116 72884 19128
rect 72936 19156 72942 19168
rect 73065 19159 73123 19165
rect 73065 19156 73077 19159
rect 72936 19128 73077 19156
rect 72936 19116 72942 19128
rect 73065 19125 73077 19128
rect 73111 19125 73123 19159
rect 73065 19119 73123 19125
rect 73154 19116 73160 19168
rect 73212 19156 73218 19168
rect 73448 19156 73476 19196
rect 75149 19193 75161 19196
rect 75195 19193 75207 19227
rect 75149 19187 75207 19193
rect 75270 19184 75276 19236
rect 75328 19233 75334 19236
rect 75328 19227 75377 19233
rect 75328 19193 75331 19227
rect 75365 19224 75377 19227
rect 75365 19196 75421 19224
rect 75365 19193 75377 19196
rect 75328 19187 75377 19193
rect 75328 19184 75334 19187
rect 73212 19128 73476 19156
rect 73212 19116 73218 19128
rect 73522 19116 73528 19168
rect 73580 19156 73586 19168
rect 74721 19159 74779 19165
rect 74721 19156 74733 19159
rect 73580 19128 74733 19156
rect 73580 19116 73586 19128
rect 74721 19125 74733 19128
rect 74767 19156 74779 19159
rect 74813 19159 74871 19165
rect 74813 19156 74825 19159
rect 74767 19128 74825 19156
rect 74767 19125 74779 19128
rect 74721 19119 74779 19125
rect 74813 19125 74825 19128
rect 74859 19125 74871 19159
rect 74994 19156 75000 19168
rect 74955 19128 75000 19156
rect 74813 19119 74871 19125
rect 74994 19116 75000 19128
rect 75052 19116 75058 19168
rect 75564 19165 75592 19264
rect 75549 19159 75607 19165
rect 75549 19125 75561 19159
rect 75595 19156 75607 19159
rect 140406 19156 140412 19168
rect 75595 19128 140412 19156
rect 75595 19125 75607 19128
rect 75549 19119 75607 19125
rect 140406 19116 140412 19128
rect 140464 19116 140470 19168
rect 1104 19066 178848 19088
rect 1104 19014 19606 19066
rect 19658 19014 19670 19066
rect 19722 19014 19734 19066
rect 19786 19014 19798 19066
rect 19850 19014 50326 19066
rect 50378 19014 50390 19066
rect 50442 19014 50454 19066
rect 50506 19014 50518 19066
rect 50570 19014 81046 19066
rect 81098 19014 81110 19066
rect 81162 19014 81174 19066
rect 81226 19014 81238 19066
rect 81290 19014 111766 19066
rect 111818 19014 111830 19066
rect 111882 19014 111894 19066
rect 111946 19014 111958 19066
rect 112010 19014 142486 19066
rect 142538 19014 142550 19066
rect 142602 19014 142614 19066
rect 142666 19014 142678 19066
rect 142730 19014 173206 19066
rect 173258 19014 173270 19066
rect 173322 19014 173334 19066
rect 173386 19014 173398 19066
rect 173450 19014 178848 19066
rect 1104 18992 178848 19014
rect 44634 18952 44640 18964
rect 44008 18924 44640 18952
rect 31757 18819 31815 18825
rect 31757 18785 31769 18819
rect 31803 18816 31815 18819
rect 33410 18816 33416 18828
rect 31803 18788 33416 18816
rect 31803 18785 31815 18788
rect 31757 18779 31815 18785
rect 33410 18776 33416 18788
rect 33468 18816 33474 18828
rect 35342 18816 35348 18828
rect 33468 18788 35348 18816
rect 33468 18776 33474 18788
rect 35342 18776 35348 18788
rect 35400 18776 35406 18828
rect 42613 18819 42671 18825
rect 42613 18785 42625 18819
rect 42659 18816 42671 18819
rect 42794 18816 42800 18828
rect 42659 18788 42800 18816
rect 42659 18785 42671 18788
rect 42613 18779 42671 18785
rect 42794 18776 42800 18788
rect 42852 18776 42858 18828
rect 44008 18825 44036 18924
rect 44634 18912 44640 18924
rect 44692 18952 44698 18964
rect 44692 18924 55214 18952
rect 44692 18912 44698 18924
rect 46845 18887 46903 18893
rect 46845 18853 46857 18887
rect 46891 18853 46903 18887
rect 46845 18847 46903 18853
rect 43993 18819 44051 18825
rect 43993 18785 44005 18819
rect 44039 18785 44051 18819
rect 43993 18779 44051 18785
rect 31941 18683 31999 18689
rect 31941 18649 31953 18683
rect 31987 18680 31999 18683
rect 32122 18680 32128 18692
rect 31987 18652 32128 18680
rect 31987 18649 31999 18652
rect 31941 18643 31999 18649
rect 32122 18640 32128 18652
rect 32180 18640 32186 18692
rect 46753 18683 46811 18689
rect 46753 18649 46765 18683
rect 46799 18680 46811 18683
rect 46860 18680 46888 18847
rect 46934 18844 46940 18896
rect 46992 18884 46998 18896
rect 47050 18887 47108 18893
rect 47050 18884 47062 18887
rect 46992 18856 47062 18884
rect 46992 18844 46998 18856
rect 47050 18853 47062 18856
rect 47096 18853 47108 18887
rect 47050 18847 47108 18853
rect 55186 18748 55214 18924
rect 73246 18844 73252 18896
rect 73304 18884 73310 18896
rect 74169 18887 74227 18893
rect 74169 18884 74181 18887
rect 73304 18856 74181 18884
rect 73304 18844 73310 18856
rect 74169 18853 74181 18856
rect 74215 18853 74227 18887
rect 74169 18847 74227 18853
rect 66070 18816 66076 18828
rect 66031 18788 66076 18816
rect 66070 18776 66076 18788
rect 66128 18776 66134 18828
rect 67818 18816 67824 18828
rect 67779 18788 67824 18816
rect 67818 18776 67824 18788
rect 67876 18776 67882 18828
rect 68462 18816 68468 18828
rect 68423 18788 68468 18816
rect 68462 18776 68468 18788
rect 68520 18776 68526 18828
rect 72234 18776 72240 18828
rect 72292 18816 72298 18828
rect 72418 18816 72424 18828
rect 72292 18788 72424 18816
rect 72292 18776 72298 18788
rect 72418 18776 72424 18788
rect 72476 18776 72482 18828
rect 72970 18776 72976 18828
rect 73028 18816 73034 18828
rect 73065 18819 73123 18825
rect 73065 18816 73077 18819
rect 73028 18788 73077 18816
rect 73028 18776 73034 18788
rect 73065 18785 73077 18788
rect 73111 18785 73123 18819
rect 73065 18779 73123 18785
rect 74077 18819 74135 18825
rect 74077 18785 74089 18819
rect 74123 18785 74135 18819
rect 74077 18779 74135 18785
rect 55582 18748 55588 18760
rect 55186 18720 55588 18748
rect 55582 18708 55588 18720
rect 55640 18708 55646 18760
rect 47854 18680 47860 18692
rect 46799 18652 47860 18680
rect 46799 18649 46811 18652
rect 46753 18643 46811 18649
rect 47854 18640 47860 18652
rect 47912 18680 47918 18692
rect 65518 18680 65524 18692
rect 47912 18652 65524 18680
rect 47912 18640 47918 18652
rect 65518 18640 65524 18652
rect 65576 18640 65582 18692
rect 67082 18640 67088 18692
rect 67140 18680 67146 18692
rect 68557 18683 68615 18689
rect 68557 18680 68569 18683
rect 67140 18652 68569 18680
rect 67140 18640 67146 18652
rect 68557 18649 68569 18652
rect 68603 18649 68615 18683
rect 68557 18643 68615 18649
rect 71130 18640 71136 18692
rect 71188 18680 71194 18692
rect 73157 18683 73215 18689
rect 73157 18680 73169 18683
rect 71188 18652 73169 18680
rect 71188 18640 71194 18652
rect 73157 18649 73169 18652
rect 73203 18649 73215 18683
rect 73157 18643 73215 18649
rect 42705 18615 42763 18621
rect 42705 18581 42717 18615
rect 42751 18612 42763 18615
rect 42886 18612 42892 18624
rect 42751 18584 42892 18612
rect 42751 18581 42763 18584
rect 42705 18575 42763 18581
rect 42886 18572 42892 18584
rect 42944 18572 42950 18624
rect 44082 18612 44088 18624
rect 44043 18584 44088 18612
rect 44082 18572 44088 18584
rect 44140 18572 44146 18624
rect 47026 18612 47032 18624
rect 46987 18584 47032 18612
rect 47026 18572 47032 18584
rect 47084 18572 47090 18624
rect 47213 18615 47271 18621
rect 47213 18581 47225 18615
rect 47259 18612 47271 18615
rect 48314 18612 48320 18624
rect 47259 18584 48320 18612
rect 47259 18581 47271 18584
rect 47213 18575 47271 18581
rect 48314 18572 48320 18584
rect 48372 18572 48378 18624
rect 66162 18612 66168 18624
rect 66123 18584 66168 18612
rect 66162 18572 66168 18584
rect 66220 18572 66226 18624
rect 66898 18572 66904 18624
rect 66956 18612 66962 18624
rect 67913 18615 67971 18621
rect 67913 18612 67925 18615
rect 66956 18584 67925 18612
rect 66956 18572 66962 18584
rect 67913 18581 67925 18584
rect 67959 18581 67971 18615
rect 67913 18575 67971 18581
rect 70854 18572 70860 18624
rect 70912 18612 70918 18624
rect 72513 18615 72571 18621
rect 72513 18612 72525 18615
rect 70912 18584 72525 18612
rect 70912 18572 70918 18584
rect 72513 18581 72525 18584
rect 72559 18581 72571 18615
rect 73890 18612 73896 18624
rect 73851 18584 73896 18612
rect 72513 18575 72571 18581
rect 73890 18572 73896 18584
rect 73948 18572 73954 18624
rect 74092 18612 74120 18779
rect 74184 18748 74212 18847
rect 74350 18844 74356 18896
rect 74408 18893 74414 18896
rect 74408 18887 74437 18893
rect 74425 18853 74437 18887
rect 74408 18847 74437 18853
rect 74408 18844 74414 18847
rect 74258 18776 74264 18828
rect 74316 18816 74322 18828
rect 74994 18816 75000 18828
rect 74316 18788 74361 18816
rect 74460 18788 75000 18816
rect 74316 18776 74322 18788
rect 74460 18748 74488 18788
rect 74994 18776 75000 18788
rect 75052 18776 75058 18828
rect 75181 18819 75239 18825
rect 75181 18785 75193 18819
rect 75227 18816 75239 18819
rect 144546 18816 144552 18828
rect 75227 18788 144552 18816
rect 75227 18785 75239 18788
rect 75181 18779 75239 18785
rect 74184 18720 74488 18748
rect 74537 18751 74595 18757
rect 74537 18717 74549 18751
rect 74583 18748 74595 18751
rect 75086 18748 75092 18760
rect 74583 18720 75092 18748
rect 74583 18717 74595 18720
rect 74537 18711 74595 18717
rect 75086 18708 75092 18720
rect 75144 18708 75150 18760
rect 74258 18640 74264 18692
rect 74316 18680 74322 18692
rect 75196 18680 75224 18779
rect 144546 18776 144552 18788
rect 144604 18776 144610 18828
rect 74316 18652 75224 18680
rect 74316 18640 74322 18652
rect 75822 18612 75828 18624
rect 74092 18584 75828 18612
rect 75822 18572 75828 18584
rect 75880 18572 75886 18624
rect 1104 18522 178848 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 34966 18522
rect 35018 18470 35030 18522
rect 35082 18470 35094 18522
rect 35146 18470 35158 18522
rect 35210 18470 65686 18522
rect 65738 18470 65750 18522
rect 65802 18470 65814 18522
rect 65866 18470 65878 18522
rect 65930 18470 96406 18522
rect 96458 18470 96470 18522
rect 96522 18470 96534 18522
rect 96586 18470 96598 18522
rect 96650 18470 127126 18522
rect 127178 18470 127190 18522
rect 127242 18470 127254 18522
rect 127306 18470 127318 18522
rect 127370 18470 157846 18522
rect 157898 18470 157910 18522
rect 157962 18470 157974 18522
rect 158026 18470 158038 18522
rect 158090 18470 178848 18522
rect 1104 18448 178848 18470
rect 31202 18368 31208 18420
rect 31260 18408 31266 18420
rect 31849 18411 31907 18417
rect 31849 18408 31861 18411
rect 31260 18380 31861 18408
rect 31260 18368 31266 18380
rect 31849 18377 31861 18380
rect 31895 18377 31907 18411
rect 31849 18371 31907 18377
rect 47026 18368 47032 18420
rect 47084 18408 47090 18420
rect 47578 18408 47584 18420
rect 47084 18380 47584 18408
rect 47084 18368 47090 18380
rect 47578 18368 47584 18380
rect 47636 18408 47642 18420
rect 60366 18408 60372 18420
rect 47636 18380 60372 18408
rect 47636 18368 47642 18380
rect 60366 18368 60372 18380
rect 60424 18368 60430 18420
rect 31481 18275 31539 18281
rect 31481 18241 31493 18275
rect 31527 18272 31539 18275
rect 33042 18272 33048 18284
rect 31527 18244 33048 18272
rect 31527 18241 31539 18244
rect 31481 18235 31539 18241
rect 33042 18232 33048 18244
rect 33100 18232 33106 18284
rect 47118 18272 47124 18284
rect 41386 18244 47124 18272
rect 41386 18216 41414 18244
rect 47118 18232 47124 18244
rect 47176 18232 47182 18284
rect 69658 18272 69664 18284
rect 51046 18244 69664 18272
rect 30650 18204 30656 18216
rect 30611 18176 30656 18204
rect 30650 18164 30656 18176
rect 30708 18164 30714 18216
rect 30837 18207 30895 18213
rect 30837 18173 30849 18207
rect 30883 18204 30895 18207
rect 31202 18204 31208 18216
rect 30883 18176 31208 18204
rect 30883 18173 30895 18176
rect 30837 18167 30895 18173
rect 31202 18164 31208 18176
rect 31260 18164 31266 18216
rect 31294 18164 31300 18216
rect 31352 18204 31358 18216
rect 31665 18207 31723 18213
rect 31665 18204 31677 18207
rect 31352 18176 31677 18204
rect 31352 18164 31358 18176
rect 31665 18173 31677 18176
rect 31711 18173 31723 18207
rect 31938 18204 31944 18216
rect 31899 18176 31944 18204
rect 31665 18167 31723 18173
rect 31938 18164 31944 18176
rect 31996 18204 32002 18216
rect 33134 18204 33140 18216
rect 31996 18176 33140 18204
rect 31996 18164 32002 18176
rect 33134 18164 33140 18176
rect 33192 18164 33198 18216
rect 37458 18164 37464 18216
rect 37516 18204 37522 18216
rect 39117 18207 39175 18213
rect 39117 18204 39129 18207
rect 37516 18176 39129 18204
rect 37516 18164 37522 18176
rect 39117 18173 39129 18176
rect 39163 18173 39175 18207
rect 39117 18167 39175 18173
rect 39209 18207 39267 18213
rect 39209 18173 39221 18207
rect 39255 18204 39267 18207
rect 40773 18207 40831 18213
rect 40773 18204 40785 18207
rect 39255 18176 40785 18204
rect 39255 18173 39267 18176
rect 39209 18167 39267 18173
rect 40773 18173 40785 18176
rect 40819 18173 40831 18207
rect 40773 18167 40831 18173
rect 41049 18207 41107 18213
rect 41049 18173 41061 18207
rect 41095 18204 41107 18207
rect 41386 18204 41420 18216
rect 41095 18176 41420 18204
rect 41095 18173 41107 18176
rect 41049 18167 41107 18173
rect 30745 18139 30803 18145
rect 30745 18105 30757 18139
rect 30791 18136 30803 18139
rect 31846 18136 31852 18148
rect 30791 18108 31852 18136
rect 30791 18105 30803 18108
rect 30745 18099 30803 18105
rect 31846 18096 31852 18108
rect 31904 18096 31910 18148
rect 40788 18068 40816 18167
rect 41414 18164 41420 18176
rect 41472 18164 41478 18216
rect 46109 18207 46167 18213
rect 46109 18173 46121 18207
rect 46155 18204 46167 18207
rect 47026 18204 47032 18216
rect 46155 18176 47032 18204
rect 46155 18173 46167 18176
rect 46109 18167 46167 18173
rect 47026 18164 47032 18176
rect 47084 18164 47090 18216
rect 48314 18164 48320 18216
rect 48372 18204 48378 18216
rect 49421 18207 49479 18213
rect 49421 18204 49433 18207
rect 48372 18176 49433 18204
rect 48372 18164 48378 18176
rect 49421 18173 49433 18176
rect 49467 18173 49479 18207
rect 49421 18167 49479 18173
rect 49510 18164 49516 18216
rect 49568 18204 49574 18216
rect 49605 18207 49663 18213
rect 49605 18204 49617 18207
rect 49568 18176 49617 18204
rect 49568 18164 49574 18176
rect 49605 18173 49617 18176
rect 49651 18204 49663 18207
rect 51046 18204 51074 18244
rect 69658 18232 69664 18244
rect 69716 18232 69722 18284
rect 49651 18176 51074 18204
rect 49651 18173 49663 18176
rect 49605 18167 49663 18173
rect 52454 18164 52460 18216
rect 52512 18204 52518 18216
rect 53098 18204 53104 18216
rect 52512 18176 53104 18204
rect 52512 18164 52518 18176
rect 53098 18164 53104 18176
rect 53156 18204 53162 18216
rect 54021 18207 54079 18213
rect 54021 18204 54033 18207
rect 53156 18176 54033 18204
rect 53156 18164 53162 18176
rect 54021 18173 54033 18176
rect 54067 18173 54079 18207
rect 54202 18204 54208 18216
rect 54163 18176 54208 18204
rect 54021 18167 54079 18173
rect 54202 18164 54208 18176
rect 54260 18164 54266 18216
rect 72142 18204 72148 18216
rect 72103 18176 72148 18204
rect 72142 18164 72148 18176
rect 72200 18164 72206 18216
rect 73522 18204 73528 18216
rect 73483 18176 73528 18204
rect 73522 18164 73528 18176
rect 73580 18164 73586 18216
rect 41138 18136 41144 18148
rect 41099 18108 41144 18136
rect 41138 18096 41144 18108
rect 41196 18096 41202 18148
rect 54386 18136 54392 18148
rect 54347 18108 54392 18136
rect 54386 18096 54392 18108
rect 54444 18096 54450 18148
rect 41322 18068 41328 18080
rect 40788 18040 41328 18068
rect 41322 18028 41328 18040
rect 41380 18028 41386 18080
rect 46201 18071 46259 18077
rect 46201 18037 46213 18071
rect 46247 18068 46259 18071
rect 46382 18068 46388 18080
rect 46247 18040 46388 18068
rect 46247 18037 46259 18040
rect 46201 18031 46259 18037
rect 46382 18028 46388 18040
rect 46440 18028 46446 18080
rect 49602 18068 49608 18080
rect 49563 18040 49608 18068
rect 49602 18028 49608 18040
rect 49660 18028 49666 18080
rect 70762 18028 70768 18080
rect 70820 18068 70826 18080
rect 72237 18071 72295 18077
rect 72237 18068 72249 18071
rect 70820 18040 72249 18068
rect 70820 18028 70826 18040
rect 72237 18037 72249 18040
rect 72283 18037 72295 18071
rect 73614 18068 73620 18080
rect 73575 18040 73620 18068
rect 72237 18031 72295 18037
rect 73614 18028 73620 18040
rect 73672 18028 73678 18080
rect 1104 17978 178848 18000
rect 1104 17926 19606 17978
rect 19658 17926 19670 17978
rect 19722 17926 19734 17978
rect 19786 17926 19798 17978
rect 19850 17926 50326 17978
rect 50378 17926 50390 17978
rect 50442 17926 50454 17978
rect 50506 17926 50518 17978
rect 50570 17926 81046 17978
rect 81098 17926 81110 17978
rect 81162 17926 81174 17978
rect 81226 17926 81238 17978
rect 81290 17926 111766 17978
rect 111818 17926 111830 17978
rect 111882 17926 111894 17978
rect 111946 17926 111958 17978
rect 112010 17926 142486 17978
rect 142538 17926 142550 17978
rect 142602 17926 142614 17978
rect 142666 17926 142678 17978
rect 142730 17926 173206 17978
rect 173258 17926 173270 17978
rect 173322 17926 173334 17978
rect 173386 17926 173398 17978
rect 173450 17926 178848 17978
rect 1104 17904 178848 17926
rect 51537 17867 51595 17873
rect 51537 17833 51549 17867
rect 51583 17864 51595 17867
rect 52454 17864 52460 17876
rect 51583 17836 52460 17864
rect 51583 17833 51595 17836
rect 51537 17827 51595 17833
rect 52454 17824 52460 17836
rect 52512 17824 52518 17876
rect 60369 17799 60427 17805
rect 60369 17796 60381 17799
rect 59464 17768 60381 17796
rect 31294 17688 31300 17740
rect 31352 17728 31358 17740
rect 31757 17731 31815 17737
rect 31757 17728 31769 17731
rect 31352 17700 31769 17728
rect 31352 17688 31358 17700
rect 31757 17697 31769 17700
rect 31803 17697 31815 17731
rect 37458 17728 37464 17740
rect 37419 17700 37464 17728
rect 31757 17691 31815 17697
rect 37458 17688 37464 17700
rect 37516 17688 37522 17740
rect 37734 17728 37740 17740
rect 37695 17700 37740 17728
rect 37734 17688 37740 17700
rect 37792 17728 37798 17740
rect 38746 17728 38752 17740
rect 37792 17700 38752 17728
rect 37792 17688 37798 17700
rect 38746 17688 38752 17700
rect 38804 17688 38810 17740
rect 49602 17688 49608 17740
rect 49660 17728 49666 17740
rect 59464 17737 59492 17768
rect 60369 17765 60381 17768
rect 60415 17796 60427 17799
rect 61102 17796 61108 17808
rect 60415 17768 61108 17796
rect 60415 17765 60427 17768
rect 60369 17759 60427 17765
rect 61102 17756 61108 17768
rect 61160 17756 61166 17808
rect 51445 17731 51503 17737
rect 51445 17728 51457 17731
rect 49660 17700 51457 17728
rect 49660 17688 49666 17700
rect 51445 17697 51457 17700
rect 51491 17697 51503 17731
rect 51445 17691 51503 17697
rect 59449 17731 59507 17737
rect 59449 17697 59461 17731
rect 59495 17697 59507 17731
rect 59449 17691 59507 17697
rect 59538 17688 59544 17740
rect 59596 17728 59602 17740
rect 59725 17731 59783 17737
rect 59725 17728 59737 17731
rect 59596 17700 59737 17728
rect 59596 17688 59602 17700
rect 59725 17697 59737 17700
rect 59771 17728 59783 17731
rect 60182 17728 60188 17740
rect 59771 17700 60188 17728
rect 59771 17697 59783 17700
rect 59725 17691 59783 17697
rect 60182 17688 60188 17700
rect 60240 17688 60246 17740
rect 35802 17620 35808 17672
rect 35860 17660 35866 17672
rect 37645 17663 37703 17669
rect 37645 17660 37657 17663
rect 35860 17632 37657 17660
rect 35860 17620 35866 17632
rect 37645 17629 37657 17632
rect 37691 17629 37703 17663
rect 37645 17623 37703 17629
rect 37277 17595 37335 17601
rect 37277 17561 37289 17595
rect 37323 17592 37335 17595
rect 38838 17592 38844 17604
rect 37323 17564 38844 17592
rect 37323 17561 37335 17564
rect 37277 17555 37335 17561
rect 38838 17552 38844 17564
rect 38896 17552 38902 17604
rect 58342 17552 58348 17604
rect 58400 17592 58406 17604
rect 59170 17592 59176 17604
rect 58400 17564 59176 17592
rect 58400 17552 58406 17564
rect 59170 17552 59176 17564
rect 59228 17592 59234 17604
rect 59633 17595 59691 17601
rect 59633 17592 59645 17595
rect 59228 17564 59645 17592
rect 59228 17552 59234 17564
rect 59633 17561 59645 17564
rect 59679 17561 59691 17595
rect 59633 17555 59691 17561
rect 31849 17527 31907 17533
rect 31849 17493 31861 17527
rect 31895 17524 31907 17527
rect 32398 17524 32404 17536
rect 31895 17496 32404 17524
rect 31895 17493 31907 17496
rect 31849 17487 31907 17493
rect 32398 17484 32404 17496
rect 32456 17484 32462 17536
rect 59265 17527 59323 17533
rect 59265 17493 59277 17527
rect 59311 17524 59323 17527
rect 59538 17524 59544 17536
rect 59311 17496 59544 17524
rect 59311 17493 59323 17496
rect 59265 17487 59323 17493
rect 59538 17484 59544 17496
rect 59596 17484 59602 17536
rect 60550 17524 60556 17536
rect 60511 17496 60556 17524
rect 60550 17484 60556 17496
rect 60608 17484 60614 17536
rect 1104 17434 178848 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 34966 17434
rect 35018 17382 35030 17434
rect 35082 17382 35094 17434
rect 35146 17382 35158 17434
rect 35210 17382 65686 17434
rect 65738 17382 65750 17434
rect 65802 17382 65814 17434
rect 65866 17382 65878 17434
rect 65930 17382 96406 17434
rect 96458 17382 96470 17434
rect 96522 17382 96534 17434
rect 96586 17382 96598 17434
rect 96650 17382 127126 17434
rect 127178 17382 127190 17434
rect 127242 17382 127254 17434
rect 127306 17382 127318 17434
rect 127370 17382 157846 17434
rect 157898 17382 157910 17434
rect 157962 17382 157974 17434
rect 158026 17382 158038 17434
rect 158090 17382 178848 17434
rect 1104 17360 178848 17382
rect 45649 17323 45707 17329
rect 45649 17289 45661 17323
rect 45695 17320 45707 17323
rect 46934 17320 46940 17332
rect 45695 17292 46940 17320
rect 45695 17289 45707 17292
rect 45649 17283 45707 17289
rect 46934 17280 46940 17292
rect 46992 17280 46998 17332
rect 48314 17280 48320 17332
rect 48372 17320 48378 17332
rect 49421 17323 49479 17329
rect 49421 17320 49433 17323
rect 48372 17292 49433 17320
rect 48372 17280 48378 17292
rect 49421 17289 49433 17292
rect 49467 17289 49479 17323
rect 49421 17283 49479 17289
rect 59430 17323 59488 17329
rect 59430 17289 59442 17323
rect 59476 17320 59488 17323
rect 60550 17320 60556 17332
rect 59476 17292 60556 17320
rect 59476 17289 59488 17292
rect 59430 17283 59488 17289
rect 60550 17280 60556 17292
rect 60608 17280 60614 17332
rect 65870 17323 65928 17329
rect 65870 17289 65882 17323
rect 65916 17320 65928 17323
rect 67269 17323 67327 17329
rect 67269 17320 67281 17323
rect 65916 17292 67281 17320
rect 65916 17289 65928 17292
rect 65870 17283 65928 17289
rect 67269 17289 67281 17292
rect 67315 17289 67327 17323
rect 67269 17283 67327 17289
rect 70029 17323 70087 17329
rect 70029 17289 70041 17323
rect 70075 17320 70087 17323
rect 70394 17320 70400 17332
rect 70075 17292 70400 17320
rect 70075 17289 70087 17292
rect 70029 17283 70087 17289
rect 70394 17280 70400 17292
rect 70452 17320 70458 17332
rect 70854 17320 70860 17332
rect 70452 17292 70860 17320
rect 70452 17280 70458 17292
rect 70854 17280 70860 17292
rect 70912 17280 70918 17332
rect 72326 17320 72332 17332
rect 72239 17292 72332 17320
rect 72326 17280 72332 17292
rect 72384 17320 72390 17332
rect 73062 17320 73068 17332
rect 72384 17292 73068 17320
rect 72384 17280 72390 17292
rect 73062 17280 73068 17292
rect 73120 17280 73126 17332
rect 43622 17212 43628 17264
rect 43680 17252 43686 17264
rect 43717 17255 43775 17261
rect 43717 17252 43729 17255
rect 43680 17224 43729 17252
rect 43680 17212 43686 17224
rect 43717 17221 43729 17224
rect 43763 17221 43775 17255
rect 43717 17215 43775 17221
rect 57238 17212 57244 17264
rect 57296 17252 57302 17264
rect 57701 17255 57759 17261
rect 57701 17252 57713 17255
rect 57296 17224 57713 17252
rect 57296 17212 57302 17224
rect 57701 17221 57713 17224
rect 57747 17252 57759 17255
rect 59541 17255 59599 17261
rect 59541 17252 59553 17255
rect 57747 17224 59553 17252
rect 57747 17221 57759 17224
rect 57701 17215 57759 17221
rect 59541 17221 59553 17224
rect 59587 17221 59599 17255
rect 59541 17215 59599 17221
rect 63586 17212 63592 17264
rect 63644 17252 63650 17264
rect 64601 17255 64659 17261
rect 64601 17252 64613 17255
rect 63644 17224 64613 17252
rect 63644 17212 63650 17224
rect 64601 17221 64613 17224
rect 64647 17252 64659 17255
rect 65978 17252 65984 17264
rect 64647 17224 65984 17252
rect 64647 17221 64659 17224
rect 64601 17215 64659 17221
rect 65978 17212 65984 17224
rect 66036 17212 66042 17264
rect 35802 17184 35808 17196
rect 34992 17156 35808 17184
rect 34992 17125 35020 17156
rect 35802 17144 35808 17156
rect 35860 17144 35866 17196
rect 49602 17184 49608 17196
rect 49252 17156 49608 17184
rect 34977 17119 35035 17125
rect 34977 17085 34989 17119
rect 35023 17085 35035 17119
rect 35250 17116 35256 17128
rect 35211 17088 35256 17116
rect 34977 17079 35035 17085
rect 35250 17076 35256 17088
rect 35308 17076 35314 17128
rect 35437 17119 35495 17125
rect 35437 17085 35449 17119
rect 35483 17116 35495 17119
rect 35894 17116 35900 17128
rect 35483 17088 35900 17116
rect 35483 17085 35495 17088
rect 35437 17079 35495 17085
rect 35894 17076 35900 17088
rect 35952 17076 35958 17128
rect 43346 17076 43352 17128
rect 43404 17116 43410 17128
rect 43625 17119 43683 17125
rect 43625 17116 43637 17119
rect 43404 17088 43637 17116
rect 43404 17076 43410 17088
rect 43625 17085 43637 17088
rect 43671 17085 43683 17119
rect 43625 17079 43683 17085
rect 43901 17119 43959 17125
rect 43901 17085 43913 17119
rect 43947 17116 43959 17119
rect 44082 17116 44088 17128
rect 43947 17088 44088 17116
rect 43947 17085 43959 17088
rect 43901 17079 43959 17085
rect 44082 17076 44088 17088
rect 44140 17076 44146 17128
rect 44361 17119 44419 17125
rect 44361 17085 44373 17119
rect 44407 17116 44419 17119
rect 45557 17119 45615 17125
rect 45557 17116 45569 17119
rect 44407 17088 45569 17116
rect 44407 17085 44419 17088
rect 44361 17079 44419 17085
rect 45557 17085 45569 17088
rect 45603 17116 45615 17119
rect 46198 17116 46204 17128
rect 45603 17088 46204 17116
rect 45603 17085 45615 17088
rect 45557 17079 45615 17085
rect 46198 17076 46204 17088
rect 46256 17076 46262 17128
rect 49252 17125 49280 17156
rect 49602 17144 49608 17156
rect 49660 17144 49666 17196
rect 59354 17184 59360 17196
rect 57900 17156 59360 17184
rect 49237 17119 49295 17125
rect 49237 17085 49249 17119
rect 49283 17085 49295 17119
rect 49510 17116 49516 17128
rect 49471 17088 49516 17116
rect 49237 17079 49295 17085
rect 49510 17076 49516 17088
rect 49568 17076 49574 17128
rect 57900 17125 57928 17156
rect 59354 17144 59360 17156
rect 59412 17184 59418 17196
rect 59633 17187 59691 17193
rect 59633 17184 59645 17187
rect 59412 17156 59645 17184
rect 59412 17144 59418 17156
rect 59633 17153 59645 17156
rect 59679 17153 59691 17187
rect 66073 17187 66131 17193
rect 66073 17184 66085 17187
rect 59633 17147 59691 17153
rect 64800 17156 66085 17184
rect 57609 17119 57667 17125
rect 57609 17085 57621 17119
rect 57655 17085 57667 17119
rect 57609 17079 57667 17085
rect 57885 17119 57943 17125
rect 57885 17085 57897 17119
rect 57931 17085 57943 17119
rect 58342 17116 58348 17128
rect 58303 17088 58348 17116
rect 57885 17079 57943 17085
rect 56686 17008 56692 17060
rect 56744 17048 56750 17060
rect 56962 17048 56968 17060
rect 56744 17020 56968 17048
rect 56744 17008 56750 17020
rect 56962 17008 56968 17020
rect 57020 17048 57026 17060
rect 57624 17048 57652 17079
rect 58342 17076 58348 17088
rect 58400 17076 58406 17128
rect 63494 17076 63500 17128
rect 63552 17116 63558 17128
rect 64800 17125 64828 17156
rect 66073 17153 66085 17156
rect 66119 17184 66131 17187
rect 66162 17184 66168 17196
rect 66119 17156 66168 17184
rect 66119 17153 66131 17156
rect 66073 17147 66131 17153
rect 66162 17144 66168 17156
rect 66220 17144 66226 17196
rect 75086 17184 75092 17196
rect 73080 17156 75092 17184
rect 64509 17119 64567 17125
rect 64509 17116 64521 17119
rect 63552 17088 64521 17116
rect 63552 17076 63558 17088
rect 64509 17085 64521 17088
rect 64555 17085 64567 17119
rect 64509 17079 64567 17085
rect 64785 17119 64843 17125
rect 64785 17085 64797 17119
rect 64831 17085 64843 17119
rect 65705 17119 65763 17125
rect 65705 17116 65717 17119
rect 64785 17079 64843 17085
rect 64892 17088 65717 17116
rect 59265 17051 59323 17057
rect 59265 17048 59277 17051
rect 57020 17020 59277 17048
rect 57020 17008 57026 17020
rect 59265 17017 59277 17020
rect 59311 17017 59323 17051
rect 64524 17048 64552 17079
rect 64892 17048 64920 17088
rect 65705 17085 65717 17088
rect 65751 17085 65763 17119
rect 66898 17116 66904 17128
rect 66859 17088 66904 17116
rect 65705 17079 65763 17085
rect 66898 17076 66904 17088
rect 66956 17076 66962 17128
rect 67082 17116 67088 17128
rect 67043 17088 67088 17116
rect 67082 17076 67088 17088
rect 67140 17076 67146 17128
rect 69842 17116 69848 17128
rect 69803 17088 69848 17116
rect 69842 17076 69848 17088
rect 69900 17076 69906 17128
rect 70029 17119 70087 17125
rect 70029 17085 70041 17119
rect 70075 17116 70087 17119
rect 70762 17116 70768 17128
rect 70075 17088 70768 17116
rect 70075 17085 70087 17088
rect 70029 17079 70087 17085
rect 70762 17076 70768 17088
rect 70820 17076 70826 17128
rect 71130 17116 71136 17128
rect 71091 17088 71136 17116
rect 71130 17076 71136 17088
rect 71188 17076 71194 17128
rect 71314 17116 71320 17128
rect 71275 17088 71320 17116
rect 71314 17076 71320 17088
rect 71372 17076 71378 17128
rect 71682 17076 71688 17128
rect 71740 17116 71746 17128
rect 73080 17125 73108 17156
rect 75086 17144 75092 17156
rect 75144 17144 75150 17196
rect 72237 17119 72295 17125
rect 72237 17116 72249 17119
rect 71740 17088 72249 17116
rect 71740 17076 71746 17088
rect 72237 17085 72249 17088
rect 72283 17085 72295 17119
rect 72237 17079 72295 17085
rect 73065 17119 73123 17125
rect 73065 17085 73077 17119
rect 73111 17085 73123 17119
rect 73246 17116 73252 17128
rect 73207 17088 73252 17116
rect 73065 17079 73123 17085
rect 73246 17076 73252 17088
rect 73304 17076 73310 17128
rect 73341 17119 73399 17125
rect 73341 17085 73353 17119
rect 73387 17116 73399 17119
rect 74258 17116 74264 17128
rect 73387 17088 74264 17116
rect 73387 17085 73399 17088
rect 73341 17079 73399 17085
rect 64524 17020 64920 17048
rect 65245 17051 65303 17057
rect 59265 17011 59323 17017
rect 65245 17017 65257 17051
rect 65291 17017 65303 17051
rect 65245 17011 65303 17017
rect 34793 16983 34851 16989
rect 34793 16949 34805 16983
rect 34839 16980 34851 16983
rect 36354 16980 36360 16992
rect 34839 16952 36360 16980
rect 34839 16949 34851 16952
rect 34793 16943 34851 16949
rect 36354 16940 36360 16952
rect 36412 16940 36418 16992
rect 49050 16980 49056 16992
rect 49011 16952 49056 16980
rect 49050 16940 49056 16952
rect 49108 16940 49114 16992
rect 59722 16940 59728 16992
rect 59780 16980 59786 16992
rect 59909 16983 59967 16989
rect 59909 16980 59921 16983
rect 59780 16952 59921 16980
rect 59780 16940 59786 16952
rect 59909 16949 59921 16952
rect 59955 16949 59967 16983
rect 65260 16980 65288 17011
rect 69934 17008 69940 17060
rect 69992 17048 69998 17060
rect 73356 17048 73384 17079
rect 74258 17076 74264 17088
rect 74316 17076 74322 17128
rect 69992 17020 73384 17048
rect 69992 17008 69998 17020
rect 66162 16980 66168 16992
rect 65260 16952 66168 16980
rect 59909 16943 59967 16949
rect 66162 16940 66168 16952
rect 66220 16940 66226 16992
rect 66346 16980 66352 16992
rect 66307 16952 66352 16980
rect 66346 16940 66352 16952
rect 66404 16940 66410 16992
rect 70210 16980 70216 16992
rect 70171 16952 70216 16980
rect 70210 16940 70216 16952
rect 70268 16940 70274 16992
rect 71498 16980 71504 16992
rect 71459 16952 71504 16980
rect 71498 16940 71504 16952
rect 71556 16940 71562 16992
rect 72510 16940 72516 16992
rect 72568 16980 72574 16992
rect 72881 16983 72939 16989
rect 72881 16980 72893 16983
rect 72568 16952 72893 16980
rect 72568 16940 72574 16952
rect 72881 16949 72893 16952
rect 72927 16949 72939 16983
rect 72881 16943 72939 16949
rect 1104 16890 178848 16912
rect 1104 16838 19606 16890
rect 19658 16838 19670 16890
rect 19722 16838 19734 16890
rect 19786 16838 19798 16890
rect 19850 16838 50326 16890
rect 50378 16838 50390 16890
rect 50442 16838 50454 16890
rect 50506 16838 50518 16890
rect 50570 16838 81046 16890
rect 81098 16838 81110 16890
rect 81162 16838 81174 16890
rect 81226 16838 81238 16890
rect 81290 16838 111766 16890
rect 111818 16838 111830 16890
rect 111882 16838 111894 16890
rect 111946 16838 111958 16890
rect 112010 16838 142486 16890
rect 142538 16838 142550 16890
rect 142602 16838 142614 16890
rect 142666 16838 142678 16890
rect 142730 16838 173206 16890
rect 173258 16838 173270 16890
rect 173322 16838 173334 16890
rect 173386 16838 173398 16890
rect 173450 16838 178848 16890
rect 1104 16816 178848 16838
rect 32122 16736 32128 16788
rect 32180 16736 32186 16788
rect 32223 16779 32281 16785
rect 32223 16745 32235 16779
rect 32269 16776 32281 16779
rect 33686 16776 33692 16788
rect 32269 16748 33692 16776
rect 32269 16745 32281 16748
rect 32223 16739 32281 16745
rect 33686 16736 33692 16748
rect 33744 16736 33750 16788
rect 42886 16776 42892 16788
rect 42847 16748 42892 16776
rect 42886 16736 42892 16748
rect 42944 16776 42950 16788
rect 43622 16776 43628 16788
rect 42944 16748 43628 16776
rect 42944 16736 42950 16748
rect 43622 16736 43628 16748
rect 43680 16736 43686 16788
rect 60090 16776 60096 16788
rect 58728 16748 60096 16776
rect 32140 16708 32168 16736
rect 32309 16711 32367 16717
rect 32309 16708 32321 16711
rect 32140 16680 32321 16708
rect 32309 16677 32321 16680
rect 32355 16677 32367 16711
rect 43806 16708 43812 16720
rect 32309 16671 32367 16677
rect 42536 16680 43812 16708
rect 32125 16643 32183 16649
rect 32125 16609 32137 16643
rect 32171 16640 32183 16643
rect 32214 16640 32220 16652
rect 32171 16612 32220 16640
rect 32171 16609 32183 16612
rect 32125 16603 32183 16609
rect 32214 16600 32220 16612
rect 32272 16600 32278 16652
rect 32398 16640 32404 16652
rect 32359 16612 32404 16640
rect 32398 16600 32404 16612
rect 32456 16600 32462 16652
rect 40954 16640 40960 16652
rect 40915 16612 40960 16640
rect 40954 16600 40960 16612
rect 41012 16600 41018 16652
rect 41138 16640 41144 16652
rect 41099 16612 41144 16640
rect 41138 16600 41144 16612
rect 41196 16640 41202 16652
rect 42536 16649 42564 16680
rect 43806 16668 43812 16680
rect 43864 16668 43870 16720
rect 48314 16708 48320 16720
rect 47412 16680 48320 16708
rect 42521 16643 42579 16649
rect 41196 16612 42472 16640
rect 41196 16600 41202 16612
rect 41322 16572 41328 16584
rect 41283 16544 41328 16572
rect 41322 16532 41328 16544
rect 41380 16532 41386 16584
rect 41414 16532 41420 16584
rect 41472 16572 41478 16584
rect 42444 16572 42472 16612
rect 42521 16609 42533 16643
rect 42567 16609 42579 16643
rect 42981 16643 43039 16649
rect 42981 16640 42993 16643
rect 42521 16603 42579 16609
rect 42628 16612 42993 16640
rect 42628 16572 42656 16612
rect 42981 16609 42993 16612
rect 43027 16640 43039 16643
rect 43346 16640 43352 16652
rect 43027 16612 43352 16640
rect 43027 16609 43039 16612
rect 42981 16603 43039 16609
rect 43346 16600 43352 16612
rect 43404 16640 43410 16652
rect 43441 16643 43499 16649
rect 43441 16640 43453 16643
rect 43404 16612 43453 16640
rect 43404 16600 43410 16612
rect 43441 16609 43453 16612
rect 43487 16609 43499 16643
rect 43622 16640 43628 16652
rect 43583 16612 43628 16640
rect 43441 16603 43499 16609
rect 43622 16600 43628 16612
rect 43680 16600 43686 16652
rect 46198 16640 46204 16652
rect 46159 16612 46204 16640
rect 46198 16600 46204 16612
rect 46256 16600 46262 16652
rect 46382 16640 46388 16652
rect 46343 16612 46388 16640
rect 46382 16600 46388 16612
rect 46440 16600 46446 16652
rect 47210 16640 47216 16652
rect 47171 16612 47216 16640
rect 47210 16600 47216 16612
rect 47268 16600 47274 16652
rect 47412 16649 47440 16680
rect 48314 16668 48320 16680
rect 48372 16668 48378 16720
rect 54386 16708 54392 16720
rect 52932 16680 54392 16708
rect 47397 16643 47455 16649
rect 47397 16609 47409 16643
rect 47443 16609 47455 16643
rect 47397 16603 47455 16609
rect 47673 16643 47731 16649
rect 47673 16609 47685 16643
rect 47719 16609 47731 16643
rect 47854 16640 47860 16652
rect 47815 16612 47860 16640
rect 47673 16603 47731 16609
rect 41472 16544 41517 16572
rect 42444 16544 42656 16572
rect 46293 16575 46351 16581
rect 41472 16532 41478 16544
rect 46293 16541 46305 16575
rect 46339 16572 46351 16575
rect 46934 16572 46940 16584
rect 46339 16544 46940 16572
rect 46339 16541 46351 16544
rect 46293 16535 46351 16541
rect 46934 16532 46940 16544
rect 46992 16572 46998 16584
rect 47688 16572 47716 16603
rect 47854 16600 47860 16612
rect 47912 16600 47918 16652
rect 52730 16640 52736 16652
rect 52691 16612 52736 16640
rect 52730 16600 52736 16612
rect 52788 16600 52794 16652
rect 52932 16649 52960 16680
rect 54386 16668 54392 16680
rect 54444 16708 54450 16720
rect 54444 16680 56732 16708
rect 54444 16668 54450 16680
rect 56704 16652 56732 16680
rect 58728 16652 58756 16748
rect 60090 16736 60096 16748
rect 60148 16736 60154 16788
rect 59633 16711 59691 16717
rect 59633 16708 59645 16711
rect 58820 16680 59645 16708
rect 52917 16643 52975 16649
rect 52917 16609 52929 16643
rect 52963 16609 52975 16643
rect 53190 16640 53196 16652
rect 53103 16612 53196 16640
rect 52917 16603 52975 16609
rect 53190 16600 53196 16612
rect 53248 16640 53254 16652
rect 54202 16640 54208 16652
rect 53248 16612 54208 16640
rect 53248 16600 53254 16612
rect 54202 16600 54208 16612
rect 54260 16600 54266 16652
rect 56686 16640 56692 16652
rect 56647 16612 56692 16640
rect 56686 16600 56692 16612
rect 56744 16600 56750 16652
rect 56870 16640 56876 16652
rect 56783 16612 56876 16640
rect 56870 16600 56876 16612
rect 56928 16640 56934 16652
rect 57238 16640 57244 16652
rect 56928 16612 57244 16640
rect 56928 16600 56934 16612
rect 57238 16600 57244 16612
rect 57296 16600 57302 16652
rect 58250 16600 58256 16652
rect 58308 16640 58314 16652
rect 58529 16643 58587 16649
rect 58529 16640 58541 16643
rect 58308 16612 58541 16640
rect 58308 16600 58314 16612
rect 58529 16609 58541 16612
rect 58575 16609 58587 16643
rect 58710 16640 58716 16652
rect 58623 16612 58716 16640
rect 58529 16603 58587 16609
rect 58710 16600 58716 16612
rect 58768 16600 58774 16652
rect 58820 16649 58848 16680
rect 59633 16677 59645 16680
rect 59679 16677 59691 16711
rect 59633 16671 59691 16677
rect 66346 16668 66352 16720
rect 66404 16708 66410 16720
rect 69842 16708 69848 16720
rect 66404 16680 69848 16708
rect 66404 16668 66410 16680
rect 58805 16643 58863 16649
rect 58805 16609 58817 16643
rect 58851 16609 58863 16643
rect 58805 16603 58863 16609
rect 59081 16643 59139 16649
rect 59081 16609 59093 16643
rect 59127 16640 59139 16643
rect 59446 16640 59452 16652
rect 59127 16612 59452 16640
rect 59127 16609 59139 16612
rect 59081 16603 59139 16609
rect 59446 16600 59452 16612
rect 59504 16600 59510 16652
rect 59541 16643 59599 16649
rect 59541 16609 59553 16643
rect 59587 16609 59599 16643
rect 59541 16603 59599 16609
rect 53098 16572 53104 16584
rect 46992 16544 47716 16572
rect 53059 16544 53104 16572
rect 46992 16532 46998 16544
rect 53098 16532 53104 16544
rect 53156 16532 53162 16584
rect 59170 16532 59176 16584
rect 59228 16572 59234 16584
rect 59556 16572 59584 16603
rect 65518 16600 65524 16652
rect 65576 16640 65582 16652
rect 65797 16643 65855 16649
rect 65797 16640 65809 16643
rect 65576 16612 65809 16640
rect 65576 16600 65582 16612
rect 65797 16609 65809 16612
rect 65843 16609 65855 16643
rect 65797 16603 65855 16609
rect 65981 16643 66039 16649
rect 65981 16609 65993 16643
rect 66027 16640 66039 16643
rect 67082 16640 67088 16652
rect 66027 16612 67088 16640
rect 66027 16609 66039 16612
rect 65981 16603 66039 16609
rect 67082 16600 67088 16612
rect 67140 16600 67146 16652
rect 68940 16649 68968 16680
rect 69842 16668 69848 16680
rect 69900 16708 69906 16720
rect 70397 16711 70455 16717
rect 70397 16708 70409 16711
rect 69900 16680 70409 16708
rect 69900 16668 69906 16680
rect 70397 16677 70409 16680
rect 70443 16677 70455 16711
rect 73246 16708 73252 16720
rect 70397 16671 70455 16677
rect 72620 16680 73252 16708
rect 68925 16643 68983 16649
rect 68925 16609 68937 16643
rect 68971 16609 68983 16643
rect 68925 16603 68983 16609
rect 69109 16643 69167 16649
rect 69109 16609 69121 16643
rect 69155 16640 69167 16643
rect 70544 16643 70602 16649
rect 69155 16612 70348 16640
rect 69155 16609 69167 16612
rect 69109 16603 69167 16609
rect 66254 16572 66260 16584
rect 59228 16544 59584 16572
rect 66167 16544 66260 16572
rect 59228 16532 59234 16544
rect 66254 16532 66260 16544
rect 66312 16572 66318 16584
rect 66898 16572 66904 16584
rect 66312 16544 66904 16572
rect 66312 16532 66318 16544
rect 66898 16532 66904 16544
rect 66956 16532 66962 16584
rect 70320 16572 70348 16612
rect 70544 16609 70556 16643
rect 70590 16640 70602 16643
rect 71498 16640 71504 16652
rect 70590 16612 71504 16640
rect 70590 16609 70602 16612
rect 70544 16603 70602 16609
rect 71498 16600 71504 16612
rect 71556 16600 71562 16652
rect 72418 16640 72424 16652
rect 72379 16612 72424 16640
rect 72418 16600 72424 16612
rect 72476 16600 72482 16652
rect 72620 16649 72648 16680
rect 73246 16668 73252 16680
rect 73304 16668 73310 16720
rect 72605 16643 72663 16649
rect 72605 16609 72617 16643
rect 72651 16609 72663 16643
rect 72878 16640 72884 16652
rect 72839 16612 72884 16640
rect 72605 16603 72663 16609
rect 72878 16600 72884 16612
rect 72936 16600 72942 16652
rect 73062 16640 73068 16652
rect 72975 16612 73068 16640
rect 73062 16600 73068 16612
rect 73120 16640 73126 16652
rect 75270 16640 75276 16652
rect 73120 16612 75276 16640
rect 73120 16600 73126 16612
rect 75270 16600 75276 16612
rect 75328 16600 75334 16652
rect 70394 16572 70400 16584
rect 70320 16544 70400 16572
rect 70394 16532 70400 16544
rect 70452 16532 70458 16584
rect 70762 16572 70768 16584
rect 70723 16544 70768 16572
rect 70762 16532 70768 16544
rect 70820 16532 70826 16584
rect 71133 16575 71191 16581
rect 71133 16541 71145 16575
rect 71179 16572 71191 16575
rect 71682 16572 71688 16584
rect 71179 16544 71688 16572
rect 71179 16541 71191 16544
rect 71133 16535 71191 16541
rect 71682 16532 71688 16544
rect 71740 16532 71746 16584
rect 70412 16504 70440 16532
rect 70673 16507 70731 16513
rect 70673 16504 70685 16507
rect 70412 16476 70685 16504
rect 70673 16473 70685 16476
rect 70719 16473 70731 16507
rect 70673 16467 70731 16473
rect 42705 16439 42763 16445
rect 42705 16405 42717 16439
rect 42751 16436 42763 16439
rect 42794 16436 42800 16448
rect 42751 16408 42800 16436
rect 42751 16405 42763 16408
rect 42705 16399 42763 16405
rect 42794 16396 42800 16408
rect 42852 16396 42858 16448
rect 56686 16436 56692 16448
rect 56647 16408 56692 16436
rect 56686 16396 56692 16408
rect 56744 16396 56750 16448
rect 58986 16436 58992 16448
rect 58947 16408 58992 16436
rect 58986 16396 58992 16408
rect 59044 16396 59050 16448
rect 66162 16436 66168 16448
rect 66123 16408 66168 16436
rect 66162 16396 66168 16408
rect 66220 16396 66226 16448
rect 68922 16436 68928 16448
rect 68883 16408 68928 16436
rect 68922 16396 68928 16408
rect 68980 16396 68986 16448
rect 1104 16346 178848 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 34966 16346
rect 35018 16294 35030 16346
rect 35082 16294 35094 16346
rect 35146 16294 35158 16346
rect 35210 16294 65686 16346
rect 65738 16294 65750 16346
rect 65802 16294 65814 16346
rect 65866 16294 65878 16346
rect 65930 16294 96406 16346
rect 96458 16294 96470 16346
rect 96522 16294 96534 16346
rect 96586 16294 96598 16346
rect 96650 16294 127126 16346
rect 127178 16294 127190 16346
rect 127242 16294 127254 16346
rect 127306 16294 127318 16346
rect 127370 16294 157846 16346
rect 157898 16294 157910 16346
rect 157962 16294 157974 16346
rect 158026 16294 158038 16346
rect 158090 16294 178848 16346
rect 1104 16272 178848 16294
rect 32033 16235 32091 16241
rect 32033 16201 32045 16235
rect 32079 16232 32091 16235
rect 32398 16232 32404 16244
rect 32079 16204 32404 16232
rect 32079 16201 32091 16204
rect 32033 16195 32091 16201
rect 32398 16192 32404 16204
rect 32456 16192 32462 16244
rect 33229 16235 33287 16241
rect 33229 16201 33241 16235
rect 33275 16201 33287 16235
rect 33229 16195 33287 16201
rect 33413 16235 33471 16241
rect 33413 16201 33425 16235
rect 33459 16232 33471 16235
rect 34514 16232 34520 16244
rect 33459 16204 34520 16232
rect 33459 16201 33471 16204
rect 33413 16195 33471 16201
rect 31481 16167 31539 16173
rect 31481 16133 31493 16167
rect 31527 16164 31539 16167
rect 31938 16164 31944 16176
rect 31527 16136 31944 16164
rect 31527 16133 31539 16136
rect 31481 16127 31539 16133
rect 31938 16124 31944 16136
rect 31996 16124 32002 16176
rect 33244 16164 33272 16195
rect 34514 16192 34520 16204
rect 34572 16232 34578 16244
rect 35250 16232 35256 16244
rect 34572 16204 35256 16232
rect 34572 16192 34578 16204
rect 35250 16192 35256 16204
rect 35308 16192 35314 16244
rect 69014 16192 69020 16244
rect 69072 16232 69078 16244
rect 71133 16235 71191 16241
rect 71133 16232 71145 16235
rect 69072 16204 71145 16232
rect 69072 16192 69078 16204
rect 71133 16201 71145 16204
rect 71179 16201 71191 16235
rect 71866 16232 71872 16244
rect 71779 16204 71872 16232
rect 71133 16195 71191 16201
rect 71866 16192 71872 16204
rect 71924 16232 71930 16244
rect 72878 16232 72884 16244
rect 71924 16204 72884 16232
rect 71924 16192 71930 16204
rect 72878 16192 72884 16204
rect 72936 16192 72942 16244
rect 32140 16136 33272 16164
rect 44085 16167 44143 16173
rect 32140 16096 32168 16136
rect 44085 16133 44097 16167
rect 44131 16164 44143 16167
rect 44726 16164 44732 16176
rect 44131 16136 44732 16164
rect 44131 16133 44143 16136
rect 44085 16127 44143 16133
rect 44726 16124 44732 16136
rect 44784 16124 44790 16176
rect 45830 16164 45836 16176
rect 45791 16136 45836 16164
rect 45830 16124 45836 16136
rect 45888 16124 45894 16176
rect 67818 16164 67824 16176
rect 65536 16136 67824 16164
rect 46934 16096 46940 16108
rect 31680 16068 32168 16096
rect 31680 16037 31708 16068
rect 32140 16040 32168 16068
rect 45848 16068 46940 16096
rect 31662 16031 31720 16037
rect 31662 15997 31674 16031
rect 31708 15997 31720 16031
rect 31662 15991 31720 15997
rect 32122 15988 32128 16040
rect 32180 16028 32186 16040
rect 32180 16000 32225 16028
rect 32180 15988 32186 16000
rect 43806 15988 43812 16040
rect 43864 16028 43870 16040
rect 45848 16037 45876 16068
rect 46934 16056 46940 16068
rect 46992 16056 46998 16108
rect 56686 16056 56692 16108
rect 56744 16096 56750 16108
rect 57425 16099 57483 16105
rect 57425 16096 57437 16099
rect 56744 16068 57437 16096
rect 56744 16056 56750 16068
rect 57425 16065 57437 16068
rect 57471 16065 57483 16099
rect 65536 16096 65564 16136
rect 67818 16124 67824 16136
rect 67876 16124 67882 16176
rect 65702 16096 65708 16108
rect 57425 16059 57483 16065
rect 65444 16068 65564 16096
rect 65663 16068 65708 16096
rect 44361 16031 44419 16037
rect 44361 16028 44373 16031
rect 43864 16000 44373 16028
rect 43864 15988 43870 16000
rect 44361 15997 44373 16000
rect 44407 15997 44419 16031
rect 44361 15991 44419 15997
rect 45833 16031 45891 16037
rect 45833 15997 45845 16031
rect 45879 15997 45891 16031
rect 45833 15991 45891 15997
rect 46109 16031 46167 16037
rect 46109 15997 46121 16031
rect 46155 16028 46167 16031
rect 46198 16028 46204 16040
rect 46155 16000 46204 16028
rect 46155 15997 46167 16000
rect 46109 15991 46167 15997
rect 46198 15988 46204 16000
rect 46256 15988 46262 16040
rect 57241 16031 57299 16037
rect 57241 15997 57253 16031
rect 57287 15997 57299 16031
rect 57241 15991 57299 15997
rect 57517 16031 57575 16037
rect 57517 15997 57529 16031
rect 57563 16028 57575 16031
rect 58066 16028 58072 16040
rect 57563 16000 58072 16028
rect 57563 15997 57575 16000
rect 57517 15991 57575 15997
rect 32214 15920 32220 15972
rect 32272 15960 32278 15972
rect 33045 15963 33103 15969
rect 33045 15960 33057 15963
rect 32272 15932 33057 15960
rect 32272 15920 32278 15932
rect 33045 15929 33057 15932
rect 33091 15960 33103 15963
rect 36078 15960 36084 15972
rect 33091 15932 36084 15960
rect 33091 15929 33103 15932
rect 33045 15923 33103 15929
rect 36078 15920 36084 15932
rect 36136 15920 36142 15972
rect 44085 15963 44143 15969
rect 44085 15929 44097 15963
rect 44131 15929 44143 15963
rect 44085 15923 44143 15929
rect 31665 15895 31723 15901
rect 31665 15861 31677 15895
rect 31711 15892 31723 15895
rect 32398 15892 32404 15904
rect 31711 15864 32404 15892
rect 31711 15861 31723 15864
rect 31665 15855 31723 15861
rect 32398 15852 32404 15864
rect 32456 15892 32462 15904
rect 33250 15895 33308 15901
rect 33250 15892 33262 15895
rect 32456 15864 33262 15892
rect 32456 15852 32462 15864
rect 33250 15861 33262 15864
rect 33296 15861 33308 15895
rect 44100 15892 44128 15923
rect 44174 15920 44180 15972
rect 44232 15960 44238 15972
rect 44269 15963 44327 15969
rect 44269 15960 44281 15963
rect 44232 15932 44281 15960
rect 44232 15920 44238 15932
rect 44269 15929 44281 15932
rect 44315 15929 44327 15963
rect 44269 15923 44327 15929
rect 46017 15963 46075 15969
rect 46017 15929 46029 15963
rect 46063 15960 46075 15963
rect 46382 15960 46388 15972
rect 46063 15932 46388 15960
rect 46063 15929 46075 15932
rect 46017 15923 46075 15929
rect 46382 15920 46388 15932
rect 46440 15920 46446 15972
rect 57256 15960 57284 15991
rect 58066 15988 58072 16000
rect 58124 15988 58130 16040
rect 63405 16031 63463 16037
rect 63405 15997 63417 16031
rect 63451 16028 63463 16031
rect 63494 16028 63500 16040
rect 63451 16000 63500 16028
rect 63451 15997 63463 16000
rect 63405 15991 63463 15997
rect 63494 15988 63500 16000
rect 63552 15988 63558 16040
rect 63586 15988 63592 16040
rect 63644 16028 63650 16040
rect 63644 16000 63689 16028
rect 63644 15988 63650 16000
rect 65334 15988 65340 16040
rect 65392 16028 65398 16040
rect 65444 16037 65472 16068
rect 65702 16056 65708 16068
rect 65760 16096 65766 16108
rect 66162 16096 66168 16108
rect 65760 16068 66168 16096
rect 65760 16056 65766 16068
rect 66162 16056 66168 16068
rect 66220 16096 66226 16108
rect 71130 16096 71136 16108
rect 66220 16068 66300 16096
rect 66220 16056 66226 16068
rect 65429 16031 65487 16037
rect 65429 16028 65441 16031
rect 65392 16000 65441 16028
rect 65392 15988 65398 16000
rect 65429 15997 65441 16000
rect 65475 15997 65487 16031
rect 65429 15991 65487 15997
rect 65521 16031 65579 16037
rect 65521 15997 65533 16031
rect 65567 15997 65579 16031
rect 65521 15991 65579 15997
rect 65797 16031 65855 16037
rect 65797 15997 65809 16031
rect 65843 16028 65855 16031
rect 66070 16028 66076 16040
rect 65843 16000 66076 16028
rect 65843 15997 65855 16000
rect 65797 15991 65855 15997
rect 58986 15960 58992 15972
rect 57256 15932 58992 15960
rect 58986 15920 58992 15932
rect 59044 15920 59050 15972
rect 65536 15960 65564 15991
rect 66070 15988 66076 16000
rect 66128 15988 66134 16040
rect 66272 16037 66300 16068
rect 70504 16068 71136 16096
rect 70504 16040 70532 16068
rect 71130 16056 71136 16068
rect 71188 16056 71194 16108
rect 66257 16031 66315 16037
rect 66257 15997 66269 16031
rect 66303 15997 66315 16031
rect 66257 15991 66315 15997
rect 70210 15988 70216 16040
rect 70268 16028 70274 16040
rect 70305 16031 70363 16037
rect 70305 16028 70317 16031
rect 70268 16000 70317 16028
rect 70268 15988 70274 16000
rect 70305 15997 70317 16000
rect 70351 15997 70363 16031
rect 70486 16028 70492 16040
rect 70399 16000 70492 16028
rect 70305 15991 70363 15997
rect 70486 15988 70492 16000
rect 70544 15988 70550 16040
rect 70673 16031 70731 16037
rect 70673 15997 70685 16031
rect 70719 16028 70731 16031
rect 71409 16031 71467 16037
rect 71409 16028 71421 16031
rect 70719 16000 71421 16028
rect 70719 15997 70731 16000
rect 70673 15991 70731 15997
rect 71409 15997 71421 16000
rect 71455 15997 71467 16031
rect 71409 15991 71467 15997
rect 66349 15963 66407 15969
rect 66349 15960 66361 15963
rect 65536 15932 66361 15960
rect 66349 15929 66361 15932
rect 66395 15929 66407 15963
rect 66349 15923 66407 15929
rect 47026 15892 47032 15904
rect 44100 15864 47032 15892
rect 33250 15855 33308 15861
rect 47026 15852 47032 15864
rect 47084 15852 47090 15904
rect 57054 15892 57060 15904
rect 57015 15864 57060 15892
rect 57054 15852 57060 15864
rect 57112 15852 57118 15904
rect 63497 15895 63555 15901
rect 63497 15861 63509 15895
rect 63543 15892 63555 15895
rect 64046 15892 64052 15904
rect 63543 15864 64052 15892
rect 63543 15861 63555 15864
rect 63497 15855 63555 15861
rect 64046 15852 64052 15864
rect 64104 15852 64110 15904
rect 65242 15892 65248 15904
rect 65203 15864 65248 15892
rect 65242 15852 65248 15864
rect 65300 15852 65306 15904
rect 69842 15852 69848 15904
rect 69900 15892 69906 15904
rect 70688 15892 70716 15991
rect 71682 15988 71688 16040
rect 71740 16028 71746 16040
rect 71869 16031 71927 16037
rect 71869 16028 71881 16031
rect 71740 16000 71881 16028
rect 71740 15988 71746 16000
rect 71869 15997 71881 16000
rect 71915 15997 71927 16031
rect 72050 16028 72056 16040
rect 71963 16000 72056 16028
rect 71869 15991 71927 15997
rect 72050 15988 72056 16000
rect 72108 16028 72114 16040
rect 73614 16028 73620 16040
rect 72108 16000 73620 16028
rect 72108 15988 72114 16000
rect 73614 15988 73620 16000
rect 73672 15988 73678 16040
rect 71133 15963 71191 15969
rect 71133 15929 71145 15963
rect 71179 15929 71191 15963
rect 71314 15960 71320 15972
rect 71275 15932 71320 15960
rect 71133 15923 71191 15929
rect 69900 15864 70716 15892
rect 71148 15892 71176 15923
rect 71314 15920 71320 15932
rect 71372 15920 71378 15972
rect 72326 15892 72332 15904
rect 71148 15864 72332 15892
rect 69900 15852 69906 15864
rect 72326 15852 72332 15864
rect 72384 15852 72390 15904
rect 1104 15802 178848 15824
rect 1104 15750 19606 15802
rect 19658 15750 19670 15802
rect 19722 15750 19734 15802
rect 19786 15750 19798 15802
rect 19850 15750 50326 15802
rect 50378 15750 50390 15802
rect 50442 15750 50454 15802
rect 50506 15750 50518 15802
rect 50570 15750 81046 15802
rect 81098 15750 81110 15802
rect 81162 15750 81174 15802
rect 81226 15750 81238 15802
rect 81290 15750 111766 15802
rect 111818 15750 111830 15802
rect 111882 15750 111894 15802
rect 111946 15750 111958 15802
rect 112010 15750 142486 15802
rect 142538 15750 142550 15802
rect 142602 15750 142614 15802
rect 142666 15750 142678 15802
rect 142730 15750 173206 15802
rect 173258 15750 173270 15802
rect 173322 15750 173334 15802
rect 173386 15750 173398 15802
rect 173450 15750 178848 15802
rect 1104 15728 178848 15750
rect 28994 15648 29000 15700
rect 29052 15688 29058 15700
rect 29273 15691 29331 15697
rect 29273 15688 29285 15691
rect 29052 15660 29285 15688
rect 29052 15648 29058 15660
rect 29273 15657 29285 15660
rect 29319 15657 29331 15691
rect 29273 15651 29331 15657
rect 31846 15648 31852 15700
rect 31904 15688 31910 15700
rect 31941 15691 31999 15697
rect 31941 15688 31953 15691
rect 31904 15660 31953 15688
rect 31904 15648 31910 15660
rect 31941 15657 31953 15660
rect 31987 15657 31999 15691
rect 56870 15688 56876 15700
rect 56831 15660 56876 15688
rect 31941 15651 31999 15657
rect 56870 15648 56876 15660
rect 56928 15648 56934 15700
rect 62669 15691 62727 15697
rect 62669 15657 62681 15691
rect 62715 15688 62727 15691
rect 63586 15688 63592 15700
rect 62715 15660 63592 15688
rect 62715 15657 62727 15660
rect 62669 15651 62727 15657
rect 63586 15648 63592 15660
rect 63644 15648 63650 15700
rect 70213 15691 70271 15697
rect 70213 15657 70225 15691
rect 70259 15688 70271 15691
rect 70486 15688 70492 15700
rect 70259 15660 70492 15688
rect 70259 15657 70271 15660
rect 70213 15651 70271 15657
rect 70486 15648 70492 15660
rect 70544 15648 70550 15700
rect 71133 15691 71191 15697
rect 71133 15657 71145 15691
rect 71179 15688 71191 15691
rect 72050 15688 72056 15700
rect 71179 15660 72056 15688
rect 71179 15657 71191 15660
rect 71133 15651 71191 15657
rect 72050 15648 72056 15660
rect 72108 15648 72114 15700
rect 32030 15620 32036 15632
rect 31864 15592 32036 15620
rect 29086 15512 29092 15564
rect 29144 15552 29150 15564
rect 29181 15555 29239 15561
rect 29181 15552 29193 15555
rect 29144 15524 29193 15552
rect 29144 15512 29150 15524
rect 29181 15521 29193 15524
rect 29227 15552 29239 15555
rect 30006 15552 30012 15564
rect 29227 15524 30012 15552
rect 29227 15521 29239 15524
rect 29181 15515 29239 15521
rect 30006 15512 30012 15524
rect 30064 15512 30070 15564
rect 31864 15561 31892 15592
rect 32030 15580 32036 15592
rect 32088 15580 32094 15632
rect 56686 15620 56692 15632
rect 56647 15592 56692 15620
rect 56686 15580 56692 15592
rect 56744 15580 56750 15632
rect 62485 15623 62543 15629
rect 62485 15589 62497 15623
rect 62531 15620 62543 15623
rect 70949 15623 71007 15629
rect 62531 15592 64092 15620
rect 62531 15589 62543 15592
rect 62485 15583 62543 15589
rect 64064 15564 64092 15592
rect 69124 15592 70256 15620
rect 31849 15555 31907 15561
rect 31849 15521 31861 15555
rect 31895 15521 31907 15555
rect 33686 15552 33692 15564
rect 33647 15524 33692 15552
rect 31849 15515 31907 15521
rect 33686 15512 33692 15524
rect 33744 15512 33750 15564
rect 33873 15555 33931 15561
rect 33873 15521 33885 15555
rect 33919 15552 33931 15555
rect 34514 15552 34520 15564
rect 33919 15524 34520 15552
rect 33919 15521 33931 15524
rect 33873 15515 33931 15521
rect 34514 15512 34520 15524
rect 34572 15512 34578 15564
rect 56962 15552 56968 15564
rect 56923 15524 56968 15552
rect 56962 15512 56968 15524
rect 57020 15512 57026 15564
rect 59722 15512 59728 15564
rect 59780 15552 59786 15564
rect 62761 15555 62819 15561
rect 59780 15524 62620 15552
rect 59780 15512 59786 15524
rect 29457 15487 29515 15493
rect 29457 15453 29469 15487
rect 29503 15484 29515 15487
rect 31202 15484 31208 15496
rect 29503 15456 31208 15484
rect 29503 15453 29515 15456
rect 29457 15447 29515 15453
rect 31202 15444 31208 15456
rect 31260 15484 31266 15496
rect 32033 15487 32091 15493
rect 32033 15484 32045 15487
rect 31260 15456 32045 15484
rect 31260 15444 31266 15456
rect 32033 15453 32045 15456
rect 32079 15453 32091 15487
rect 62592 15484 62620 15524
rect 62761 15521 62773 15555
rect 62807 15552 62819 15555
rect 63494 15552 63500 15564
rect 62807 15524 63500 15552
rect 62807 15521 62819 15524
rect 62761 15515 62819 15521
rect 62776 15484 62804 15515
rect 63494 15512 63500 15524
rect 63552 15512 63558 15564
rect 63865 15555 63923 15561
rect 63865 15521 63877 15555
rect 63911 15521 63923 15555
rect 64046 15552 64052 15564
rect 64007 15524 64052 15552
rect 63865 15515 63923 15521
rect 62592 15456 62804 15484
rect 32033 15447 32091 15453
rect 63880 15416 63908 15515
rect 64046 15512 64052 15524
rect 64104 15512 64110 15564
rect 64141 15555 64199 15561
rect 64141 15521 64153 15555
rect 64187 15552 64199 15555
rect 65978 15552 65984 15564
rect 64187 15524 65984 15552
rect 64187 15521 64199 15524
rect 64141 15515 64199 15521
rect 63954 15444 63960 15496
rect 64012 15484 64018 15496
rect 64156 15484 64184 15515
rect 65978 15512 65984 15524
rect 66036 15512 66042 15564
rect 69124 15561 69152 15592
rect 70228 15564 70256 15592
rect 70949 15589 70961 15623
rect 70995 15620 71007 15623
rect 71866 15620 71872 15632
rect 70995 15592 71872 15620
rect 70995 15589 71007 15592
rect 70949 15583 71007 15589
rect 71866 15580 71872 15592
rect 71924 15580 71930 15632
rect 69109 15555 69167 15561
rect 69109 15521 69121 15555
rect 69155 15521 69167 15555
rect 69842 15552 69848 15564
rect 69803 15524 69848 15552
rect 69109 15515 69167 15521
rect 69842 15512 69848 15524
rect 69900 15512 69906 15564
rect 70210 15512 70216 15564
rect 70268 15552 70274 15564
rect 70305 15555 70363 15561
rect 70305 15552 70317 15555
rect 70268 15524 70317 15552
rect 70268 15512 70274 15524
rect 70305 15521 70317 15524
rect 70351 15521 70363 15555
rect 70305 15515 70363 15521
rect 71225 15555 71283 15561
rect 71225 15521 71237 15555
rect 71271 15552 71283 15555
rect 71682 15552 71688 15564
rect 71271 15524 71688 15552
rect 71271 15521 71283 15524
rect 71225 15515 71283 15521
rect 71682 15512 71688 15524
rect 71740 15512 71746 15564
rect 64012 15456 64184 15484
rect 64012 15444 64018 15456
rect 68922 15444 68928 15496
rect 68980 15484 68986 15496
rect 69293 15487 69351 15493
rect 69293 15484 69305 15487
rect 68980 15456 69305 15484
rect 68980 15444 68986 15456
rect 69293 15453 69305 15456
rect 69339 15453 69351 15487
rect 69293 15447 69351 15453
rect 69382 15444 69388 15496
rect 69440 15484 69446 15496
rect 72142 15484 72148 15496
rect 69440 15456 72148 15484
rect 69440 15444 69446 15456
rect 72142 15444 72148 15456
rect 72200 15444 72206 15496
rect 65702 15416 65708 15428
rect 63880 15388 65708 15416
rect 65702 15376 65708 15388
rect 65760 15376 65766 15428
rect 28810 15348 28816 15360
rect 28771 15320 28816 15348
rect 28810 15308 28816 15320
rect 28868 15308 28874 15360
rect 31478 15348 31484 15360
rect 31439 15320 31484 15348
rect 31478 15308 31484 15320
rect 31536 15308 31542 15360
rect 33689 15351 33747 15357
rect 33689 15317 33701 15351
rect 33735 15348 33747 15351
rect 34790 15348 34796 15360
rect 33735 15320 34796 15348
rect 33735 15317 33747 15320
rect 33689 15311 33747 15317
rect 34790 15308 34796 15320
rect 34848 15308 34854 15360
rect 55306 15308 55312 15360
rect 55364 15348 55370 15360
rect 56689 15351 56747 15357
rect 56689 15348 56701 15351
rect 55364 15320 56701 15348
rect 55364 15308 55370 15320
rect 56689 15317 56701 15320
rect 56735 15317 56747 15351
rect 62482 15348 62488 15360
rect 62443 15320 62488 15348
rect 56689 15311 56747 15317
rect 62482 15308 62488 15320
rect 62540 15308 62546 15360
rect 63678 15348 63684 15360
rect 63639 15320 63684 15348
rect 63678 15308 63684 15320
rect 63736 15308 63742 15360
rect 67634 15308 67640 15360
rect 67692 15348 67698 15360
rect 68925 15351 68983 15357
rect 68925 15348 68937 15351
rect 67692 15320 68937 15348
rect 67692 15308 67698 15320
rect 68925 15317 68937 15320
rect 68971 15317 68983 15351
rect 70026 15348 70032 15360
rect 69987 15320 70032 15348
rect 68925 15311 68983 15317
rect 70026 15308 70032 15320
rect 70084 15308 70090 15360
rect 70118 15308 70124 15360
rect 70176 15348 70182 15360
rect 70949 15351 71007 15357
rect 70949 15348 70961 15351
rect 70176 15320 70961 15348
rect 70176 15308 70182 15320
rect 70949 15317 70961 15320
rect 70995 15317 71007 15351
rect 70949 15311 71007 15317
rect 1104 15258 178848 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 34966 15258
rect 35018 15206 35030 15258
rect 35082 15206 35094 15258
rect 35146 15206 35158 15258
rect 35210 15206 65686 15258
rect 65738 15206 65750 15258
rect 65802 15206 65814 15258
rect 65866 15206 65878 15258
rect 65930 15206 96406 15258
rect 96458 15206 96470 15258
rect 96522 15206 96534 15258
rect 96586 15206 96598 15258
rect 96650 15206 127126 15258
rect 127178 15206 127190 15258
rect 127242 15206 127254 15258
rect 127306 15206 127318 15258
rect 127370 15206 157846 15258
rect 157898 15206 157910 15258
rect 157962 15206 157974 15258
rect 158026 15206 158038 15258
rect 158090 15206 178848 15258
rect 1104 15184 178848 15206
rect 30653 15079 30711 15085
rect 30653 15045 30665 15079
rect 30699 15076 30711 15079
rect 32490 15076 32496 15088
rect 30699 15048 32496 15076
rect 30699 15045 30711 15048
rect 30653 15039 30711 15045
rect 32490 15036 32496 15048
rect 32548 15036 32554 15088
rect 28902 14968 28908 15020
rect 28960 15008 28966 15020
rect 31113 15011 31171 15017
rect 31113 15008 31125 15011
rect 28960 14980 31125 15008
rect 28960 14968 28966 14980
rect 31113 14977 31125 14980
rect 31159 14977 31171 15011
rect 31113 14971 31171 14977
rect 31202 14968 31208 15020
rect 31260 15008 31266 15020
rect 31260 14980 31305 15008
rect 31260 14968 31266 14980
rect 63494 14968 63500 15020
rect 63552 15008 63558 15020
rect 65981 15011 66039 15017
rect 65981 15008 65993 15011
rect 63552 14980 65993 15008
rect 63552 14968 63558 14980
rect 65981 14977 65993 14980
rect 66027 14977 66039 15011
rect 65981 14971 66039 14977
rect 33502 14940 33508 14952
rect 33463 14912 33508 14940
rect 33502 14900 33508 14912
rect 33560 14900 33566 14952
rect 33778 14940 33784 14952
rect 33739 14912 33784 14940
rect 33778 14900 33784 14912
rect 33836 14900 33842 14952
rect 59538 14900 59544 14952
rect 59596 14940 59602 14952
rect 59909 14943 59967 14949
rect 59909 14940 59921 14943
rect 59596 14912 59921 14940
rect 59596 14900 59602 14912
rect 59909 14909 59921 14912
rect 59955 14909 59967 14943
rect 59909 14903 59967 14909
rect 65518 14900 65524 14952
rect 65576 14940 65582 14952
rect 65797 14943 65855 14949
rect 65797 14940 65809 14943
rect 65576 14912 65809 14940
rect 65576 14900 65582 14912
rect 65797 14909 65809 14912
rect 65843 14909 65855 14943
rect 68373 14943 68431 14949
rect 68373 14940 68385 14943
rect 65797 14903 65855 14909
rect 68020 14912 68385 14940
rect 35161 14875 35219 14881
rect 35161 14841 35173 14875
rect 35207 14872 35219 14875
rect 35342 14872 35348 14884
rect 35207 14844 35348 14872
rect 35207 14841 35219 14844
rect 35161 14835 35219 14841
rect 35342 14832 35348 14844
rect 35400 14832 35406 14884
rect 59722 14872 59728 14884
rect 59683 14844 59728 14872
rect 59722 14832 59728 14844
rect 59780 14832 59786 14884
rect 60090 14872 60096 14884
rect 60051 14844 60096 14872
rect 60090 14832 60096 14844
rect 60148 14832 60154 14884
rect 65613 14875 65671 14881
rect 65613 14841 65625 14875
rect 65659 14872 65671 14875
rect 66346 14872 66352 14884
rect 65659 14844 66352 14872
rect 65659 14841 65671 14844
rect 65613 14835 65671 14841
rect 66346 14832 66352 14844
rect 66404 14872 66410 14884
rect 68020 14872 68048 14912
rect 68373 14909 68385 14912
rect 68419 14909 68431 14943
rect 68373 14903 68431 14909
rect 68554 14900 68560 14952
rect 68612 14940 68618 14952
rect 68612 14912 70394 14940
rect 68612 14900 68618 14912
rect 66404 14844 68048 14872
rect 68097 14875 68155 14881
rect 66404 14832 66410 14844
rect 68097 14841 68109 14875
rect 68143 14872 68155 14875
rect 68922 14872 68928 14884
rect 68143 14844 68928 14872
rect 68143 14841 68155 14844
rect 68097 14835 68155 14841
rect 68922 14832 68928 14844
rect 68980 14832 68986 14884
rect 70366 14872 70394 14912
rect 73522 14872 73528 14884
rect 70366 14844 73528 14872
rect 73522 14832 73528 14844
rect 73580 14832 73586 14884
rect 31018 14804 31024 14816
rect 30931 14776 31024 14804
rect 31018 14764 31024 14776
rect 31076 14804 31082 14816
rect 32214 14804 32220 14816
rect 31076 14776 32220 14804
rect 31076 14764 31082 14776
rect 32214 14764 32220 14776
rect 32272 14764 32278 14816
rect 65518 14764 65524 14816
rect 65576 14804 65582 14816
rect 68195 14807 68253 14813
rect 68195 14804 68207 14807
rect 65576 14776 68207 14804
rect 65576 14764 65582 14776
rect 68195 14773 68207 14776
rect 68241 14773 68253 14807
rect 68195 14767 68253 14773
rect 68281 14807 68339 14813
rect 68281 14773 68293 14807
rect 68327 14804 68339 14807
rect 70394 14804 70400 14816
rect 68327 14776 70400 14804
rect 68327 14773 68339 14776
rect 68281 14767 68339 14773
rect 70394 14764 70400 14776
rect 70452 14764 70458 14816
rect 1104 14714 178848 14736
rect 1104 14662 19606 14714
rect 19658 14662 19670 14714
rect 19722 14662 19734 14714
rect 19786 14662 19798 14714
rect 19850 14662 50326 14714
rect 50378 14662 50390 14714
rect 50442 14662 50454 14714
rect 50506 14662 50518 14714
rect 50570 14662 81046 14714
rect 81098 14662 81110 14714
rect 81162 14662 81174 14714
rect 81226 14662 81238 14714
rect 81290 14662 111766 14714
rect 111818 14662 111830 14714
rect 111882 14662 111894 14714
rect 111946 14662 111958 14714
rect 112010 14662 142486 14714
rect 142538 14662 142550 14714
rect 142602 14662 142614 14714
rect 142666 14662 142678 14714
rect 142730 14662 173206 14714
rect 173258 14662 173270 14714
rect 173322 14662 173334 14714
rect 173386 14662 173398 14714
rect 173450 14662 178848 14714
rect 1104 14640 178848 14662
rect 33042 14560 33048 14612
rect 33100 14600 33106 14612
rect 33229 14603 33287 14609
rect 33229 14600 33241 14603
rect 33100 14572 33241 14600
rect 33100 14560 33106 14572
rect 33229 14569 33241 14572
rect 33275 14569 33287 14603
rect 33229 14563 33287 14569
rect 68649 14603 68707 14609
rect 68649 14569 68661 14603
rect 68695 14600 68707 14603
rect 70118 14600 70124 14612
rect 68695 14572 70124 14600
rect 68695 14569 68707 14572
rect 68649 14563 68707 14569
rect 70118 14560 70124 14572
rect 70176 14560 70182 14612
rect 31754 14492 31760 14544
rect 31812 14532 31818 14544
rect 31849 14535 31907 14541
rect 31849 14532 31861 14535
rect 31812 14504 31861 14532
rect 31812 14492 31818 14504
rect 31849 14501 31861 14504
rect 31895 14501 31907 14535
rect 34057 14535 34115 14541
rect 34057 14532 34069 14535
rect 31849 14495 31907 14501
rect 33060 14504 34069 14532
rect 31110 14464 31116 14476
rect 31071 14436 31116 14464
rect 31110 14424 31116 14436
rect 31168 14464 31174 14476
rect 33060 14464 33088 14504
rect 34057 14501 34069 14504
rect 34103 14532 34115 14535
rect 39666 14532 39672 14544
rect 34103 14504 39672 14532
rect 34103 14501 34115 14504
rect 34057 14495 34115 14501
rect 39666 14492 39672 14504
rect 39724 14532 39730 14544
rect 46845 14535 46903 14541
rect 46845 14532 46857 14535
rect 39724 14504 46857 14532
rect 39724 14492 39730 14504
rect 46845 14501 46857 14504
rect 46891 14532 46903 14535
rect 69845 14535 69903 14541
rect 46891 14504 51074 14532
rect 46891 14501 46903 14504
rect 46845 14495 46903 14501
rect 31168 14436 33088 14464
rect 31168 14424 31174 14436
rect 33134 14424 33140 14476
rect 33192 14464 33198 14476
rect 34606 14464 34612 14476
rect 33192 14436 34612 14464
rect 33192 14424 33198 14436
rect 34606 14424 34612 14436
rect 34664 14424 34670 14476
rect 51046 14464 51074 14504
rect 69845 14501 69857 14535
rect 69891 14532 69903 14535
rect 73890 14532 73896 14544
rect 69891 14504 73896 14532
rect 69891 14501 69903 14504
rect 69845 14495 69903 14501
rect 73890 14492 73896 14504
rect 73948 14492 73954 14544
rect 68554 14464 68560 14476
rect 51046 14436 55214 14464
rect 68515 14436 68560 14464
rect 31202 14356 31208 14408
rect 31260 14396 31266 14408
rect 33413 14399 33471 14405
rect 33413 14396 33425 14399
rect 31260 14368 33425 14396
rect 31260 14356 31266 14368
rect 33413 14365 33425 14368
rect 33459 14396 33471 14399
rect 33962 14396 33968 14408
rect 33459 14368 33968 14396
rect 33459 14365 33471 14368
rect 33413 14359 33471 14365
rect 33962 14356 33968 14368
rect 34020 14356 34026 14408
rect 55186 14340 55214 14436
rect 68554 14424 68560 14436
rect 68612 14424 68618 14476
rect 69750 14464 69756 14476
rect 69711 14436 69756 14464
rect 69750 14424 69756 14436
rect 69808 14464 69814 14476
rect 74350 14464 74356 14476
rect 69808 14436 74356 14464
rect 69808 14424 69814 14436
rect 74350 14424 74356 14436
rect 74408 14424 74414 14476
rect 68833 14399 68891 14405
rect 68833 14365 68845 14399
rect 68879 14396 68891 14399
rect 69106 14396 69112 14408
rect 68879 14368 69112 14396
rect 68879 14365 68891 14368
rect 68833 14359 68891 14365
rect 69106 14356 69112 14368
rect 69164 14356 69170 14408
rect 70029 14399 70087 14405
rect 70029 14365 70041 14399
rect 70075 14396 70087 14399
rect 70302 14396 70308 14408
rect 70075 14368 70308 14396
rect 70075 14365 70087 14368
rect 70029 14359 70087 14365
rect 70302 14356 70308 14368
rect 70360 14356 70366 14408
rect 34238 14328 34244 14340
rect 34199 14300 34244 14328
rect 34238 14288 34244 14300
rect 34296 14288 34302 14340
rect 55186 14300 55220 14340
rect 55214 14288 55220 14300
rect 55272 14328 55278 14340
rect 101306 14328 101312 14340
rect 55272 14300 101312 14328
rect 55272 14288 55278 14300
rect 101306 14288 101312 14300
rect 101364 14288 101370 14340
rect 32769 14263 32827 14269
rect 32769 14229 32781 14263
rect 32815 14260 32827 14263
rect 33134 14260 33140 14272
rect 32815 14232 33140 14260
rect 32815 14229 32827 14232
rect 32769 14223 32827 14229
rect 33134 14220 33140 14232
rect 33192 14220 33198 14272
rect 46934 14260 46940 14272
rect 46895 14232 46940 14260
rect 46934 14220 46940 14232
rect 46992 14220 46998 14272
rect 68186 14260 68192 14272
rect 68147 14232 68192 14260
rect 68186 14220 68192 14232
rect 68244 14220 68250 14272
rect 68278 14220 68284 14272
rect 68336 14260 68342 14272
rect 69385 14263 69443 14269
rect 69385 14260 69397 14263
rect 68336 14232 69397 14260
rect 68336 14220 68342 14232
rect 69385 14229 69397 14232
rect 69431 14229 69443 14263
rect 69385 14223 69443 14229
rect 1104 14170 178848 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 34966 14170
rect 35018 14118 35030 14170
rect 35082 14118 35094 14170
rect 35146 14118 35158 14170
rect 35210 14118 65686 14170
rect 65738 14118 65750 14170
rect 65802 14118 65814 14170
rect 65866 14118 65878 14170
rect 65930 14118 96406 14170
rect 96458 14118 96470 14170
rect 96522 14118 96534 14170
rect 96586 14118 96598 14170
rect 96650 14118 127126 14170
rect 127178 14118 127190 14170
rect 127242 14118 127254 14170
rect 127306 14118 127318 14170
rect 127370 14118 157846 14170
rect 157898 14118 157910 14170
rect 157962 14118 157974 14170
rect 158026 14118 158038 14170
rect 158090 14118 178848 14170
rect 1104 14096 178848 14118
rect 30006 14016 30012 14068
rect 30064 14056 30070 14068
rect 30469 14059 30527 14065
rect 30469 14056 30481 14059
rect 30064 14028 30481 14056
rect 30064 14016 30070 14028
rect 30469 14025 30481 14028
rect 30515 14025 30527 14059
rect 30469 14019 30527 14025
rect 40681 14059 40739 14065
rect 40681 14025 40693 14059
rect 40727 14056 40739 14059
rect 41138 14056 41144 14068
rect 40727 14028 41144 14056
rect 40727 14025 40739 14028
rect 40681 14019 40739 14025
rect 41138 14016 41144 14028
rect 41196 14016 41202 14068
rect 46845 14059 46903 14065
rect 46845 14025 46857 14059
rect 46891 14056 46903 14059
rect 48038 14056 48044 14068
rect 46891 14028 48044 14056
rect 46891 14025 46903 14028
rect 46845 14019 46903 14025
rect 48038 14016 48044 14028
rect 48096 14016 48102 14068
rect 57238 14016 57244 14068
rect 57296 14056 57302 14068
rect 60553 14059 60611 14065
rect 60553 14056 60565 14059
rect 57296 14028 60565 14056
rect 57296 14016 57302 14028
rect 60553 14025 60565 14028
rect 60599 14025 60611 14059
rect 60553 14019 60611 14025
rect 62390 14016 62396 14068
rect 62448 14056 62454 14068
rect 65061 14059 65119 14065
rect 65061 14056 65073 14059
rect 62448 14028 65073 14056
rect 62448 14016 62454 14028
rect 65061 14025 65073 14028
rect 65107 14025 65119 14059
rect 65061 14019 65119 14025
rect 33413 13991 33471 13997
rect 33413 13957 33425 13991
rect 33459 13988 33471 13991
rect 35250 13988 35256 14000
rect 33459 13960 35256 13988
rect 33459 13957 33471 13960
rect 33413 13951 33471 13957
rect 35250 13948 35256 13960
rect 35308 13948 35314 14000
rect 35897 13991 35955 13997
rect 35897 13957 35909 13991
rect 35943 13988 35955 13991
rect 36630 13988 36636 14000
rect 35943 13960 36636 13988
rect 35943 13957 35955 13960
rect 35897 13951 35955 13957
rect 36630 13948 36636 13960
rect 36688 13948 36694 14000
rect 38381 13991 38439 13997
rect 38381 13957 38393 13991
rect 38427 13988 38439 13991
rect 39574 13988 39580 14000
rect 38427 13960 39580 13988
rect 38427 13957 38439 13960
rect 38381 13951 38439 13957
rect 39574 13948 39580 13960
rect 39632 13948 39638 14000
rect 39684 13960 41368 13988
rect 29089 13923 29147 13929
rect 29089 13889 29101 13923
rect 29135 13920 29147 13923
rect 30834 13920 30840 13932
rect 29135 13892 30840 13920
rect 29135 13889 29147 13892
rect 29089 13883 29147 13889
rect 30834 13880 30840 13892
rect 30892 13880 30898 13932
rect 31938 13880 31944 13932
rect 31996 13920 32002 13932
rect 33873 13923 33931 13929
rect 33873 13920 33885 13923
rect 31996 13892 33885 13920
rect 31996 13880 32002 13892
rect 33873 13889 33885 13892
rect 33919 13889 33931 13923
rect 33873 13883 33931 13889
rect 34057 13923 34115 13929
rect 34057 13889 34069 13923
rect 34103 13889 34115 13923
rect 36354 13920 36360 13932
rect 36315 13892 36360 13920
rect 34057 13883 34115 13889
rect 29365 13855 29423 13861
rect 29365 13821 29377 13855
rect 29411 13852 29423 13855
rect 31662 13852 31668 13864
rect 29411 13824 31668 13852
rect 29411 13821 29423 13824
rect 29365 13815 29423 13821
rect 31662 13812 31668 13824
rect 31720 13812 31726 13864
rect 33962 13812 33968 13864
rect 34020 13852 34026 13864
rect 34072 13852 34100 13883
rect 36354 13880 36360 13892
rect 36412 13880 36418 13932
rect 36449 13923 36507 13929
rect 36449 13889 36461 13923
rect 36495 13889 36507 13923
rect 38838 13920 38844 13932
rect 38799 13892 38844 13920
rect 36449 13883 36507 13889
rect 36464 13852 36492 13883
rect 38838 13880 38844 13892
rect 38896 13880 38902 13932
rect 39025 13923 39083 13929
rect 39025 13889 39037 13923
rect 39071 13920 39083 13923
rect 39684 13920 39712 13960
rect 39071 13892 39712 13920
rect 39071 13889 39083 13892
rect 39025 13883 39083 13889
rect 39040 13852 39068 13883
rect 40954 13880 40960 13932
rect 41012 13920 41018 13932
rect 41340 13929 41368 13960
rect 47854 13948 47860 14000
rect 47912 13988 47918 14000
rect 48777 13991 48835 13997
rect 48777 13988 48789 13991
rect 47912 13960 48789 13988
rect 47912 13948 47918 13960
rect 48777 13957 48789 13960
rect 48823 13957 48835 13991
rect 48777 13951 48835 13957
rect 56594 13948 56600 14000
rect 56652 13988 56658 14000
rect 59265 13991 59323 13997
rect 59265 13988 59277 13991
rect 56652 13960 59277 13988
rect 56652 13948 56658 13960
rect 59265 13957 59277 13960
rect 59311 13957 59323 13991
rect 60090 13988 60096 14000
rect 59265 13951 59323 13957
rect 59740 13960 60096 13988
rect 41141 13923 41199 13929
rect 41141 13920 41153 13923
rect 41012 13892 41153 13920
rect 41012 13880 41018 13892
rect 41141 13889 41153 13892
rect 41187 13889 41199 13923
rect 41141 13883 41199 13889
rect 41325 13923 41383 13929
rect 41325 13889 41337 13923
rect 41371 13920 41383 13923
rect 43622 13920 43628 13932
rect 41371 13892 43628 13920
rect 41371 13889 41383 13892
rect 41325 13883 41383 13889
rect 43622 13880 43628 13892
rect 43680 13920 43686 13932
rect 44913 13923 44971 13929
rect 44913 13920 44925 13923
rect 43680 13892 44925 13920
rect 43680 13880 43686 13892
rect 44913 13889 44925 13892
rect 44959 13889 44971 13923
rect 44913 13883 44971 13889
rect 47210 13880 47216 13932
rect 47268 13920 47274 13932
rect 47305 13923 47363 13929
rect 47305 13920 47317 13923
rect 47268 13892 47317 13920
rect 47268 13880 47274 13892
rect 47305 13889 47317 13892
rect 47351 13889 47363 13923
rect 47305 13883 47363 13889
rect 47489 13923 47547 13929
rect 47489 13889 47501 13923
rect 47535 13889 47547 13923
rect 47489 13883 47547 13889
rect 39666 13852 39672 13864
rect 34020 13824 36492 13852
rect 34020 13812 34026 13824
rect 35894 13744 35900 13796
rect 35952 13784 35958 13796
rect 36265 13787 36323 13793
rect 36265 13784 36277 13787
rect 35952 13756 36277 13784
rect 35952 13744 35958 13756
rect 36265 13753 36277 13756
rect 36311 13753 36323 13787
rect 36464 13784 36492 13824
rect 36648 13824 39068 13852
rect 39627 13824 39672 13852
rect 36538 13784 36544 13796
rect 36451 13756 36544 13784
rect 36265 13747 36323 13753
rect 36538 13744 36544 13756
rect 36596 13784 36602 13796
rect 36648 13784 36676 13824
rect 39666 13812 39672 13824
rect 39724 13812 39730 13864
rect 39850 13852 39856 13864
rect 39811 13824 39856 13852
rect 39850 13812 39856 13824
rect 39908 13812 39914 13864
rect 44729 13855 44787 13861
rect 44729 13821 44741 13855
rect 44775 13852 44787 13855
rect 44818 13852 44824 13864
rect 44775 13824 44824 13852
rect 44775 13821 44787 13824
rect 44729 13815 44787 13821
rect 44818 13812 44824 13824
rect 44876 13852 44882 13864
rect 47026 13852 47032 13864
rect 44876 13824 47032 13852
rect 44876 13812 44882 13824
rect 47026 13812 47032 13824
rect 47084 13852 47090 13864
rect 47504 13852 47532 13883
rect 49050 13880 49056 13932
rect 49108 13920 49114 13932
rect 49237 13923 49295 13929
rect 49237 13920 49249 13923
rect 49108 13892 49249 13920
rect 49108 13880 49114 13892
rect 49237 13889 49249 13892
rect 49283 13889 49295 13923
rect 49418 13920 49424 13932
rect 49379 13892 49424 13920
rect 49237 13883 49295 13889
rect 49418 13880 49424 13892
rect 49476 13880 49482 13932
rect 59740 13929 59768 13960
rect 60090 13948 60096 13960
rect 60148 13948 60154 14000
rect 64966 13948 64972 14000
rect 65024 13988 65030 14000
rect 66257 13991 66315 13997
rect 66257 13988 66269 13991
rect 65024 13960 66269 13988
rect 65024 13948 65030 13960
rect 66257 13957 66269 13960
rect 66303 13957 66315 13991
rect 66257 13951 66315 13957
rect 66898 13948 66904 14000
rect 66956 13988 66962 14000
rect 68097 13991 68155 13997
rect 68097 13988 68109 13991
rect 66956 13960 68109 13988
rect 66956 13948 66962 13960
rect 68097 13957 68109 13960
rect 68143 13957 68155 13991
rect 68097 13951 68155 13957
rect 69566 13948 69572 14000
rect 69624 13988 69630 14000
rect 69753 13991 69811 13997
rect 69753 13988 69765 13991
rect 69624 13960 69765 13988
rect 69624 13948 69630 13960
rect 69753 13957 69765 13960
rect 69799 13957 69811 13991
rect 70210 13988 70216 14000
rect 69753 13951 69811 13957
rect 69860 13960 70216 13988
rect 59725 13923 59783 13929
rect 59725 13889 59737 13923
rect 59771 13889 59783 13923
rect 59906 13920 59912 13932
rect 59819 13892 59912 13920
rect 59725 13883 59783 13889
rect 59906 13880 59912 13892
rect 59964 13920 59970 13932
rect 61197 13923 61255 13929
rect 61197 13920 61209 13923
rect 59964 13892 61209 13920
rect 59964 13880 59970 13892
rect 61197 13889 61209 13892
rect 61243 13920 61255 13923
rect 65518 13920 65524 13932
rect 61243 13892 63448 13920
rect 65479 13892 65524 13920
rect 61243 13889 61255 13892
rect 61197 13883 61255 13889
rect 49436 13852 49464 13880
rect 63420 13864 63448 13892
rect 65518 13880 65524 13892
rect 65576 13880 65582 13932
rect 65705 13923 65763 13929
rect 65705 13889 65717 13923
rect 65751 13920 65763 13923
rect 66809 13923 66867 13929
rect 66809 13920 66821 13923
rect 65751 13892 66821 13920
rect 65751 13889 65763 13892
rect 65705 13883 65763 13889
rect 66809 13889 66821 13892
rect 66855 13920 66867 13923
rect 68741 13923 68799 13929
rect 68741 13920 68753 13923
rect 66855 13892 68753 13920
rect 66855 13889 66867 13892
rect 66809 13883 66867 13889
rect 68741 13889 68753 13892
rect 68787 13920 68799 13923
rect 69106 13920 69112 13932
rect 68787 13892 69112 13920
rect 68787 13889 68799 13892
rect 68741 13883 68799 13889
rect 47084 13824 49464 13852
rect 47084 13812 47090 13824
rect 55214 13812 55220 13864
rect 55272 13852 55278 13864
rect 55398 13852 55404 13864
rect 55272 13824 55317 13852
rect 55359 13824 55404 13852
rect 55272 13812 55278 13824
rect 55398 13812 55404 13824
rect 55456 13812 55462 13864
rect 56965 13855 57023 13861
rect 56965 13821 56977 13855
rect 57011 13852 57023 13855
rect 60366 13852 60372 13864
rect 57011 13824 60372 13852
rect 57011 13821 57023 13824
rect 56965 13815 57023 13821
rect 60366 13812 60372 13824
rect 60424 13812 60430 13864
rect 61013 13855 61071 13861
rect 61013 13821 61025 13855
rect 61059 13852 61071 13855
rect 62482 13852 62488 13864
rect 61059 13824 62488 13852
rect 61059 13821 61071 13824
rect 61013 13815 61071 13821
rect 62482 13812 62488 13824
rect 62540 13812 62546 13864
rect 63402 13812 63408 13864
rect 63460 13852 63466 13864
rect 65720 13852 65748 13883
rect 69106 13880 69112 13892
rect 69164 13920 69170 13932
rect 69860 13920 69888 13960
rect 70210 13948 70216 13960
rect 70268 13948 70274 14000
rect 70302 13920 70308 13932
rect 69164 13892 69888 13920
rect 70263 13892 70308 13920
rect 69164 13880 69170 13892
rect 70302 13880 70308 13892
rect 70360 13880 70366 13932
rect 63460 13824 65748 13852
rect 66717 13855 66775 13861
rect 63460 13812 63466 13824
rect 66717 13821 66729 13855
rect 66763 13852 66775 13855
rect 67634 13852 67640 13864
rect 66763 13824 67640 13852
rect 66763 13821 66775 13824
rect 66717 13815 66775 13821
rect 67634 13812 67640 13824
rect 67692 13812 67698 13864
rect 68557 13855 68615 13861
rect 68557 13821 68569 13855
rect 68603 13852 68615 13855
rect 69014 13852 69020 13864
rect 68603 13824 69020 13852
rect 68603 13821 68615 13824
rect 68557 13815 68615 13821
rect 69014 13812 69020 13824
rect 69072 13812 69078 13864
rect 69842 13812 69848 13864
rect 69900 13852 69906 13864
rect 70121 13855 70179 13861
rect 70121 13852 70133 13855
rect 69900 13824 70133 13852
rect 69900 13812 69906 13824
rect 70121 13821 70133 13824
rect 70167 13821 70179 13855
rect 70121 13815 70179 13821
rect 70213 13855 70271 13861
rect 70213 13821 70225 13855
rect 70259 13852 70271 13855
rect 72510 13852 72516 13864
rect 70259 13824 72516 13852
rect 70259 13821 70271 13824
rect 70213 13815 70271 13821
rect 72510 13812 72516 13824
rect 72568 13812 72574 13864
rect 38746 13784 38752 13796
rect 36596 13756 36676 13784
rect 38707 13756 38752 13784
rect 36596 13744 36602 13756
rect 38746 13744 38752 13756
rect 38804 13744 38810 13796
rect 41049 13787 41107 13793
rect 41049 13753 41061 13787
rect 41095 13784 41107 13787
rect 41414 13784 41420 13796
rect 41095 13756 41420 13784
rect 41095 13753 41107 13756
rect 41049 13747 41107 13753
rect 41414 13744 41420 13756
rect 41472 13744 41478 13796
rect 47213 13787 47271 13793
rect 47213 13753 47225 13787
rect 47259 13784 47271 13787
rect 47762 13784 47768 13796
rect 47259 13756 47768 13784
rect 47259 13753 47271 13756
rect 47213 13747 47271 13753
rect 47762 13744 47768 13756
rect 47820 13784 47826 13796
rect 48406 13784 48412 13796
rect 47820 13756 48412 13784
rect 47820 13744 47826 13756
rect 48406 13744 48412 13756
rect 48464 13744 48470 13796
rect 33781 13719 33839 13725
rect 33781 13685 33793 13719
rect 33827 13716 33839 13719
rect 35342 13716 35348 13728
rect 33827 13688 35348 13716
rect 33827 13685 33839 13688
rect 33781 13679 33839 13685
rect 35342 13676 35348 13688
rect 35400 13716 35406 13728
rect 40126 13716 40132 13728
rect 35400 13688 40132 13716
rect 35400 13676 35406 13688
rect 40126 13676 40132 13688
rect 40184 13676 40190 13728
rect 49145 13719 49203 13725
rect 49145 13685 49157 13719
rect 49191 13716 49203 13719
rect 49510 13716 49516 13728
rect 49191 13688 49516 13716
rect 49191 13685 49203 13688
rect 49145 13679 49203 13685
rect 49510 13676 49516 13688
rect 49568 13716 49574 13728
rect 50614 13716 50620 13728
rect 49568 13688 50620 13716
rect 49568 13676 49574 13688
rect 50614 13676 50620 13688
rect 50672 13676 50678 13728
rect 56686 13676 56692 13728
rect 56744 13716 56750 13728
rect 56781 13719 56839 13725
rect 56781 13716 56793 13719
rect 56744 13688 56793 13716
rect 56744 13676 56750 13688
rect 56781 13685 56793 13688
rect 56827 13685 56839 13719
rect 56781 13679 56839 13685
rect 59633 13719 59691 13725
rect 59633 13685 59645 13719
rect 59679 13716 59691 13719
rect 60826 13716 60832 13728
rect 59679 13688 60832 13716
rect 59679 13685 59691 13688
rect 59633 13679 59691 13685
rect 60826 13676 60832 13688
rect 60884 13676 60890 13728
rect 60921 13719 60979 13725
rect 60921 13685 60933 13719
rect 60967 13716 60979 13719
rect 62482 13716 62488 13728
rect 60967 13688 62488 13716
rect 60967 13685 60979 13688
rect 60921 13679 60979 13685
rect 62482 13676 62488 13688
rect 62540 13716 62546 13728
rect 65150 13716 65156 13728
rect 62540 13688 65156 13716
rect 62540 13676 62546 13688
rect 65150 13676 65156 13688
rect 65208 13676 65214 13728
rect 65429 13719 65487 13725
rect 65429 13685 65441 13719
rect 65475 13716 65487 13719
rect 66254 13716 66260 13728
rect 65475 13688 66260 13716
rect 65475 13685 65487 13688
rect 65429 13679 65487 13685
rect 66254 13676 66260 13688
rect 66312 13676 66318 13728
rect 66625 13719 66683 13725
rect 66625 13685 66637 13719
rect 66671 13716 66683 13719
rect 68002 13716 68008 13728
rect 66671 13688 68008 13716
rect 66671 13685 66683 13688
rect 66625 13679 66683 13685
rect 68002 13676 68008 13688
rect 68060 13676 68066 13728
rect 68465 13719 68523 13725
rect 68465 13685 68477 13719
rect 68511 13716 68523 13719
rect 68646 13716 68652 13728
rect 68511 13688 68652 13716
rect 68511 13685 68523 13688
rect 68465 13679 68523 13685
rect 68646 13676 68652 13688
rect 68704 13676 68710 13728
rect 1104 13626 178848 13648
rect 1104 13574 19606 13626
rect 19658 13574 19670 13626
rect 19722 13574 19734 13626
rect 19786 13574 19798 13626
rect 19850 13574 50326 13626
rect 50378 13574 50390 13626
rect 50442 13574 50454 13626
rect 50506 13574 50518 13626
rect 50570 13574 81046 13626
rect 81098 13574 81110 13626
rect 81162 13574 81174 13626
rect 81226 13574 81238 13626
rect 81290 13574 111766 13626
rect 111818 13574 111830 13626
rect 111882 13574 111894 13626
rect 111946 13574 111958 13626
rect 112010 13574 142486 13626
rect 142538 13574 142550 13626
rect 142602 13574 142614 13626
rect 142666 13574 142678 13626
rect 142730 13574 173206 13626
rect 173258 13574 173270 13626
rect 173322 13574 173334 13626
rect 173386 13574 173398 13626
rect 173450 13574 178848 13626
rect 1104 13552 178848 13574
rect 32214 13512 32220 13524
rect 32175 13484 32220 13512
rect 32214 13472 32220 13484
rect 32272 13472 32278 13524
rect 33413 13515 33471 13521
rect 33413 13481 33425 13515
rect 33459 13512 33471 13515
rect 38194 13512 38200 13524
rect 33459 13484 38200 13512
rect 33459 13481 33471 13484
rect 33413 13475 33471 13481
rect 38194 13472 38200 13484
rect 38252 13472 38258 13524
rect 42794 13472 42800 13524
rect 42852 13512 42858 13524
rect 43533 13515 43591 13521
rect 43533 13512 43545 13515
rect 42852 13484 43545 13512
rect 42852 13472 42858 13484
rect 43533 13481 43545 13484
rect 43579 13481 43591 13515
rect 44726 13512 44732 13524
rect 44687 13484 44732 13512
rect 43533 13475 43591 13481
rect 44726 13472 44732 13484
rect 44784 13472 44790 13524
rect 47578 13512 47584 13524
rect 47539 13484 47584 13512
rect 47578 13472 47584 13484
rect 47636 13472 47642 13524
rect 51905 13515 51963 13521
rect 51905 13481 51917 13515
rect 51951 13512 51963 13515
rect 52730 13512 52736 13524
rect 51951 13484 52736 13512
rect 51951 13481 51963 13484
rect 51905 13475 51963 13481
rect 52730 13472 52736 13484
rect 52788 13472 52794 13524
rect 55306 13512 55312 13524
rect 55267 13484 55312 13512
rect 55306 13472 55312 13484
rect 55364 13472 55370 13524
rect 57609 13515 57667 13521
rect 57609 13481 57621 13515
rect 57655 13512 57667 13515
rect 58250 13512 58256 13524
rect 57655 13484 58256 13512
rect 57655 13481 57667 13484
rect 57609 13475 57667 13481
rect 58250 13472 58256 13484
rect 58308 13472 58314 13524
rect 59906 13512 59912 13524
rect 58360 13484 59912 13512
rect 42613 13447 42671 13453
rect 33152 13416 34008 13444
rect 30834 13376 30840 13388
rect 30795 13348 30840 13376
rect 30834 13336 30840 13348
rect 30892 13336 30898 13388
rect 33152 13385 33180 13416
rect 33980 13388 34008 13416
rect 42613 13413 42625 13447
rect 42659 13444 42671 13447
rect 43438 13444 43444 13456
rect 42659 13416 43444 13444
rect 42659 13413 42671 13416
rect 42613 13407 42671 13413
rect 42812 13388 42840 13416
rect 43438 13404 43444 13416
rect 43496 13404 43502 13456
rect 44634 13444 44640 13456
rect 44595 13416 44640 13444
rect 44634 13404 44640 13416
rect 44692 13404 44698 13456
rect 58360 13444 58388 13484
rect 59906 13472 59912 13484
rect 59964 13472 59970 13524
rect 63313 13515 63371 13521
rect 63313 13481 63325 13515
rect 63359 13512 63371 13515
rect 65242 13512 65248 13524
rect 63359 13484 65248 13512
rect 63359 13481 63371 13484
rect 63313 13475 63371 13481
rect 65242 13472 65248 13484
rect 65300 13472 65306 13524
rect 66254 13472 66260 13524
rect 66312 13512 66318 13524
rect 71225 13515 71283 13521
rect 66312 13484 70394 13512
rect 66312 13472 66318 13484
rect 57900 13416 58388 13444
rect 70366 13444 70394 13484
rect 71225 13481 71237 13515
rect 71271 13512 71283 13515
rect 72418 13512 72424 13524
rect 71271 13484 72424 13512
rect 71271 13481 71283 13484
rect 71225 13475 71283 13481
rect 72418 13472 72424 13484
rect 72476 13472 72482 13524
rect 72234 13444 72240 13456
rect 70366 13416 72240 13444
rect 33137 13379 33195 13385
rect 33137 13345 33149 13379
rect 33183 13345 33195 13379
rect 33137 13339 33195 13345
rect 33226 13336 33232 13388
rect 33284 13376 33290 13388
rect 33597 13379 33655 13385
rect 33597 13376 33609 13379
rect 33284 13348 33609 13376
rect 33284 13336 33290 13348
rect 33597 13345 33609 13348
rect 33643 13345 33655 13379
rect 33962 13376 33968 13388
rect 33923 13348 33968 13376
rect 33597 13339 33655 13345
rect 31113 13311 31171 13317
rect 31113 13277 31125 13311
rect 31159 13308 31171 13311
rect 33045 13311 33103 13317
rect 31159 13280 32536 13308
rect 31159 13277 31171 13280
rect 31113 13271 31171 13277
rect 32508 13240 32536 13280
rect 33045 13277 33057 13311
rect 33091 13308 33103 13311
rect 33244 13308 33272 13336
rect 33091 13280 33272 13308
rect 33612 13308 33640 13339
rect 33962 13336 33968 13348
rect 34020 13336 34026 13388
rect 42794 13336 42800 13388
rect 42852 13336 42858 13388
rect 45462 13336 45468 13388
rect 45520 13376 45526 13388
rect 46201 13379 46259 13385
rect 46201 13376 46213 13379
rect 45520 13348 46213 13376
rect 45520 13336 45526 13348
rect 46201 13345 46213 13348
rect 46247 13376 46259 13379
rect 48501 13379 48559 13385
rect 46247 13348 46612 13376
rect 46247 13345 46259 13348
rect 46201 13339 46259 13345
rect 34514 13308 34520 13320
rect 33612 13280 34520 13308
rect 33091 13277 33103 13280
rect 33045 13271 33103 13277
rect 34514 13268 34520 13280
rect 34572 13268 34578 13320
rect 36170 13268 36176 13320
rect 36228 13308 36234 13320
rect 36265 13311 36323 13317
rect 36265 13308 36277 13311
rect 36228 13280 36277 13308
rect 36228 13268 36234 13280
rect 36265 13277 36277 13280
rect 36311 13277 36323 13311
rect 36265 13271 36323 13277
rect 36541 13311 36599 13317
rect 36541 13277 36553 13311
rect 36587 13308 36599 13311
rect 38562 13308 38568 13320
rect 36587 13280 38568 13308
rect 36587 13277 36599 13280
rect 36541 13271 36599 13277
rect 38562 13268 38568 13280
rect 38620 13268 38626 13320
rect 40954 13308 40960 13320
rect 40915 13280 40960 13308
rect 40954 13268 40960 13280
rect 41012 13268 41018 13320
rect 41233 13311 41291 13317
rect 41233 13277 41245 13311
rect 41279 13308 41291 13311
rect 41598 13308 41604 13320
rect 41279 13280 41604 13308
rect 41279 13277 41291 13280
rect 41233 13271 41291 13277
rect 41598 13268 41604 13280
rect 41656 13268 41662 13320
rect 43622 13308 43628 13320
rect 43583 13280 43628 13308
rect 43622 13268 43628 13280
rect 43680 13268 43686 13320
rect 44818 13308 44824 13320
rect 44779 13280 44824 13308
rect 44818 13268 44824 13280
rect 44876 13268 44882 13320
rect 46474 13308 46480 13320
rect 46435 13280 46480 13308
rect 46474 13268 46480 13280
rect 46532 13268 46538 13320
rect 46584 13308 46612 13348
rect 48501 13345 48513 13379
rect 48547 13376 48559 13379
rect 48774 13376 48780 13388
rect 48547 13348 48780 13376
rect 48547 13345 48559 13348
rect 48501 13339 48559 13345
rect 48774 13336 48780 13348
rect 48832 13336 48838 13388
rect 51813 13379 51871 13385
rect 51813 13345 51825 13379
rect 51859 13376 51871 13379
rect 52270 13376 52276 13388
rect 51859 13348 52276 13376
rect 51859 13345 51871 13348
rect 51813 13339 51871 13345
rect 52270 13336 52276 13348
rect 52328 13376 52334 13388
rect 53190 13376 53196 13388
rect 52328 13348 53196 13376
rect 52328 13336 52334 13348
rect 53190 13336 53196 13348
rect 53248 13336 53254 13388
rect 55214 13336 55220 13388
rect 55272 13376 55278 13388
rect 57146 13376 57152 13388
rect 55272 13348 57152 13376
rect 55272 13336 55278 13348
rect 57146 13336 57152 13348
rect 57204 13336 57210 13388
rect 57514 13376 57520 13388
rect 57475 13348 57520 13376
rect 57514 13336 57520 13348
rect 57572 13336 57578 13388
rect 48869 13311 48927 13317
rect 48869 13308 48881 13311
rect 46584 13280 48881 13308
rect 48869 13277 48881 13280
rect 48915 13277 48927 13311
rect 48869 13271 48927 13277
rect 49418 13268 49424 13320
rect 49476 13308 49482 13320
rect 52089 13311 52147 13317
rect 52089 13308 52101 13311
rect 49476 13280 52101 13308
rect 49476 13268 49482 13280
rect 52089 13277 52101 13280
rect 52135 13308 52147 13311
rect 55493 13311 55551 13317
rect 55493 13308 55505 13311
rect 52135 13280 55505 13308
rect 52135 13277 52147 13280
rect 52089 13271 52147 13277
rect 55493 13277 55505 13280
rect 55539 13308 55551 13311
rect 57606 13308 57612 13320
rect 55539 13280 57612 13308
rect 55539 13277 55551 13280
rect 55493 13271 55551 13277
rect 57606 13268 57612 13280
rect 57664 13308 57670 13320
rect 57793 13311 57851 13317
rect 57793 13308 57805 13311
rect 57664 13280 57805 13308
rect 57664 13268 57670 13280
rect 57793 13277 57805 13280
rect 57839 13308 57851 13311
rect 57900 13308 57928 13416
rect 72234 13404 72240 13416
rect 72292 13404 72298 13456
rect 57974 13336 57980 13388
rect 58032 13376 58038 13388
rect 58621 13379 58679 13385
rect 58621 13376 58633 13379
rect 58032 13348 58633 13376
rect 58032 13336 58038 13348
rect 58621 13345 58633 13348
rect 58667 13345 58679 13379
rect 58621 13339 58679 13345
rect 63221 13379 63279 13385
rect 63221 13345 63233 13379
rect 63267 13376 63279 13379
rect 65334 13376 65340 13388
rect 63267 13348 65340 13376
rect 63267 13345 63279 13348
rect 63221 13339 63279 13345
rect 65334 13336 65340 13348
rect 65392 13336 65398 13388
rect 69477 13379 69535 13385
rect 69477 13345 69489 13379
rect 69523 13376 69535 13379
rect 70302 13376 70308 13388
rect 69523 13348 70308 13376
rect 69523 13345 69535 13348
rect 69477 13339 69535 13345
rect 70302 13336 70308 13348
rect 70360 13376 70366 13388
rect 71130 13376 71136 13388
rect 70360 13336 70394 13376
rect 71043 13348 71136 13376
rect 71130 13336 71136 13348
rect 71188 13376 71194 13388
rect 73062 13376 73068 13388
rect 71188 13348 73068 13376
rect 71188 13336 71194 13348
rect 73062 13336 73068 13348
rect 73120 13336 73126 13388
rect 57839 13280 57928 13308
rect 58345 13311 58403 13317
rect 57839 13277 57851 13280
rect 57793 13271 57851 13277
rect 58345 13277 58357 13311
rect 58391 13277 58403 13311
rect 58345 13271 58403 13277
rect 60001 13311 60059 13317
rect 60001 13277 60013 13311
rect 60047 13308 60059 13311
rect 60826 13308 60832 13320
rect 60047 13280 60832 13308
rect 60047 13277 60059 13280
rect 60001 13271 60059 13277
rect 33226 13240 33232 13252
rect 32508 13212 33232 13240
rect 33226 13200 33232 13212
rect 33284 13200 33290 13252
rect 41966 13200 41972 13252
rect 42024 13240 42030 13252
rect 43073 13243 43131 13249
rect 43073 13240 43085 13243
rect 42024 13212 43085 13240
rect 42024 13200 42030 13212
rect 43073 13209 43085 13212
rect 43119 13209 43131 13243
rect 43073 13203 43131 13209
rect 56686 13200 56692 13252
rect 56744 13240 56750 13252
rect 57882 13240 57888 13252
rect 56744 13212 57888 13240
rect 56744 13200 56750 13212
rect 57882 13200 57888 13212
rect 57940 13240 57946 13252
rect 58360 13240 58388 13271
rect 60826 13268 60832 13280
rect 60884 13308 60890 13320
rect 61838 13308 61844 13320
rect 60884 13280 61844 13308
rect 60884 13268 60890 13280
rect 61838 13268 61844 13280
rect 61896 13268 61902 13320
rect 63402 13308 63408 13320
rect 63363 13280 63408 13308
rect 63402 13268 63408 13280
rect 63460 13268 63466 13320
rect 64598 13308 64604 13320
rect 64559 13280 64604 13308
rect 64598 13268 64604 13280
rect 64656 13268 64662 13320
rect 64874 13308 64880 13320
rect 64835 13280 64880 13308
rect 64874 13268 64880 13280
rect 64932 13268 64938 13320
rect 66622 13268 66628 13320
rect 66680 13308 66686 13320
rect 67177 13311 67235 13317
rect 67177 13308 67189 13311
rect 66680 13280 67189 13308
rect 66680 13268 66686 13280
rect 67177 13277 67189 13280
rect 67223 13277 67235 13311
rect 67450 13308 67456 13320
rect 67411 13280 67456 13308
rect 67177 13271 67235 13277
rect 67450 13268 67456 13280
rect 67508 13268 67514 13320
rect 70121 13311 70179 13317
rect 70121 13277 70133 13311
rect 70167 13308 70179 13311
rect 70210 13308 70216 13320
rect 70167 13280 70216 13308
rect 70167 13277 70179 13280
rect 70121 13271 70179 13277
rect 70210 13268 70216 13280
rect 70268 13268 70274 13320
rect 60274 13240 60280 13252
rect 57940 13212 58388 13240
rect 59280 13212 60280 13240
rect 57940 13200 57946 13212
rect 35894 13132 35900 13184
rect 35952 13172 35958 13184
rect 37645 13175 37703 13181
rect 37645 13172 37657 13175
rect 35952 13144 37657 13172
rect 35952 13132 35958 13144
rect 37645 13141 37657 13144
rect 37691 13141 37703 13175
rect 37645 13135 37703 13141
rect 44269 13175 44327 13181
rect 44269 13141 44281 13175
rect 44315 13172 44327 13175
rect 44450 13172 44456 13184
rect 44315 13144 44456 13172
rect 44315 13141 44327 13144
rect 44269 13135 44327 13141
rect 44450 13132 44456 13144
rect 44508 13132 44514 13184
rect 48590 13132 48596 13184
rect 48648 13172 48654 13184
rect 51445 13175 51503 13181
rect 51445 13172 51457 13175
rect 48648 13144 51457 13172
rect 48648 13132 48654 13144
rect 51445 13141 51457 13144
rect 51491 13141 51503 13175
rect 51445 13135 51503 13141
rect 54662 13132 54668 13184
rect 54720 13172 54726 13184
rect 54849 13175 54907 13181
rect 54849 13172 54861 13175
rect 54720 13144 54861 13172
rect 54720 13132 54726 13144
rect 54849 13141 54861 13144
rect 54895 13141 54907 13175
rect 54849 13135 54907 13141
rect 54938 13132 54944 13184
rect 54996 13172 55002 13184
rect 57149 13175 57207 13181
rect 57149 13172 57161 13175
rect 54996 13144 57161 13172
rect 54996 13132 55002 13144
rect 57149 13141 57161 13144
rect 57195 13141 57207 13175
rect 57149 13135 57207 13141
rect 57514 13132 57520 13184
rect 57572 13172 57578 13184
rect 58710 13172 58716 13184
rect 57572 13144 58716 13172
rect 57572 13132 57578 13144
rect 58710 13132 58716 13144
rect 58768 13172 58774 13184
rect 59280 13172 59308 13212
rect 60274 13200 60280 13212
rect 60332 13200 60338 13252
rect 69750 13240 69756 13252
rect 68664 13212 69756 13240
rect 58768 13144 59308 13172
rect 58768 13132 58774 13144
rect 60090 13132 60096 13184
rect 60148 13172 60154 13184
rect 62853 13175 62911 13181
rect 62853 13172 62865 13175
rect 60148 13144 62865 13172
rect 60148 13132 60154 13144
rect 62853 13141 62865 13144
rect 62899 13141 62911 13175
rect 62853 13135 62911 13141
rect 66165 13175 66223 13181
rect 66165 13141 66177 13175
rect 66211 13172 66223 13175
rect 67082 13172 67088 13184
rect 66211 13144 67088 13172
rect 66211 13141 66223 13144
rect 66165 13135 66223 13141
rect 67082 13132 67088 13144
rect 67140 13172 67146 13184
rect 68664 13172 68692 13212
rect 69750 13200 69756 13212
rect 69808 13200 69814 13252
rect 70366 13240 70394 13336
rect 71409 13311 71467 13317
rect 71409 13277 71421 13311
rect 71455 13308 71467 13311
rect 73890 13308 73896 13320
rect 71455 13280 73896 13308
rect 71455 13277 71467 13280
rect 71409 13271 71467 13277
rect 71424 13240 71452 13271
rect 73890 13268 73896 13280
rect 73948 13268 73954 13320
rect 70366 13212 71452 13240
rect 67140 13144 68692 13172
rect 68741 13175 68799 13181
rect 67140 13132 67146 13144
rect 68741 13141 68753 13175
rect 68787 13172 68799 13175
rect 70118 13172 70124 13184
rect 68787 13144 70124 13172
rect 68787 13141 68799 13144
rect 68741 13135 68799 13141
rect 70118 13132 70124 13144
rect 70176 13132 70182 13184
rect 70670 13132 70676 13184
rect 70728 13172 70734 13184
rect 70765 13175 70823 13181
rect 70765 13172 70777 13175
rect 70728 13144 70777 13172
rect 70728 13132 70734 13144
rect 70765 13141 70777 13144
rect 70811 13141 70823 13175
rect 70765 13135 70823 13141
rect 1104 13082 178848 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 34966 13082
rect 35018 13030 35030 13082
rect 35082 13030 35094 13082
rect 35146 13030 35158 13082
rect 35210 13030 65686 13082
rect 65738 13030 65750 13082
rect 65802 13030 65814 13082
rect 65866 13030 65878 13082
rect 65930 13030 96406 13082
rect 96458 13030 96470 13082
rect 96522 13030 96534 13082
rect 96586 13030 96598 13082
rect 96650 13030 127126 13082
rect 127178 13030 127190 13082
rect 127242 13030 127254 13082
rect 127306 13030 127318 13082
rect 127370 13030 157846 13082
rect 157898 13030 157910 13082
rect 157962 13030 157974 13082
rect 158026 13030 158038 13082
rect 158090 13030 178848 13082
rect 1104 13008 178848 13030
rect 32030 12968 32036 12980
rect 31991 12940 32036 12968
rect 32030 12928 32036 12940
rect 32088 12928 32094 12980
rect 34606 12968 34612 12980
rect 34567 12940 34612 12968
rect 34606 12928 34612 12940
rect 34664 12928 34670 12980
rect 36078 12928 36084 12980
rect 36136 12968 36142 12980
rect 36817 12971 36875 12977
rect 36817 12968 36829 12971
rect 36136 12940 36829 12968
rect 36136 12928 36142 12940
rect 36817 12937 36829 12940
rect 36863 12937 36875 12971
rect 36817 12931 36875 12937
rect 38746 12928 38752 12980
rect 38804 12968 38810 12980
rect 39206 12968 39212 12980
rect 38804 12940 39212 12968
rect 38804 12928 38810 12940
rect 39206 12928 39212 12940
rect 39264 12968 39270 12980
rect 39853 12971 39911 12977
rect 39853 12968 39865 12971
rect 39264 12940 39865 12968
rect 39264 12928 39270 12940
rect 39853 12937 39865 12940
rect 39899 12937 39911 12971
rect 39853 12931 39911 12937
rect 41506 12928 41512 12980
rect 41564 12968 41570 12980
rect 41969 12971 42027 12977
rect 41969 12968 41981 12971
rect 41564 12940 41981 12968
rect 41564 12928 41570 12940
rect 41969 12937 41981 12940
rect 42015 12968 42027 12971
rect 42610 12968 42616 12980
rect 42015 12940 42616 12968
rect 42015 12937 42027 12940
rect 41969 12931 42027 12937
rect 42610 12928 42616 12940
rect 42668 12928 42674 12980
rect 44634 12928 44640 12980
rect 44692 12968 44698 12980
rect 45646 12968 45652 12980
rect 44692 12940 45652 12968
rect 44692 12928 44698 12940
rect 45646 12928 45652 12940
rect 45704 12928 45710 12980
rect 56413 12971 56471 12977
rect 56413 12937 56425 12971
rect 56459 12968 56471 12971
rect 57146 12968 57152 12980
rect 56459 12940 57152 12968
rect 56459 12937 56471 12940
rect 56413 12931 56471 12937
rect 57146 12928 57152 12940
rect 57204 12928 57210 12980
rect 58526 12928 58532 12980
rect 58584 12968 58590 12980
rect 61657 12971 61715 12977
rect 61657 12968 61669 12971
rect 58584 12940 61669 12968
rect 58584 12928 58590 12940
rect 61657 12937 61669 12940
rect 61703 12937 61715 12971
rect 63954 12968 63960 12980
rect 61657 12931 61715 12937
rect 62040 12940 63960 12968
rect 30469 12835 30527 12841
rect 30469 12801 30481 12835
rect 30515 12832 30527 12835
rect 30834 12832 30840 12844
rect 30515 12804 30840 12832
rect 30515 12801 30527 12804
rect 30469 12795 30527 12801
rect 30834 12792 30840 12804
rect 30892 12832 30898 12844
rect 33045 12835 33103 12841
rect 33045 12832 33057 12835
rect 30892 12804 33057 12832
rect 30892 12792 30898 12804
rect 33045 12801 33057 12804
rect 33091 12832 33103 12835
rect 33502 12832 33508 12844
rect 33091 12804 33508 12832
rect 33091 12801 33103 12804
rect 33045 12795 33103 12801
rect 33502 12792 33508 12804
rect 33560 12832 33566 12844
rect 35437 12835 35495 12841
rect 35437 12832 35449 12835
rect 33560 12804 35449 12832
rect 33560 12792 33566 12804
rect 35437 12801 35449 12804
rect 35483 12832 35495 12835
rect 36170 12832 36176 12844
rect 35483 12804 36176 12832
rect 35483 12801 35495 12804
rect 35437 12795 35495 12801
rect 36170 12792 36176 12804
rect 36228 12832 36234 12844
rect 36998 12832 37004 12844
rect 36228 12804 37004 12832
rect 36228 12792 36234 12804
rect 36998 12792 37004 12804
rect 37056 12832 37062 12844
rect 38473 12835 38531 12841
rect 38473 12832 38485 12835
rect 37056 12804 38485 12832
rect 37056 12792 37062 12804
rect 38473 12801 38485 12804
rect 38519 12832 38531 12835
rect 40589 12835 40647 12841
rect 40589 12832 40601 12835
rect 38519 12804 40601 12832
rect 38519 12801 38531 12804
rect 38473 12795 38531 12801
rect 40589 12801 40601 12804
rect 40635 12832 40647 12835
rect 40954 12832 40960 12844
rect 40635 12804 40960 12832
rect 40635 12801 40647 12804
rect 40589 12795 40647 12801
rect 40954 12792 40960 12804
rect 41012 12832 41018 12844
rect 44269 12835 44327 12841
rect 44269 12832 44281 12835
rect 41012 12804 44281 12832
rect 41012 12792 41018 12804
rect 44269 12801 44281 12804
rect 44315 12832 44327 12835
rect 45462 12832 45468 12844
rect 44315 12804 45468 12832
rect 44315 12801 44327 12804
rect 44269 12795 44327 12801
rect 45462 12792 45468 12804
rect 45520 12792 45526 12844
rect 45830 12792 45836 12844
rect 45888 12832 45894 12844
rect 46845 12835 46903 12841
rect 46845 12832 46857 12835
rect 45888 12804 46857 12832
rect 45888 12792 45894 12804
rect 46845 12801 46857 12804
rect 46891 12801 46903 12835
rect 47026 12832 47032 12844
rect 46987 12804 47032 12832
rect 46845 12795 46903 12801
rect 47026 12792 47032 12804
rect 47084 12792 47090 12844
rect 47946 12792 47952 12844
rect 48004 12832 48010 12844
rect 49053 12835 49111 12841
rect 49053 12832 49065 12835
rect 48004 12804 49065 12832
rect 48004 12792 48010 12804
rect 49053 12801 49065 12804
rect 49099 12801 49111 12835
rect 54849 12835 54907 12841
rect 54849 12832 54861 12835
rect 49053 12795 49111 12801
rect 50908 12804 54861 12832
rect 30745 12767 30803 12773
rect 30745 12733 30757 12767
rect 30791 12764 30803 12767
rect 32950 12764 32956 12776
rect 30791 12736 32956 12764
rect 30791 12733 30803 12736
rect 30745 12727 30803 12733
rect 32950 12724 32956 12736
rect 33008 12724 33014 12776
rect 33318 12764 33324 12776
rect 33279 12736 33324 12764
rect 33318 12724 33324 12736
rect 33376 12724 33382 12776
rect 35713 12767 35771 12773
rect 35713 12733 35725 12767
rect 35759 12764 35771 12767
rect 37182 12764 37188 12776
rect 35759 12736 37188 12764
rect 35759 12733 35771 12736
rect 35713 12727 35771 12733
rect 37182 12724 37188 12736
rect 37240 12724 37246 12776
rect 38746 12764 38752 12776
rect 38707 12736 38752 12764
rect 38746 12724 38752 12736
rect 38804 12724 38810 12776
rect 40862 12764 40868 12776
rect 40823 12736 40868 12764
rect 40862 12724 40868 12736
rect 40920 12724 40926 12776
rect 44542 12764 44548 12776
rect 44503 12736 44548 12764
rect 44542 12724 44548 12736
rect 44600 12724 44606 12776
rect 46753 12767 46811 12773
rect 46753 12733 46765 12767
rect 46799 12764 46811 12767
rect 47118 12764 47124 12776
rect 46799 12736 47124 12764
rect 46799 12733 46811 12736
rect 46753 12727 46811 12733
rect 47118 12724 47124 12736
rect 47176 12764 47182 12776
rect 47578 12764 47584 12776
rect 47176 12736 47584 12764
rect 47176 12724 47182 12736
rect 47578 12724 47584 12736
rect 47636 12724 47642 12776
rect 48774 12764 48780 12776
rect 48735 12736 48780 12764
rect 48774 12724 48780 12736
rect 48832 12764 48838 12776
rect 50908 12773 50936 12804
rect 54849 12801 54861 12804
rect 54895 12832 54907 12835
rect 56686 12832 56692 12844
rect 54895 12804 56692 12832
rect 54895 12801 54907 12804
rect 54849 12795 54907 12801
rect 56686 12792 56692 12804
rect 56744 12792 56750 12844
rect 57054 12792 57060 12844
rect 57112 12832 57118 12844
rect 57425 12835 57483 12841
rect 57425 12832 57437 12835
rect 57112 12804 57437 12832
rect 57112 12792 57118 12804
rect 57425 12801 57437 12804
rect 57471 12801 57483 12835
rect 57606 12832 57612 12844
rect 57567 12804 57612 12832
rect 57425 12795 57483 12801
rect 57606 12792 57612 12804
rect 57664 12792 57670 12844
rect 57882 12792 57888 12844
rect 57940 12832 57946 12844
rect 59541 12835 59599 12841
rect 59541 12832 59553 12835
rect 57940 12804 59553 12832
rect 57940 12792 57946 12804
rect 59541 12801 59553 12804
rect 59587 12801 59599 12835
rect 59541 12795 59599 12801
rect 50893 12767 50951 12773
rect 50893 12764 50905 12767
rect 48832 12736 50905 12764
rect 48832 12724 48838 12736
rect 50893 12733 50905 12736
rect 50939 12733 50951 12767
rect 50893 12727 50951 12733
rect 50982 12724 50988 12776
rect 51040 12764 51046 12776
rect 51169 12767 51227 12773
rect 51169 12764 51181 12767
rect 51040 12736 51181 12764
rect 51040 12724 51046 12736
rect 51169 12733 51181 12736
rect 51215 12733 51227 12767
rect 55122 12764 55128 12776
rect 55083 12736 55128 12764
rect 51169 12727 51227 12733
rect 55122 12724 55128 12736
rect 55180 12724 55186 12776
rect 59814 12764 59820 12776
rect 59775 12736 59820 12764
rect 59814 12724 59820 12736
rect 59872 12724 59878 12776
rect 62040 12773 62068 12940
rect 63954 12928 63960 12940
rect 64012 12928 64018 12980
rect 67266 12928 67272 12980
rect 67324 12968 67330 12980
rect 69753 12971 69811 12977
rect 69753 12968 69765 12971
rect 67324 12940 69765 12968
rect 67324 12928 67330 12940
rect 69753 12937 69765 12940
rect 69799 12937 69811 12971
rect 69753 12931 69811 12937
rect 62301 12835 62359 12841
rect 62301 12801 62313 12835
rect 62347 12832 62359 12835
rect 63402 12832 63408 12844
rect 62347 12804 63408 12832
rect 62347 12801 62359 12804
rect 62301 12795 62359 12801
rect 63402 12792 63408 12804
rect 63460 12792 63466 12844
rect 66622 12832 66628 12844
rect 66583 12804 66628 12832
rect 66622 12792 66628 12804
rect 66680 12792 66686 12844
rect 68002 12792 68008 12844
rect 68060 12832 68066 12844
rect 68281 12835 68339 12841
rect 68281 12832 68293 12835
rect 68060 12804 68293 12832
rect 68060 12792 68066 12804
rect 68281 12801 68293 12804
rect 68327 12832 68339 12835
rect 69382 12832 69388 12844
rect 68327 12804 69388 12832
rect 68327 12801 68339 12804
rect 68281 12795 68339 12801
rect 69382 12792 69388 12804
rect 69440 12792 69446 12844
rect 70210 12792 70216 12844
rect 70268 12832 70274 12844
rect 70351 12835 70409 12841
rect 70351 12832 70363 12835
rect 70268 12804 70363 12832
rect 70268 12792 70274 12804
rect 70351 12801 70363 12804
rect 70397 12801 70409 12835
rect 70351 12795 70409 12801
rect 62025 12767 62083 12773
rect 62025 12733 62037 12767
rect 62071 12733 62083 12767
rect 62025 12727 62083 12733
rect 62117 12767 62175 12773
rect 62117 12733 62129 12767
rect 62163 12764 62175 12767
rect 63678 12764 63684 12776
rect 62163 12736 63684 12764
rect 62163 12733 62175 12736
rect 62117 12727 62175 12733
rect 63678 12724 63684 12736
rect 63736 12724 63742 12776
rect 64046 12724 64052 12776
rect 64104 12764 64110 12776
rect 64509 12767 64567 12773
rect 64509 12764 64521 12767
rect 64104 12736 64521 12764
rect 64104 12724 64110 12736
rect 64509 12733 64521 12736
rect 64555 12764 64567 12767
rect 64598 12764 64604 12776
rect 64555 12736 64604 12764
rect 64555 12733 64567 12736
rect 64509 12727 64567 12733
rect 64598 12724 64604 12736
rect 64656 12724 64662 12776
rect 64782 12764 64788 12776
rect 64743 12736 64788 12764
rect 64782 12724 64788 12736
rect 64840 12724 64846 12776
rect 65518 12724 65524 12776
rect 65576 12764 65582 12776
rect 66901 12767 66959 12773
rect 66901 12764 66913 12767
rect 65576 12736 66913 12764
rect 65576 12724 65582 12736
rect 66901 12733 66913 12736
rect 66947 12733 66959 12767
rect 70118 12764 70124 12776
rect 70079 12736 70124 12764
rect 66901 12727 66959 12733
rect 70118 12724 70124 12736
rect 70176 12764 70182 12776
rect 72970 12764 72976 12776
rect 70176 12736 72976 12764
rect 70176 12724 70182 12736
rect 72970 12724 72976 12736
rect 73028 12724 73034 12776
rect 50433 12699 50491 12705
rect 50433 12665 50445 12699
rect 50479 12696 50491 12699
rect 50614 12696 50620 12708
rect 50479 12668 50620 12696
rect 50479 12665 50491 12668
rect 50433 12659 50491 12665
rect 50614 12656 50620 12668
rect 50672 12656 50678 12708
rect 61197 12699 61255 12705
rect 61197 12665 61209 12699
rect 61243 12696 61255 12699
rect 62482 12696 62488 12708
rect 61243 12668 62488 12696
rect 61243 12665 61255 12668
rect 61197 12659 61255 12665
rect 62482 12656 62488 12668
rect 62540 12656 62546 12708
rect 63313 12699 63371 12705
rect 63313 12665 63325 12699
rect 63359 12696 63371 12699
rect 63494 12696 63500 12708
rect 63359 12668 63500 12696
rect 63359 12665 63371 12668
rect 63313 12659 63371 12665
rect 63494 12656 63500 12668
rect 63552 12656 63558 12708
rect 70026 12656 70032 12708
rect 70084 12696 70090 12708
rect 70213 12699 70271 12705
rect 70213 12696 70225 12699
rect 70084 12668 70225 12696
rect 70084 12656 70090 12668
rect 70213 12665 70225 12668
rect 70259 12665 70271 12699
rect 70213 12659 70271 12665
rect 46106 12588 46112 12640
rect 46164 12628 46170 12640
rect 46385 12631 46443 12637
rect 46385 12628 46397 12631
rect 46164 12600 46397 12628
rect 46164 12588 46170 12600
rect 46385 12597 46397 12600
rect 46431 12597 46443 12631
rect 52270 12628 52276 12640
rect 52231 12600 52276 12628
rect 46385 12591 46443 12597
rect 52270 12588 52276 12600
rect 52328 12588 52334 12640
rect 56962 12628 56968 12640
rect 56923 12600 56968 12628
rect 56962 12588 56968 12600
rect 57020 12588 57026 12640
rect 57333 12631 57391 12637
rect 57333 12597 57345 12631
rect 57379 12628 57391 12631
rect 58066 12628 58072 12640
rect 57379 12600 58072 12628
rect 57379 12597 57391 12600
rect 57333 12591 57391 12597
rect 58066 12588 58072 12600
rect 58124 12588 58130 12640
rect 61286 12588 61292 12640
rect 61344 12628 61350 12640
rect 62853 12631 62911 12637
rect 62853 12628 62865 12631
rect 61344 12600 62865 12628
rect 61344 12588 61350 12600
rect 62853 12597 62865 12600
rect 62899 12597 62911 12631
rect 62853 12591 62911 12597
rect 63221 12631 63279 12637
rect 63221 12597 63233 12631
rect 63267 12628 63279 12631
rect 65058 12628 65064 12640
rect 63267 12600 65064 12628
rect 63267 12597 63279 12600
rect 63221 12591 63279 12597
rect 65058 12588 65064 12600
rect 65116 12628 65122 12640
rect 66073 12631 66131 12637
rect 66073 12628 66085 12631
rect 65116 12600 66085 12628
rect 65116 12588 65122 12600
rect 66073 12597 66085 12600
rect 66119 12628 66131 12631
rect 68462 12628 68468 12640
rect 66119 12600 68468 12628
rect 66119 12597 66131 12600
rect 66073 12591 66131 12597
rect 68462 12588 68468 12600
rect 68520 12588 68526 12640
rect 1104 12538 178848 12560
rect 1104 12486 19606 12538
rect 19658 12486 19670 12538
rect 19722 12486 19734 12538
rect 19786 12486 19798 12538
rect 19850 12486 50326 12538
rect 50378 12486 50390 12538
rect 50442 12486 50454 12538
rect 50506 12486 50518 12538
rect 50570 12486 81046 12538
rect 81098 12486 81110 12538
rect 81162 12486 81174 12538
rect 81226 12486 81238 12538
rect 81290 12486 111766 12538
rect 111818 12486 111830 12538
rect 111882 12486 111894 12538
rect 111946 12486 111958 12538
rect 112010 12486 142486 12538
rect 142538 12486 142550 12538
rect 142602 12486 142614 12538
rect 142666 12486 142678 12538
rect 142730 12486 173206 12538
rect 173258 12486 173270 12538
rect 173322 12486 173334 12538
rect 173386 12486 173398 12538
rect 173450 12486 178848 12538
rect 1104 12464 178848 12486
rect 34790 12384 34796 12436
rect 34848 12424 34854 12436
rect 36173 12427 36231 12433
rect 36173 12424 36185 12427
rect 34848 12396 36185 12424
rect 34848 12384 34854 12396
rect 36173 12393 36185 12396
rect 36219 12393 36231 12427
rect 38381 12427 38439 12433
rect 38381 12424 38393 12427
rect 36173 12387 36231 12393
rect 36280 12396 38393 12424
rect 34514 12316 34520 12368
rect 34572 12356 34578 12368
rect 35434 12356 35440 12368
rect 34572 12328 35440 12356
rect 34572 12316 34578 12328
rect 35434 12316 35440 12328
rect 35492 12356 35498 12368
rect 36280 12356 36308 12396
rect 38381 12393 38393 12396
rect 38427 12393 38439 12427
rect 60366 12424 60372 12436
rect 60327 12396 60372 12424
rect 38381 12387 38439 12393
rect 60366 12384 60372 12396
rect 60424 12384 60430 12436
rect 60706 12396 70394 12424
rect 35492 12328 36308 12356
rect 35492 12316 35498 12328
rect 36078 12288 36084 12300
rect 36039 12260 36084 12288
rect 36078 12248 36084 12260
rect 36136 12248 36142 12300
rect 36998 12288 37004 12300
rect 36959 12260 37004 12288
rect 36998 12248 37004 12260
rect 37056 12248 37062 12300
rect 44910 12248 44916 12300
rect 44968 12288 44974 12300
rect 45462 12288 45468 12300
rect 44968 12260 45468 12288
rect 44968 12248 44974 12260
rect 45462 12248 45468 12260
rect 45520 12288 45526 12300
rect 46845 12291 46903 12297
rect 46845 12288 46857 12291
rect 45520 12260 46857 12288
rect 45520 12248 45526 12260
rect 46845 12257 46857 12260
rect 46891 12257 46903 12291
rect 56686 12288 56692 12300
rect 56647 12260 56692 12288
rect 46845 12251 46903 12257
rect 56686 12248 56692 12260
rect 56744 12248 56750 12300
rect 59081 12291 59139 12297
rect 59081 12257 59093 12291
rect 59127 12288 59139 12291
rect 60706 12288 60734 12396
rect 62942 12316 62948 12368
rect 63000 12356 63006 12368
rect 63000 12328 64184 12356
rect 63000 12316 63006 12328
rect 59127 12260 60734 12288
rect 59127 12257 59139 12260
rect 59081 12251 59139 12257
rect 36357 12223 36415 12229
rect 36357 12189 36369 12223
rect 36403 12220 36415 12223
rect 36538 12220 36544 12232
rect 36403 12192 36544 12220
rect 36403 12189 36415 12192
rect 36357 12183 36415 12189
rect 36538 12180 36544 12192
rect 36596 12180 36602 12232
rect 37277 12223 37335 12229
rect 37277 12189 37289 12223
rect 37323 12220 37335 12223
rect 42426 12220 42432 12232
rect 37323 12192 42432 12220
rect 37323 12189 37335 12192
rect 37277 12183 37335 12189
rect 42426 12180 42432 12192
rect 42484 12180 42490 12232
rect 47121 12223 47179 12229
rect 47121 12189 47133 12223
rect 47167 12220 47179 12223
rect 47210 12220 47216 12232
rect 47167 12192 47216 12220
rect 47167 12189 47179 12192
rect 47121 12183 47179 12189
rect 47210 12180 47216 12192
rect 47268 12180 47274 12232
rect 55766 12180 55772 12232
rect 55824 12220 55830 12232
rect 56965 12223 57023 12229
rect 56965 12220 56977 12223
rect 55824 12192 56977 12220
rect 55824 12180 55830 12192
rect 56965 12189 56977 12192
rect 57011 12189 57023 12223
rect 56965 12183 57023 12189
rect 61933 12223 61991 12229
rect 61933 12189 61945 12223
rect 61979 12189 61991 12223
rect 61933 12183 61991 12189
rect 36556 12152 36584 12180
rect 36998 12152 37004 12164
rect 36556 12124 37004 12152
rect 36998 12112 37004 12124
rect 37056 12112 37062 12164
rect 35526 12044 35532 12096
rect 35584 12084 35590 12096
rect 35713 12087 35771 12093
rect 35713 12084 35725 12087
rect 35584 12056 35725 12084
rect 35584 12044 35590 12056
rect 35713 12053 35725 12056
rect 35759 12053 35771 12087
rect 48406 12084 48412 12096
rect 48367 12056 48412 12084
rect 35713 12047 35771 12053
rect 48406 12044 48412 12056
rect 48464 12044 48470 12096
rect 58066 12084 58072 12096
rect 58027 12056 58072 12084
rect 58066 12044 58072 12056
rect 58124 12044 58130 12096
rect 61654 12044 61660 12096
rect 61712 12084 61718 12096
rect 61948 12084 61976 12183
rect 62114 12180 62120 12232
rect 62172 12220 62178 12232
rect 62209 12223 62267 12229
rect 62209 12220 62221 12223
rect 62172 12192 62221 12220
rect 62172 12180 62178 12192
rect 62209 12189 62221 12192
rect 62255 12189 62267 12223
rect 64046 12220 64052 12232
rect 64007 12192 64052 12220
rect 62209 12183 62267 12189
rect 64046 12180 64052 12192
rect 64104 12180 64110 12232
rect 64156 12220 64184 12328
rect 66070 12316 66076 12368
rect 66128 12356 66134 12368
rect 66128 12328 67404 12356
rect 66128 12316 66134 12328
rect 64325 12223 64383 12229
rect 64325 12220 64337 12223
rect 64156 12192 64337 12220
rect 64325 12189 64337 12192
rect 64371 12189 64383 12223
rect 64325 12183 64383 12189
rect 66622 12180 66628 12232
rect 66680 12220 66686 12232
rect 67269 12223 67327 12229
rect 67269 12220 67281 12223
rect 66680 12192 67281 12220
rect 66680 12180 66686 12192
rect 64064 12152 64092 12180
rect 62868 12124 64092 12152
rect 62868 12084 62896 12124
rect 67192 12096 67220 12192
rect 67269 12189 67281 12192
rect 67315 12189 67327 12223
rect 67376 12220 67404 12328
rect 70366 12288 70394 12396
rect 93946 12288 93952 12300
rect 70366 12260 93952 12288
rect 93946 12248 93952 12260
rect 94004 12248 94010 12300
rect 67545 12223 67603 12229
rect 67545 12220 67557 12223
rect 67376 12192 67557 12220
rect 67269 12183 67327 12189
rect 67545 12189 67557 12192
rect 67591 12189 67603 12223
rect 69385 12223 69443 12229
rect 69385 12220 69397 12223
rect 67545 12183 67603 12189
rect 68204 12192 69397 12220
rect 61712 12056 62896 12084
rect 63497 12087 63555 12093
rect 61712 12044 61718 12056
rect 63497 12053 63509 12087
rect 63543 12084 63555 12087
rect 63862 12084 63868 12096
rect 63543 12056 63868 12084
rect 63543 12053 63555 12056
rect 63497 12047 63555 12053
rect 63862 12044 63868 12056
rect 63920 12044 63926 12096
rect 65150 12044 65156 12096
rect 65208 12084 65214 12096
rect 65334 12084 65340 12096
rect 65208 12056 65340 12084
rect 65208 12044 65214 12056
rect 65334 12044 65340 12056
rect 65392 12084 65398 12096
rect 65429 12087 65487 12093
rect 65429 12084 65441 12087
rect 65392 12056 65441 12084
rect 65392 12044 65398 12056
rect 65429 12053 65441 12056
rect 65475 12053 65487 12087
rect 67174 12084 67180 12096
rect 67087 12056 67180 12084
rect 65429 12047 65487 12053
rect 67174 12044 67180 12056
rect 67232 12084 67238 12096
rect 68204 12084 68232 12192
rect 69385 12189 69397 12192
rect 69431 12189 69443 12223
rect 69658 12220 69664 12232
rect 69619 12192 69664 12220
rect 69385 12183 69443 12189
rect 69658 12180 69664 12192
rect 69716 12180 69722 12232
rect 68646 12084 68652 12096
rect 67232 12056 68232 12084
rect 68607 12056 68652 12084
rect 67232 12044 67238 12056
rect 68646 12044 68652 12056
rect 68704 12044 68710 12096
rect 69842 12044 69848 12096
rect 69900 12084 69906 12096
rect 70946 12084 70952 12096
rect 69900 12056 70952 12084
rect 69900 12044 69906 12056
rect 70946 12044 70952 12056
rect 71004 12044 71010 12096
rect 1104 11994 178848 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 34966 11994
rect 35018 11942 35030 11994
rect 35082 11942 35094 11994
rect 35146 11942 35158 11994
rect 35210 11942 65686 11994
rect 65738 11942 65750 11994
rect 65802 11942 65814 11994
rect 65866 11942 65878 11994
rect 65930 11942 96406 11994
rect 96458 11942 96470 11994
rect 96522 11942 96534 11994
rect 96586 11942 96598 11994
rect 96650 11942 127126 11994
rect 127178 11942 127190 11994
rect 127242 11942 127254 11994
rect 127306 11942 127318 11994
rect 127370 11942 157846 11994
rect 157898 11942 157910 11994
rect 157962 11942 157974 11994
rect 158026 11942 158038 11994
rect 158090 11942 178848 11994
rect 1104 11920 178848 11942
rect 61654 11880 61660 11892
rect 61615 11852 61660 11880
rect 61654 11840 61660 11852
rect 61712 11840 61718 11892
rect 57882 11704 57888 11756
rect 57940 11744 57946 11756
rect 59265 11747 59323 11753
rect 59265 11744 59277 11747
rect 57940 11716 59277 11744
rect 57940 11704 57946 11716
rect 59265 11713 59277 11716
rect 59311 11713 59323 11747
rect 59265 11707 59323 11713
rect 63586 11704 63592 11756
rect 63644 11744 63650 11756
rect 65337 11747 65395 11753
rect 65337 11744 65349 11747
rect 63644 11716 65349 11744
rect 63644 11704 63650 11716
rect 65337 11713 65349 11716
rect 65383 11713 65395 11747
rect 65337 11707 65395 11713
rect 65978 11704 65984 11756
rect 66036 11744 66042 11756
rect 67453 11747 67511 11753
rect 67453 11744 67465 11747
rect 66036 11716 67465 11744
rect 66036 11704 66042 11716
rect 67453 11713 67465 11716
rect 67499 11713 67511 11747
rect 67453 11707 67511 11713
rect 59538 11676 59544 11688
rect 59499 11648 59544 11676
rect 59538 11636 59544 11648
rect 59596 11636 59602 11688
rect 60366 11636 60372 11688
rect 60424 11676 60430 11688
rect 61841 11679 61899 11685
rect 61841 11676 61853 11679
rect 60424 11648 61853 11676
rect 60424 11636 60430 11648
rect 61841 11645 61853 11648
rect 61887 11645 61899 11679
rect 61841 11639 61899 11645
rect 64046 11636 64052 11688
rect 64104 11676 64110 11688
rect 65061 11679 65119 11685
rect 65061 11676 65073 11679
rect 64104 11648 65073 11676
rect 64104 11636 64110 11648
rect 65061 11645 65073 11648
rect 65107 11676 65119 11679
rect 67174 11676 67180 11688
rect 65107 11648 67180 11676
rect 65107 11645 65119 11648
rect 65061 11639 65119 11645
rect 67174 11636 67180 11648
rect 67232 11636 67238 11688
rect 60274 11500 60280 11552
rect 60332 11540 60338 11552
rect 60550 11540 60556 11552
rect 60332 11512 60556 11540
rect 60332 11500 60338 11512
rect 60550 11500 60556 11512
rect 60608 11540 60614 11552
rect 60829 11543 60887 11549
rect 60829 11540 60841 11543
rect 60608 11512 60841 11540
rect 60608 11500 60614 11512
rect 60829 11509 60841 11512
rect 60875 11509 60887 11543
rect 60829 11503 60887 11509
rect 66254 11500 66260 11552
rect 66312 11540 66318 11552
rect 66441 11543 66499 11549
rect 66441 11540 66453 11543
rect 66312 11512 66453 11540
rect 66312 11500 66318 11512
rect 66441 11509 66453 11512
rect 66487 11509 66499 11543
rect 68554 11540 68560 11552
rect 68515 11512 68560 11540
rect 66441 11503 66499 11509
rect 68554 11500 68560 11512
rect 68612 11500 68618 11552
rect 1104 11450 178848 11472
rect 1104 11398 19606 11450
rect 19658 11398 19670 11450
rect 19722 11398 19734 11450
rect 19786 11398 19798 11450
rect 19850 11398 50326 11450
rect 50378 11398 50390 11450
rect 50442 11398 50454 11450
rect 50506 11398 50518 11450
rect 50570 11398 81046 11450
rect 81098 11398 81110 11450
rect 81162 11398 81174 11450
rect 81226 11398 81238 11450
rect 81290 11398 111766 11450
rect 111818 11398 111830 11450
rect 111882 11398 111894 11450
rect 111946 11398 111958 11450
rect 112010 11398 142486 11450
rect 142538 11398 142550 11450
rect 142602 11398 142614 11450
rect 142666 11398 142678 11450
rect 142730 11398 173206 11450
rect 173258 11398 173270 11450
rect 173322 11398 173334 11450
rect 173386 11398 173398 11450
rect 173450 11398 178848 11450
rect 1104 11376 178848 11398
rect 68925 11339 68983 11345
rect 68925 11305 68937 11339
rect 68971 11336 68983 11339
rect 70394 11336 70400 11348
rect 68971 11308 70400 11336
rect 68971 11305 68983 11308
rect 68925 11299 68983 11305
rect 70394 11296 70400 11308
rect 70452 11336 70458 11348
rect 71130 11336 71136 11348
rect 70452 11308 71136 11336
rect 70452 11296 70458 11308
rect 71130 11296 71136 11308
rect 71188 11296 71194 11348
rect 67174 11160 67180 11212
rect 67232 11200 67238 11212
rect 67361 11203 67419 11209
rect 67361 11200 67373 11203
rect 67232 11172 67373 11200
rect 67232 11160 67238 11172
rect 67361 11169 67373 11172
rect 67407 11169 67419 11203
rect 67361 11163 67419 11169
rect 67542 11092 67548 11144
rect 67600 11132 67606 11144
rect 67637 11135 67695 11141
rect 67637 11132 67649 11135
rect 67600 11104 67649 11132
rect 67600 11092 67606 11104
rect 67637 11101 67649 11104
rect 67683 11101 67695 11135
rect 67637 11095 67695 11101
rect 1104 10906 178848 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 34966 10906
rect 35018 10854 35030 10906
rect 35082 10854 35094 10906
rect 35146 10854 35158 10906
rect 35210 10854 65686 10906
rect 65738 10854 65750 10906
rect 65802 10854 65814 10906
rect 65866 10854 65878 10906
rect 65930 10854 96406 10906
rect 96458 10854 96470 10906
rect 96522 10854 96534 10906
rect 96586 10854 96598 10906
rect 96650 10854 127126 10906
rect 127178 10854 127190 10906
rect 127242 10854 127254 10906
rect 127306 10854 127318 10906
rect 127370 10854 157846 10906
rect 157898 10854 157910 10906
rect 157962 10854 157974 10906
rect 158026 10854 158038 10906
rect 158090 10854 178848 10906
rect 1104 10832 178848 10854
rect 33226 10752 33232 10804
rect 33284 10792 33290 10804
rect 33413 10795 33471 10801
rect 33413 10792 33425 10795
rect 33284 10764 33425 10792
rect 33284 10752 33290 10764
rect 33413 10761 33425 10764
rect 33459 10761 33471 10795
rect 33413 10755 33471 10761
rect 33778 10752 33784 10804
rect 33836 10792 33842 10804
rect 34517 10795 34575 10801
rect 34517 10792 34529 10795
rect 33836 10764 34529 10792
rect 33836 10752 33842 10764
rect 34517 10761 34529 10764
rect 34563 10761 34575 10795
rect 34517 10755 34575 10761
rect 33229 10591 33287 10597
rect 33229 10557 33241 10591
rect 33275 10588 33287 10591
rect 33594 10588 33600 10600
rect 33275 10560 33600 10588
rect 33275 10557 33287 10560
rect 33229 10551 33287 10557
rect 33594 10548 33600 10560
rect 33652 10588 33658 10600
rect 34238 10588 34244 10600
rect 33652 10560 34244 10588
rect 33652 10548 33658 10560
rect 34238 10548 34244 10560
rect 34296 10588 34302 10600
rect 34333 10591 34391 10597
rect 34333 10588 34345 10591
rect 34296 10560 34345 10588
rect 34296 10548 34302 10560
rect 34333 10557 34345 10560
rect 34379 10557 34391 10591
rect 60366 10588 60372 10600
rect 60327 10560 60372 10588
rect 34333 10551 34391 10557
rect 60366 10548 60372 10560
rect 60424 10548 60430 10600
rect 60645 10591 60703 10597
rect 60645 10557 60657 10591
rect 60691 10588 60703 10591
rect 65426 10588 65432 10600
rect 60691 10560 65432 10588
rect 60691 10557 60703 10560
rect 60645 10551 60703 10557
rect 65426 10548 65432 10560
rect 65484 10548 65490 10600
rect 33045 10523 33103 10529
rect 33045 10489 33057 10523
rect 33091 10520 33103 10523
rect 33778 10520 33784 10532
rect 33091 10492 33784 10520
rect 33091 10489 33103 10492
rect 33045 10483 33103 10489
rect 33778 10480 33784 10492
rect 33836 10480 33842 10532
rect 34149 10523 34207 10529
rect 34149 10489 34161 10523
rect 34195 10520 34207 10523
rect 35802 10520 35808 10532
rect 34195 10492 35808 10520
rect 34195 10489 34207 10492
rect 34149 10483 34207 10489
rect 35802 10480 35808 10492
rect 35860 10480 35866 10532
rect 1104 10362 178848 10384
rect 1104 10310 19606 10362
rect 19658 10310 19670 10362
rect 19722 10310 19734 10362
rect 19786 10310 19798 10362
rect 19850 10310 50326 10362
rect 50378 10310 50390 10362
rect 50442 10310 50454 10362
rect 50506 10310 50518 10362
rect 50570 10310 81046 10362
rect 81098 10310 81110 10362
rect 81162 10310 81174 10362
rect 81226 10310 81238 10362
rect 81290 10310 111766 10362
rect 111818 10310 111830 10362
rect 111882 10310 111894 10362
rect 111946 10310 111958 10362
rect 112010 10310 142486 10362
rect 142538 10310 142550 10362
rect 142602 10310 142614 10362
rect 142666 10310 142678 10362
rect 142730 10310 173206 10362
rect 173258 10310 173270 10362
rect 173322 10310 173334 10362
rect 173386 10310 173398 10362
rect 173450 10310 178848 10362
rect 1104 10288 178848 10310
rect 32674 10248 32680 10260
rect 31404 10220 32680 10248
rect 31404 10189 31432 10220
rect 32674 10208 32680 10220
rect 32732 10208 32738 10260
rect 33594 10248 33600 10260
rect 32784 10220 33600 10248
rect 31389 10183 31447 10189
rect 31389 10149 31401 10183
rect 31435 10149 31447 10183
rect 31389 10143 31447 10149
rect 31662 10140 31668 10192
rect 31720 10180 31726 10192
rect 31757 10183 31815 10189
rect 31757 10180 31769 10183
rect 31720 10152 31769 10180
rect 31720 10140 31726 10152
rect 31757 10149 31769 10152
rect 31803 10149 31815 10183
rect 32784 10180 32812 10220
rect 33594 10208 33600 10220
rect 33652 10208 33658 10260
rect 32950 10180 32956 10192
rect 31757 10143 31815 10149
rect 32508 10152 32812 10180
rect 32911 10152 32956 10180
rect 31573 10115 31631 10121
rect 31573 10081 31585 10115
rect 31619 10112 31631 10115
rect 32508 10112 32536 10152
rect 32784 10121 32812 10152
rect 32950 10140 32956 10152
rect 33008 10140 33014 10192
rect 33318 10140 33324 10192
rect 33376 10180 33382 10192
rect 33781 10183 33839 10189
rect 33781 10180 33793 10183
rect 33376 10152 33793 10180
rect 33376 10140 33382 10152
rect 33781 10149 33793 10152
rect 33827 10149 33839 10183
rect 33781 10143 33839 10149
rect 38746 10140 38752 10192
rect 38804 10180 38810 10192
rect 39945 10183 40003 10189
rect 39945 10180 39957 10183
rect 38804 10152 39957 10180
rect 38804 10140 38810 10152
rect 39945 10149 39957 10152
rect 39991 10149 40003 10183
rect 41598 10180 41604 10192
rect 39945 10143 40003 10149
rect 40052 10152 41460 10180
rect 41559 10152 41604 10180
rect 31619 10084 32536 10112
rect 32585 10115 32643 10121
rect 31619 10081 31631 10084
rect 31573 10075 31631 10081
rect 32585 10081 32597 10115
rect 32631 10081 32643 10115
rect 32585 10075 32643 10081
rect 32769 10115 32827 10121
rect 32769 10081 32781 10115
rect 32815 10081 32827 10115
rect 32769 10075 32827 10081
rect 33413 10115 33471 10121
rect 33413 10081 33425 10115
rect 33459 10081 33471 10115
rect 33594 10112 33600 10124
rect 33555 10084 33600 10112
rect 33413 10075 33471 10081
rect 32600 9976 32628 10075
rect 33428 10044 33456 10075
rect 33594 10072 33600 10084
rect 33652 10072 33658 10124
rect 39577 10115 39635 10121
rect 39577 10081 39589 10115
rect 39623 10081 39635 10115
rect 39758 10112 39764 10124
rect 39719 10084 39764 10112
rect 39577 10075 39635 10081
rect 34698 10044 34704 10056
rect 33428 10016 34704 10044
rect 34698 10004 34704 10016
rect 34756 10004 34762 10056
rect 39592 10044 39620 10075
rect 39758 10072 39764 10084
rect 39816 10112 39822 10124
rect 40052 10112 40080 10152
rect 41432 10121 41460 10152
rect 41598 10140 41604 10152
rect 41656 10140 41662 10192
rect 44542 10140 44548 10192
rect 44600 10180 44606 10192
rect 45281 10183 45339 10189
rect 45281 10180 45293 10183
rect 44600 10152 45293 10180
rect 44600 10140 44606 10152
rect 45281 10149 45293 10152
rect 45327 10149 45339 10183
rect 45281 10143 45339 10149
rect 46474 10140 46480 10192
rect 46532 10180 46538 10192
rect 46569 10183 46627 10189
rect 46569 10180 46581 10183
rect 46532 10152 46581 10180
rect 46532 10140 46538 10152
rect 46569 10149 46581 10152
rect 46615 10149 46627 10183
rect 47946 10180 47952 10192
rect 47907 10152 47952 10180
rect 46569 10143 46627 10149
rect 47946 10140 47952 10152
rect 48004 10140 48010 10192
rect 60366 10180 60372 10192
rect 58728 10152 60372 10180
rect 39816 10084 40080 10112
rect 41233 10115 41291 10121
rect 39816 10072 39822 10084
rect 41233 10081 41245 10115
rect 41279 10081 41291 10115
rect 41233 10075 41291 10081
rect 41417 10115 41475 10121
rect 41417 10081 41429 10115
rect 41463 10081 41475 10115
rect 41417 10075 41475 10081
rect 44913 10115 44971 10121
rect 44913 10081 44925 10115
rect 44959 10081 44971 10115
rect 44913 10075 44971 10081
rect 45097 10115 45155 10121
rect 45097 10081 45109 10115
rect 45143 10081 45155 10115
rect 46198 10112 46204 10124
rect 46159 10084 46204 10112
rect 45097 10075 45155 10081
rect 40770 10044 40776 10056
rect 39592 10016 40776 10044
rect 40770 10004 40776 10016
rect 40828 10004 40834 10056
rect 41248 10044 41276 10075
rect 42518 10044 42524 10056
rect 41248 10016 42524 10044
rect 42518 10004 42524 10016
rect 42576 10004 42582 10056
rect 34422 9976 34428 9988
rect 32600 9948 34428 9976
rect 34422 9936 34428 9948
rect 34480 9936 34486 9988
rect 44928 9976 44956 10075
rect 45112 10044 45140 10075
rect 46198 10072 46204 10084
rect 46256 10072 46262 10124
rect 46385 10115 46443 10121
rect 46385 10081 46397 10115
rect 46431 10081 46443 10115
rect 46385 10075 46443 10081
rect 46400 10044 46428 10075
rect 47026 10072 47032 10124
rect 47084 10112 47090 10124
rect 47581 10115 47639 10121
rect 47581 10112 47593 10115
rect 47084 10084 47593 10112
rect 47084 10072 47090 10084
rect 47581 10081 47593 10084
rect 47627 10081 47639 10115
rect 47762 10112 47768 10124
rect 47723 10084 47768 10112
rect 47581 10075 47639 10081
rect 47762 10072 47768 10084
rect 47820 10072 47826 10124
rect 56502 10072 56508 10124
rect 56560 10112 56566 10124
rect 58728 10121 58756 10152
rect 60366 10140 60372 10152
rect 60424 10180 60430 10192
rect 62761 10183 62819 10189
rect 60424 10152 62620 10180
rect 60424 10140 60430 10152
rect 62592 10121 62620 10152
rect 62761 10149 62773 10183
rect 62807 10180 62819 10183
rect 64874 10180 64880 10192
rect 62807 10152 64880 10180
rect 62807 10149 62819 10152
rect 62761 10143 62819 10149
rect 64874 10140 64880 10152
rect 64932 10140 64938 10192
rect 66257 10183 66315 10189
rect 66257 10149 66269 10183
rect 66303 10180 66315 10183
rect 67542 10180 67548 10192
rect 66303 10152 67548 10180
rect 66303 10149 66315 10152
rect 66257 10143 66315 10149
rect 67542 10140 67548 10152
rect 67600 10140 67606 10192
rect 56689 10115 56747 10121
rect 56689 10112 56701 10115
rect 56560 10084 56701 10112
rect 56560 10072 56566 10084
rect 56689 10081 56701 10084
rect 56735 10112 56747 10115
rect 58713 10115 58771 10121
rect 58713 10112 58725 10115
rect 56735 10084 58725 10112
rect 56735 10081 56747 10084
rect 56689 10075 56747 10081
rect 58713 10081 58725 10084
rect 58759 10081 58771 10115
rect 58713 10075 58771 10081
rect 62393 10115 62451 10121
rect 62393 10081 62405 10115
rect 62439 10081 62451 10115
rect 62393 10075 62451 10081
rect 62577 10115 62635 10121
rect 62577 10081 62589 10115
rect 62623 10081 62635 10115
rect 62577 10075 62635 10081
rect 46934 10044 46940 10056
rect 45112 10016 46940 10044
rect 46934 10004 46940 10016
rect 46992 10044 46998 10056
rect 47780 10044 47808 10072
rect 46992 10016 47808 10044
rect 62408 10044 62436 10075
rect 63678 10072 63684 10124
rect 63736 10112 63742 10124
rect 65889 10115 65947 10121
rect 65889 10112 65901 10115
rect 63736 10084 65901 10112
rect 63736 10072 63742 10084
rect 65889 10081 65901 10084
rect 65935 10081 65947 10115
rect 65889 10075 65947 10081
rect 66073 10115 66131 10121
rect 66073 10081 66085 10115
rect 66119 10081 66131 10115
rect 66073 10075 66131 10081
rect 64598 10044 64604 10056
rect 62408 10016 64604 10044
rect 46992 10004 46998 10016
rect 64598 10004 64604 10016
rect 64656 10004 64662 10056
rect 65426 10004 65432 10056
rect 65484 10044 65490 10056
rect 66088 10044 66116 10075
rect 65484 10016 66116 10044
rect 65484 10004 65490 10016
rect 45278 9976 45284 9988
rect 44928 9948 45284 9976
rect 45278 9936 45284 9948
rect 45336 9936 45342 9988
rect 58897 9979 58955 9985
rect 58897 9945 58909 9979
rect 58943 9976 58955 9979
rect 60090 9976 60096 9988
rect 58943 9948 60096 9976
rect 58943 9945 58955 9948
rect 58897 9939 58955 9945
rect 60090 9936 60096 9948
rect 60148 9936 60154 9988
rect 56870 9908 56876 9920
rect 56831 9880 56876 9908
rect 56870 9868 56876 9880
rect 56928 9868 56934 9920
rect 1104 9818 178848 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 34966 9818
rect 35018 9766 35030 9818
rect 35082 9766 35094 9818
rect 35146 9766 35158 9818
rect 35210 9766 65686 9818
rect 65738 9766 65750 9818
rect 65802 9766 65814 9818
rect 65866 9766 65878 9818
rect 65930 9766 96406 9818
rect 96458 9766 96470 9818
rect 96522 9766 96534 9818
rect 96586 9766 96598 9818
rect 96650 9766 127126 9818
rect 127178 9766 127190 9818
rect 127242 9766 127254 9818
rect 127306 9766 127318 9818
rect 127370 9766 157846 9818
rect 157898 9766 157910 9818
rect 157962 9766 157974 9818
rect 158026 9766 158038 9818
rect 158090 9766 178848 9818
rect 1104 9744 178848 9766
rect 37182 9596 37188 9648
rect 37240 9636 37246 9648
rect 37369 9639 37427 9645
rect 37369 9636 37381 9639
rect 37240 9608 37381 9636
rect 37240 9596 37246 9608
rect 37369 9605 37381 9608
rect 37415 9605 37427 9639
rect 37369 9599 37427 9605
rect 38562 9596 38568 9648
rect 38620 9636 38626 9648
rect 38657 9639 38715 9645
rect 38657 9636 38669 9639
rect 38620 9608 38669 9636
rect 38620 9596 38626 9608
rect 38657 9605 38669 9608
rect 38703 9605 38715 9639
rect 40862 9636 40868 9648
rect 40823 9608 40868 9636
rect 38657 9599 38715 9605
rect 40862 9596 40868 9608
rect 40920 9596 40926 9648
rect 42426 9636 42432 9648
rect 42387 9608 42432 9636
rect 42426 9596 42432 9608
rect 42484 9596 42490 9648
rect 47210 9636 47216 9648
rect 47171 9608 47216 9636
rect 47210 9596 47216 9608
rect 47268 9596 47274 9648
rect 49145 9639 49203 9645
rect 49145 9605 49157 9639
rect 49191 9636 49203 9639
rect 50982 9636 50988 9648
rect 49191 9608 50988 9636
rect 49191 9605 49203 9608
rect 49145 9599 49203 9605
rect 50982 9596 50988 9608
rect 51040 9596 51046 9648
rect 55122 9596 55128 9648
rect 55180 9636 55186 9648
rect 55217 9639 55275 9645
rect 55217 9636 55229 9639
rect 55180 9608 55229 9636
rect 55180 9596 55186 9608
rect 55217 9605 55229 9608
rect 55263 9605 55275 9639
rect 55217 9599 55275 9605
rect 57425 9639 57483 9645
rect 57425 9605 57437 9639
rect 57471 9636 57483 9639
rect 57974 9636 57980 9648
rect 57471 9608 57980 9636
rect 57471 9605 57483 9608
rect 57425 9599 57483 9605
rect 57974 9596 57980 9608
rect 58032 9596 58038 9648
rect 58345 9639 58403 9645
rect 58345 9605 58357 9639
rect 58391 9636 58403 9639
rect 59814 9636 59820 9648
rect 58391 9608 59820 9636
rect 58391 9605 58403 9608
rect 58345 9599 58403 9605
rect 59814 9596 59820 9608
rect 59872 9596 59878 9648
rect 72510 9636 72516 9648
rect 60706 9608 72516 9636
rect 42260 9540 49096 9568
rect 29086 9460 29092 9512
rect 29144 9500 29150 9512
rect 32030 9500 32036 9512
rect 29144 9472 32036 9500
rect 29144 9460 29150 9472
rect 32030 9460 32036 9472
rect 32088 9500 32094 9512
rect 36262 9500 36268 9512
rect 32088 9472 36268 9500
rect 32088 9460 32094 9472
rect 36262 9460 36268 9472
rect 36320 9460 36326 9512
rect 37185 9503 37243 9509
rect 37185 9469 37197 9503
rect 37231 9500 37243 9503
rect 38473 9503 38531 9509
rect 38473 9500 38485 9503
rect 37231 9472 38485 9500
rect 37231 9469 37243 9472
rect 37185 9463 37243 9469
rect 38473 9469 38485 9472
rect 38519 9500 38531 9503
rect 39758 9500 39764 9512
rect 38519 9472 39764 9500
rect 38519 9469 38531 9472
rect 38473 9463 38531 9469
rect 39758 9460 39764 9472
rect 39816 9500 39822 9512
rect 42260 9509 42288 9540
rect 40681 9503 40739 9509
rect 40681 9500 40693 9503
rect 39816 9472 40693 9500
rect 39816 9460 39822 9472
rect 40681 9469 40693 9472
rect 40727 9469 40739 9503
rect 40681 9463 40739 9469
rect 42245 9503 42303 9509
rect 42245 9469 42257 9503
rect 42291 9469 42303 9503
rect 42245 9463 42303 9469
rect 47029 9503 47087 9509
rect 47029 9469 47041 9503
rect 47075 9500 47087 9503
rect 47762 9500 47768 9512
rect 47075 9472 47768 9500
rect 47075 9469 47087 9472
rect 47029 9463 47087 9469
rect 47762 9460 47768 9472
rect 47820 9500 47826 9512
rect 48961 9503 49019 9509
rect 48961 9500 48973 9503
rect 47820 9472 48973 9500
rect 47820 9460 47826 9472
rect 48961 9469 48973 9472
rect 49007 9469 49019 9503
rect 49068 9500 49096 9540
rect 49694 9528 49700 9580
rect 49752 9568 49758 9580
rect 50614 9568 50620 9580
rect 49752 9540 50620 9568
rect 49752 9528 49758 9540
rect 50614 9528 50620 9540
rect 50672 9568 50678 9580
rect 54478 9568 54484 9580
rect 50672 9540 54484 9568
rect 50672 9528 50678 9540
rect 54478 9528 54484 9540
rect 54536 9528 54542 9580
rect 55398 9568 55404 9580
rect 54956 9540 55404 9568
rect 54956 9500 54984 9540
rect 55398 9528 55404 9540
rect 55456 9568 55462 9580
rect 56502 9568 56508 9580
rect 55456 9540 56508 9568
rect 55456 9528 55462 9540
rect 56502 9528 56508 9540
rect 56560 9528 56566 9580
rect 56597 9571 56655 9577
rect 56597 9537 56609 9571
rect 56643 9568 56655 9571
rect 59538 9568 59544 9580
rect 56643 9540 59544 9568
rect 56643 9537 56655 9540
rect 56597 9531 56655 9537
rect 59538 9528 59544 9540
rect 59596 9528 59602 9580
rect 60706 9568 60734 9608
rect 72510 9596 72516 9608
rect 72568 9596 72574 9648
rect 63586 9568 63592 9580
rect 59648 9540 60734 9568
rect 63547 9540 63592 9568
rect 49068 9472 54984 9500
rect 55033 9503 55091 9509
rect 48961 9463 49019 9469
rect 55033 9469 55045 9503
rect 55079 9500 55091 9503
rect 56413 9503 56471 9509
rect 56413 9500 56425 9503
rect 55079 9472 56425 9500
rect 55079 9469 55091 9472
rect 55033 9463 55091 9469
rect 56413 9469 56425 9472
rect 56459 9500 56471 9503
rect 56870 9500 56876 9512
rect 56459 9472 56876 9500
rect 56459 9469 56471 9472
rect 56413 9463 56471 9469
rect 56870 9460 56876 9472
rect 56928 9500 56934 9512
rect 57241 9503 57299 9509
rect 57241 9500 57253 9503
rect 56928 9472 57253 9500
rect 56928 9460 56934 9472
rect 57241 9469 57253 9472
rect 57287 9500 57299 9503
rect 58161 9503 58219 9509
rect 58161 9500 58173 9503
rect 57287 9472 58173 9500
rect 57287 9469 57299 9472
rect 57241 9463 57299 9469
rect 58161 9469 58173 9472
rect 58207 9469 58219 9503
rect 58161 9463 58219 9469
rect 30190 9392 30196 9444
rect 30248 9432 30254 9444
rect 36078 9432 36084 9444
rect 30248 9404 36084 9432
rect 30248 9392 30254 9404
rect 36078 9392 36084 9404
rect 36136 9392 36142 9444
rect 37001 9435 37059 9441
rect 37001 9401 37013 9435
rect 37047 9432 37059 9435
rect 37366 9432 37372 9444
rect 37047 9404 37372 9432
rect 37047 9401 37059 9404
rect 37001 9395 37059 9401
rect 37366 9392 37372 9404
rect 37424 9392 37430 9444
rect 38289 9435 38347 9441
rect 38289 9401 38301 9435
rect 38335 9432 38347 9435
rect 38378 9432 38384 9444
rect 38335 9404 38384 9432
rect 38335 9401 38347 9404
rect 38289 9395 38347 9401
rect 38378 9392 38384 9404
rect 38436 9392 38442 9444
rect 40497 9435 40555 9441
rect 40497 9401 40509 9435
rect 40543 9401 40555 9435
rect 40497 9395 40555 9401
rect 36096 9364 36124 9392
rect 37734 9364 37740 9376
rect 36096 9336 37740 9364
rect 37734 9324 37740 9336
rect 37792 9324 37798 9376
rect 40512 9364 40540 9395
rect 40586 9392 40592 9444
rect 40644 9432 40650 9444
rect 42061 9435 42119 9441
rect 42061 9432 42073 9435
rect 40644 9404 42073 9432
rect 40644 9392 40650 9404
rect 42061 9401 42073 9404
rect 42107 9401 42119 9435
rect 42061 9395 42119 9401
rect 46658 9392 46664 9444
rect 46716 9432 46722 9444
rect 46845 9435 46903 9441
rect 46845 9432 46857 9435
rect 46716 9404 46857 9432
rect 46716 9392 46722 9404
rect 46845 9401 46857 9404
rect 46891 9401 46903 9435
rect 46845 9395 46903 9401
rect 48777 9435 48835 9441
rect 48777 9401 48789 9435
rect 48823 9432 48835 9435
rect 49418 9432 49424 9444
rect 48823 9404 49424 9432
rect 48823 9401 48835 9404
rect 48777 9395 48835 9401
rect 49418 9392 49424 9404
rect 49476 9392 49482 9444
rect 53466 9392 53472 9444
rect 53524 9432 53530 9444
rect 54849 9435 54907 9441
rect 54849 9432 54861 9435
rect 53524 9404 54861 9432
rect 53524 9392 53530 9404
rect 54849 9401 54861 9404
rect 54895 9401 54907 9435
rect 56226 9432 56232 9444
rect 56187 9404 56232 9432
rect 54849 9395 54907 9401
rect 56226 9392 56232 9404
rect 56284 9392 56290 9444
rect 57054 9432 57060 9444
rect 57015 9404 57060 9432
rect 57054 9392 57060 9404
rect 57112 9392 57118 9444
rect 57974 9432 57980 9444
rect 57935 9404 57980 9432
rect 57974 9392 57980 9404
rect 58032 9392 58038 9444
rect 42426 9364 42432 9376
rect 40512 9336 42432 9364
rect 42426 9324 42432 9336
rect 42484 9324 42490 9376
rect 54754 9324 54760 9376
rect 54812 9364 54818 9376
rect 59648 9364 59676 9540
rect 63586 9528 63592 9540
rect 63644 9528 63650 9580
rect 65613 9571 65671 9577
rect 65613 9537 65625 9571
rect 65659 9568 65671 9571
rect 65978 9568 65984 9580
rect 65659 9540 65984 9568
rect 65659 9537 65671 9540
rect 65613 9531 65671 9537
rect 65978 9528 65984 9540
rect 66036 9528 66042 9580
rect 66441 9571 66499 9577
rect 66441 9537 66453 9571
rect 66487 9568 66499 9571
rect 67269 9571 67327 9577
rect 66487 9540 67220 9568
rect 66487 9537 66499 9540
rect 66441 9531 66499 9537
rect 60090 9460 60096 9512
rect 60148 9500 60154 9512
rect 60642 9500 60648 9512
rect 60148 9472 60648 9500
rect 60148 9460 60154 9472
rect 60642 9460 60648 9472
rect 60700 9500 60706 9512
rect 62025 9503 62083 9509
rect 62025 9500 62037 9503
rect 60700 9472 62037 9500
rect 60700 9460 60706 9472
rect 62025 9469 62037 9472
rect 62071 9500 62083 9503
rect 63405 9503 63463 9509
rect 63405 9500 63417 9503
rect 62071 9472 63417 9500
rect 62071 9469 62083 9472
rect 62025 9463 62083 9469
rect 63405 9469 63417 9472
rect 63451 9469 63463 9503
rect 63405 9463 63463 9469
rect 64506 9460 64512 9512
rect 64564 9500 64570 9512
rect 64564 9472 65380 9500
rect 64564 9460 64570 9472
rect 61838 9432 61844 9444
rect 61799 9404 61844 9432
rect 61838 9392 61844 9404
rect 61896 9392 61902 9444
rect 62209 9435 62267 9441
rect 62209 9401 62221 9435
rect 62255 9401 62267 9435
rect 63218 9432 63224 9444
rect 63179 9404 63224 9432
rect 62209 9395 62267 9401
rect 54812 9336 59676 9364
rect 62224 9364 62252 9395
rect 63218 9392 63224 9404
rect 63276 9392 63282 9444
rect 65242 9432 65248 9444
rect 65203 9404 65248 9432
rect 65242 9392 65248 9404
rect 65300 9392 65306 9444
rect 65352 9432 65380 9472
rect 65426 9460 65432 9512
rect 65484 9500 65490 9512
rect 65794 9500 65800 9512
rect 65484 9472 65800 9500
rect 65484 9460 65490 9472
rect 65794 9460 65800 9472
rect 65852 9500 65858 9512
rect 66257 9503 66315 9509
rect 66257 9500 66269 9503
rect 65852 9472 66269 9500
rect 65852 9460 65858 9472
rect 66257 9469 66269 9472
rect 66303 9500 66315 9503
rect 67085 9503 67143 9509
rect 67085 9500 67097 9503
rect 66303 9472 67097 9500
rect 66303 9469 66315 9472
rect 66257 9463 66315 9469
rect 67085 9469 67097 9472
rect 67131 9469 67143 9503
rect 67192 9500 67220 9540
rect 67269 9537 67281 9571
rect 67315 9568 67327 9571
rect 67450 9568 67456 9580
rect 67315 9540 67456 9568
rect 67315 9537 67327 9540
rect 67269 9531 67327 9537
rect 67450 9528 67456 9540
rect 67508 9528 67514 9580
rect 69658 9500 69664 9512
rect 67192 9472 69664 9500
rect 67085 9463 67143 9469
rect 69658 9460 69664 9472
rect 69716 9460 69722 9512
rect 66073 9435 66131 9441
rect 66073 9432 66085 9435
rect 65352 9404 66085 9432
rect 66073 9401 66085 9404
rect 66119 9401 66131 9435
rect 66073 9395 66131 9401
rect 66901 9435 66959 9441
rect 66901 9401 66913 9435
rect 66947 9401 66959 9435
rect 66901 9395 66959 9401
rect 64782 9364 64788 9376
rect 62224 9336 64788 9364
rect 54812 9324 54818 9336
rect 64782 9324 64788 9336
rect 64840 9324 64846 9376
rect 65334 9324 65340 9376
rect 65392 9364 65398 9376
rect 66916 9364 66944 9395
rect 65392 9336 66944 9364
rect 65392 9324 65398 9336
rect 1104 9274 178848 9296
rect 1104 9222 19606 9274
rect 19658 9222 19670 9274
rect 19722 9222 19734 9274
rect 19786 9222 19798 9274
rect 19850 9222 50326 9274
rect 50378 9222 50390 9274
rect 50442 9222 50454 9274
rect 50506 9222 50518 9274
rect 50570 9222 81046 9274
rect 81098 9222 81110 9274
rect 81162 9222 81174 9274
rect 81226 9222 81238 9274
rect 81290 9222 111766 9274
rect 111818 9222 111830 9274
rect 111882 9222 111894 9274
rect 111946 9222 111958 9274
rect 112010 9222 142486 9274
rect 142538 9222 142550 9274
rect 142602 9222 142614 9274
rect 142666 9222 142678 9274
rect 142730 9222 173206 9274
rect 173258 9222 173270 9274
rect 173322 9222 173334 9274
rect 173386 9222 173398 9274
rect 173450 9222 178848 9274
rect 1104 9200 178848 9222
rect 48406 9160 48412 9172
rect 32784 9132 48412 9160
rect 32784 9101 32812 9132
rect 48406 9120 48412 9132
rect 48464 9160 48470 9172
rect 52086 9160 52092 9172
rect 48464 9132 52092 9160
rect 48464 9120 48470 9132
rect 52086 9120 52092 9132
rect 52144 9120 52150 9172
rect 61654 9160 61660 9172
rect 57946 9132 61660 9160
rect 32769 9095 32827 9101
rect 32769 9061 32781 9095
rect 32815 9061 32827 9095
rect 32769 9055 32827 9061
rect 41046 9052 41052 9104
rect 41104 9092 41110 9104
rect 57946 9092 57974 9132
rect 61654 9120 61660 9132
rect 61712 9120 61718 9172
rect 63681 9095 63739 9101
rect 41104 9064 57974 9092
rect 61396 9064 63540 9092
rect 41104 9052 41110 9064
rect 32582 9024 32588 9036
rect 32543 8996 32588 9024
rect 32582 8984 32588 8996
rect 32640 8984 32646 9036
rect 32861 9027 32919 9033
rect 32861 8993 32873 9027
rect 32907 8993 32919 9027
rect 32861 8987 32919 8993
rect 32953 9027 33011 9033
rect 32953 8993 32965 9027
rect 32999 9024 33011 9027
rect 33870 9024 33876 9036
rect 32999 8996 33876 9024
rect 32999 8993 33011 8996
rect 32953 8987 33011 8993
rect 30926 8916 30932 8968
rect 30984 8956 30990 8968
rect 32876 8956 32904 8987
rect 30984 8928 32904 8956
rect 30984 8916 30990 8928
rect 31386 8848 31392 8900
rect 31444 8888 31450 8900
rect 32968 8888 32996 8987
rect 33870 8984 33876 8996
rect 33928 8984 33934 9036
rect 40678 8984 40684 9036
rect 40736 9024 40742 9036
rect 54754 9024 54760 9036
rect 40736 8996 54760 9024
rect 40736 8984 40742 8996
rect 54754 8984 54760 8996
rect 54812 8984 54818 9036
rect 55030 8984 55036 9036
rect 55088 9024 55094 9036
rect 55401 9027 55459 9033
rect 55401 9024 55413 9027
rect 55088 8996 55413 9024
rect 55088 8984 55094 8996
rect 55401 8993 55413 8996
rect 55447 8993 55459 9027
rect 55401 8987 55459 8993
rect 55585 9027 55643 9033
rect 55585 8993 55597 9027
rect 55631 9024 55643 9027
rect 56870 9024 56876 9036
rect 55631 8996 56876 9024
rect 55631 8993 55643 8996
rect 55585 8987 55643 8993
rect 56870 8984 56876 8996
rect 56928 8984 56934 9036
rect 59538 8984 59544 9036
rect 59596 9024 59602 9036
rect 60553 9027 60611 9033
rect 60553 9024 60565 9027
rect 59596 8996 60565 9024
rect 59596 8984 59602 8996
rect 60553 8993 60565 8996
rect 60599 8993 60611 9027
rect 60553 8987 60611 8993
rect 60642 8984 60648 9036
rect 60700 9024 60706 9036
rect 60737 9027 60795 9033
rect 60737 9024 60749 9027
rect 60700 8996 60749 9024
rect 60700 8984 60706 8996
rect 60737 8993 60749 8996
rect 60783 9024 60795 9027
rect 61396 9024 61424 9064
rect 60783 8996 61424 9024
rect 60783 8993 60795 8996
rect 60737 8987 60795 8993
rect 61470 8984 61476 9036
rect 61528 9024 61534 9036
rect 62132 9033 62160 9064
rect 61933 9027 61991 9033
rect 61933 9024 61945 9027
rect 61528 8996 61945 9024
rect 61528 8984 61534 8996
rect 61933 8993 61945 8996
rect 61979 8993 61991 9027
rect 61933 8987 61991 8993
rect 62117 9027 62175 9033
rect 62117 8993 62129 9027
rect 62163 8993 62175 9027
rect 63310 9024 63316 9036
rect 63271 8996 63316 9024
rect 62117 8987 62175 8993
rect 63310 8984 63316 8996
rect 63368 8984 63374 9036
rect 63512 9033 63540 9064
rect 63681 9061 63693 9095
rect 63727 9092 63739 9095
rect 65518 9092 65524 9104
rect 63727 9064 65524 9092
rect 63727 9061 63739 9064
rect 63681 9055 63739 9061
rect 65518 9052 65524 9064
rect 65576 9052 65582 9104
rect 65981 9095 66039 9101
rect 65981 9061 65993 9095
rect 66027 9092 66039 9095
rect 66070 9092 66076 9104
rect 66027 9064 66076 9092
rect 66027 9061 66039 9064
rect 65981 9055 66039 9061
rect 66070 9052 66076 9064
rect 66128 9052 66134 9104
rect 63497 9027 63555 9033
rect 63497 8993 63509 9027
rect 63543 8993 63555 9027
rect 63497 8987 63555 8993
rect 63586 8984 63592 9036
rect 63644 9024 63650 9036
rect 65613 9027 65671 9033
rect 65613 9024 65625 9027
rect 63644 8996 65625 9024
rect 63644 8984 63650 8996
rect 65613 8993 65625 8996
rect 65659 8993 65671 9027
rect 65794 9024 65800 9036
rect 65755 8996 65800 9024
rect 65613 8987 65671 8993
rect 65794 8984 65800 8996
rect 65852 8984 65858 9036
rect 55766 8956 55772 8968
rect 55727 8928 55772 8956
rect 55766 8916 55772 8928
rect 55824 8916 55830 8968
rect 60921 8959 60979 8965
rect 60921 8925 60933 8959
rect 60967 8956 60979 8959
rect 62022 8956 62028 8968
rect 60967 8928 62028 8956
rect 60967 8925 60979 8928
rect 60921 8919 60979 8925
rect 62022 8916 62028 8928
rect 62080 8916 62086 8968
rect 62301 8959 62359 8965
rect 62301 8925 62313 8959
rect 62347 8956 62359 8959
rect 62942 8956 62948 8968
rect 62347 8928 62948 8956
rect 62347 8925 62359 8928
rect 62301 8919 62359 8925
rect 62942 8916 62948 8928
rect 63000 8916 63006 8968
rect 65058 8916 65064 8968
rect 65116 8956 65122 8968
rect 66990 8956 66996 8968
rect 65116 8928 66996 8956
rect 65116 8916 65122 8928
rect 66990 8916 66996 8928
rect 67048 8916 67054 8968
rect 31444 8860 32996 8888
rect 31444 8848 31450 8860
rect 38470 8848 38476 8900
rect 38528 8888 38534 8900
rect 41414 8888 41420 8900
rect 38528 8860 41420 8888
rect 38528 8848 38534 8860
rect 41414 8848 41420 8860
rect 41472 8848 41478 8900
rect 33137 8823 33195 8829
rect 33137 8789 33149 8823
rect 33183 8820 33195 8823
rect 33226 8820 33232 8832
rect 33183 8792 33232 8820
rect 33183 8789 33195 8792
rect 33137 8783 33195 8789
rect 33226 8780 33232 8792
rect 33284 8780 33290 8832
rect 33410 8780 33416 8832
rect 33468 8820 33474 8832
rect 49694 8820 49700 8832
rect 33468 8792 49700 8820
rect 33468 8780 33474 8792
rect 49694 8780 49700 8792
rect 49752 8780 49758 8832
rect 1104 8730 178848 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 34966 8730
rect 35018 8678 35030 8730
rect 35082 8678 35094 8730
rect 35146 8678 35158 8730
rect 35210 8678 65686 8730
rect 65738 8678 65750 8730
rect 65802 8678 65814 8730
rect 65866 8678 65878 8730
rect 65930 8678 96406 8730
rect 96458 8678 96470 8730
rect 96522 8678 96534 8730
rect 96586 8678 96598 8730
rect 96650 8678 127126 8730
rect 127178 8678 127190 8730
rect 127242 8678 127254 8730
rect 127306 8678 127318 8730
rect 127370 8678 157846 8730
rect 157898 8678 157910 8730
rect 157962 8678 157974 8730
rect 158026 8678 158038 8730
rect 158090 8678 178848 8730
rect 1104 8656 178848 8678
rect 33594 8576 33600 8628
rect 33652 8616 33658 8628
rect 41322 8616 41328 8628
rect 33652 8588 41328 8616
rect 33652 8576 33658 8588
rect 41322 8576 41328 8588
rect 41380 8576 41386 8628
rect 41414 8576 41420 8628
rect 41472 8616 41478 8628
rect 41472 8588 41517 8616
rect 41472 8576 41478 8588
rect 41598 8576 41604 8628
rect 41656 8616 41662 8628
rect 67634 8616 67640 8628
rect 41656 8588 67640 8616
rect 41656 8576 41662 8588
rect 67634 8576 67640 8588
rect 67692 8576 67698 8628
rect 33686 8508 33692 8560
rect 33744 8548 33750 8560
rect 33781 8551 33839 8557
rect 33781 8548 33793 8551
rect 33744 8520 33793 8548
rect 33744 8508 33750 8520
rect 33781 8517 33793 8520
rect 33827 8517 33839 8551
rect 33781 8511 33839 8517
rect 35618 8508 35624 8560
rect 35676 8548 35682 8560
rect 70026 8548 70032 8560
rect 35676 8520 70032 8548
rect 35676 8508 35682 8520
rect 70026 8508 70032 8520
rect 70084 8508 70090 8560
rect 31662 8440 31668 8492
rect 31720 8480 31726 8492
rect 31720 8452 35204 8480
rect 31720 8440 31726 8452
rect 31846 8372 31852 8424
rect 31904 8412 31910 8424
rect 32582 8412 32588 8424
rect 31904 8384 32588 8412
rect 31904 8372 31910 8384
rect 32582 8372 32588 8384
rect 32640 8412 32646 8424
rect 33042 8412 33048 8424
rect 32640 8384 33048 8412
rect 32640 8372 32646 8384
rect 33042 8372 33048 8384
rect 33100 8412 33106 8424
rect 33229 8415 33287 8421
rect 33229 8412 33241 8415
rect 33100 8384 33241 8412
rect 33100 8372 33106 8384
rect 33229 8381 33241 8384
rect 33275 8381 33287 8415
rect 33410 8412 33416 8424
rect 33371 8384 33416 8412
rect 33229 8375 33287 8381
rect 33410 8372 33416 8384
rect 33468 8372 33474 8424
rect 33597 8415 33655 8421
rect 33597 8381 33609 8415
rect 33643 8412 33655 8415
rect 33870 8412 33876 8424
rect 33643 8384 33876 8412
rect 33643 8381 33655 8384
rect 33597 8375 33655 8381
rect 33870 8372 33876 8384
rect 33928 8372 33934 8424
rect 35176 8421 35204 8452
rect 35894 8440 35900 8492
rect 35952 8480 35958 8492
rect 38286 8480 38292 8492
rect 35952 8452 38292 8480
rect 35952 8440 35958 8452
rect 38286 8440 38292 8452
rect 38344 8440 38350 8492
rect 39850 8440 39856 8492
rect 39908 8480 39914 8492
rect 65058 8480 65064 8492
rect 39908 8452 41184 8480
rect 39908 8440 39914 8452
rect 35161 8415 35219 8421
rect 35161 8381 35173 8415
rect 35207 8381 35219 8415
rect 35161 8375 35219 8381
rect 35345 8415 35403 8421
rect 35345 8381 35357 8415
rect 35391 8412 35403 8415
rect 39298 8412 39304 8424
rect 35391 8384 39304 8412
rect 35391 8381 35403 8384
rect 35345 8375 35403 8381
rect 39298 8372 39304 8384
rect 39356 8412 39362 8424
rect 40862 8412 40868 8424
rect 39356 8384 40868 8412
rect 39356 8372 39362 8384
rect 40862 8372 40868 8384
rect 40920 8372 40926 8424
rect 41046 8412 41052 8424
rect 41007 8384 41052 8412
rect 41046 8372 41052 8384
rect 41104 8372 41110 8424
rect 41156 8421 41184 8452
rect 46124 8452 65064 8480
rect 41141 8415 41199 8421
rect 41141 8381 41153 8415
rect 41187 8381 41199 8415
rect 41141 8375 41199 8381
rect 41230 8372 41236 8424
rect 41288 8412 41294 8424
rect 45554 8412 45560 8424
rect 41288 8384 41333 8412
rect 41432 8384 45560 8412
rect 41288 8372 41294 8384
rect 31938 8304 31944 8356
rect 31996 8344 32002 8356
rect 33505 8347 33563 8353
rect 33505 8344 33517 8347
rect 31996 8316 33517 8344
rect 31996 8304 32002 8316
rect 33505 8313 33517 8316
rect 33551 8313 33563 8347
rect 35894 8344 35900 8356
rect 35855 8316 35900 8344
rect 33505 8307 33563 8313
rect 35894 8304 35900 8316
rect 35952 8304 35958 8356
rect 36081 8347 36139 8353
rect 36081 8313 36093 8347
rect 36127 8344 36139 8347
rect 38654 8344 38660 8356
rect 36127 8316 38660 8344
rect 36127 8313 36139 8316
rect 36081 8307 36139 8313
rect 38654 8304 38660 8316
rect 38712 8304 38718 8356
rect 39482 8304 39488 8356
rect 39540 8344 39546 8356
rect 39540 8316 41368 8344
rect 39540 8304 39546 8316
rect 27798 8236 27804 8288
rect 27856 8276 27862 8288
rect 41046 8276 41052 8288
rect 27856 8248 41052 8276
rect 27856 8236 27862 8248
rect 41046 8236 41052 8248
rect 41104 8236 41110 8288
rect 41340 8276 41368 8316
rect 41432 8276 41460 8384
rect 45554 8372 45560 8384
rect 45612 8372 45618 8424
rect 45925 8415 45983 8421
rect 45925 8381 45937 8415
rect 45971 8412 45983 8415
rect 46014 8412 46020 8424
rect 45971 8384 46020 8412
rect 45971 8381 45983 8384
rect 45925 8375 45983 8381
rect 46014 8372 46020 8384
rect 46072 8372 46078 8424
rect 46124 8421 46152 8452
rect 65058 8440 65064 8452
rect 65116 8440 65122 8492
rect 46109 8415 46167 8421
rect 46109 8381 46121 8415
rect 46155 8381 46167 8415
rect 46290 8412 46296 8424
rect 46251 8384 46296 8412
rect 46109 8375 46167 8381
rect 46290 8372 46296 8384
rect 46348 8372 46354 8424
rect 63126 8372 63132 8424
rect 63184 8412 63190 8424
rect 67266 8412 67272 8424
rect 63184 8384 67272 8412
rect 63184 8372 63190 8384
rect 67266 8372 67272 8384
rect 67324 8372 67330 8424
rect 43254 8304 43260 8356
rect 43312 8344 43318 8356
rect 46201 8347 46259 8353
rect 46201 8344 46213 8347
rect 43312 8316 46213 8344
rect 43312 8304 43318 8316
rect 46201 8313 46213 8316
rect 46247 8313 46259 8347
rect 46201 8307 46259 8313
rect 54294 8304 54300 8356
rect 54352 8344 54358 8356
rect 56962 8344 56968 8356
rect 54352 8316 56968 8344
rect 54352 8304 54358 8316
rect 56962 8304 56968 8316
rect 57020 8304 57026 8356
rect 64414 8344 64420 8356
rect 62224 8316 64420 8344
rect 41340 8248 41460 8276
rect 45922 8236 45928 8288
rect 45980 8276 45986 8288
rect 46477 8279 46535 8285
rect 46477 8276 46489 8279
rect 45980 8248 46489 8276
rect 45980 8236 45986 8248
rect 46477 8245 46489 8248
rect 46523 8245 46535 8279
rect 46477 8239 46535 8245
rect 46566 8236 46572 8288
rect 46624 8276 46630 8288
rect 55674 8276 55680 8288
rect 46624 8248 55680 8276
rect 46624 8236 46630 8248
rect 55674 8236 55680 8248
rect 55732 8236 55738 8288
rect 55766 8236 55772 8288
rect 55824 8276 55830 8288
rect 62224 8276 62252 8316
rect 64414 8304 64420 8316
rect 64472 8304 64478 8356
rect 55824 8248 62252 8276
rect 55824 8236 55830 8248
rect 62298 8236 62304 8288
rect 62356 8276 62362 8288
rect 68646 8276 68652 8288
rect 62356 8248 68652 8276
rect 62356 8236 62362 8248
rect 68646 8236 68652 8248
rect 68704 8276 68710 8288
rect 71314 8276 71320 8288
rect 68704 8248 71320 8276
rect 68704 8236 68710 8248
rect 71314 8236 71320 8248
rect 71372 8236 71378 8288
rect 1104 8186 178848 8208
rect 1104 8134 19606 8186
rect 19658 8134 19670 8186
rect 19722 8134 19734 8186
rect 19786 8134 19798 8186
rect 19850 8134 50326 8186
rect 50378 8134 50390 8186
rect 50442 8134 50454 8186
rect 50506 8134 50518 8186
rect 50570 8134 81046 8186
rect 81098 8134 81110 8186
rect 81162 8134 81174 8186
rect 81226 8134 81238 8186
rect 81290 8134 111766 8186
rect 111818 8134 111830 8186
rect 111882 8134 111894 8186
rect 111946 8134 111958 8186
rect 112010 8134 142486 8186
rect 142538 8134 142550 8186
rect 142602 8134 142614 8186
rect 142666 8134 142678 8186
rect 142730 8134 173206 8186
rect 173258 8134 173270 8186
rect 173322 8134 173334 8186
rect 173386 8134 173398 8186
rect 173450 8134 178848 8186
rect 1104 8112 178848 8134
rect 31570 8072 31576 8084
rect 25792 8044 31576 8072
rect 20990 8004 20996 8016
rect 20951 7976 20996 8004
rect 20990 7964 20996 7976
rect 21048 7964 21054 8016
rect 21085 8007 21143 8013
rect 21085 7973 21097 8007
rect 21131 8004 21143 8007
rect 21266 8004 21272 8016
rect 21131 7976 21272 8004
rect 21131 7973 21143 7976
rect 21085 7967 21143 7973
rect 21266 7964 21272 7976
rect 21324 7964 21330 8016
rect 24210 7964 24216 8016
rect 24268 8004 24274 8016
rect 25792 8013 25820 8044
rect 31570 8032 31576 8044
rect 31628 8032 31634 8084
rect 33594 8072 33600 8084
rect 31726 8044 33456 8072
rect 33555 8044 33600 8072
rect 25777 8007 25835 8013
rect 24268 7976 25728 8004
rect 24268 7964 24274 7976
rect 20809 7939 20867 7945
rect 20809 7905 20821 7939
rect 20855 7905 20867 7939
rect 20809 7899 20867 7905
rect 20824 7868 20852 7899
rect 21174 7896 21180 7948
rect 21232 7936 21238 7948
rect 25590 7936 25596 7948
rect 21232 7908 21277 7936
rect 25551 7908 25596 7936
rect 21232 7896 21238 7908
rect 25590 7896 25596 7908
rect 25648 7896 25654 7948
rect 25700 7936 25728 7976
rect 25777 7973 25789 8007
rect 25823 7973 25835 8007
rect 27798 8004 27804 8016
rect 27759 7976 27804 8004
rect 25777 7967 25835 7973
rect 27798 7964 27804 7976
rect 27856 7964 27862 8016
rect 28166 7964 28172 8016
rect 28224 8004 28230 8016
rect 29914 8004 29920 8016
rect 28224 7976 29920 8004
rect 28224 7964 28230 7976
rect 29914 7964 29920 7976
rect 29972 7964 29978 8016
rect 30374 7964 30380 8016
rect 30432 8004 30438 8016
rect 30653 8007 30711 8013
rect 30432 7976 30604 8004
rect 30432 7964 30438 7976
rect 25869 7939 25927 7945
rect 25869 7936 25881 7939
rect 25700 7908 25881 7936
rect 25869 7905 25881 7908
rect 25915 7905 25927 7939
rect 25869 7899 25927 7905
rect 25958 7896 25964 7948
rect 26016 7936 26022 7948
rect 26016 7908 26061 7936
rect 26016 7896 26022 7908
rect 26418 7896 26424 7948
rect 26476 7936 26482 7948
rect 27614 7936 27620 7948
rect 26476 7908 27620 7936
rect 26476 7896 26482 7908
rect 27614 7896 27620 7908
rect 27672 7936 27678 7948
rect 27890 7936 27896 7948
rect 27672 7908 27717 7936
rect 27851 7908 27896 7936
rect 27672 7896 27678 7908
rect 27890 7896 27896 7908
rect 27948 7896 27954 7948
rect 27985 7939 28043 7945
rect 27985 7905 27997 7939
rect 28031 7905 28043 7939
rect 27985 7899 28043 7905
rect 20990 7868 20996 7880
rect 20824 7840 20996 7868
rect 20990 7828 20996 7840
rect 21048 7828 21054 7880
rect 25976 7868 26004 7896
rect 28000 7868 28028 7899
rect 28258 7896 28264 7948
rect 28316 7936 28322 7948
rect 28721 7939 28779 7945
rect 28721 7936 28733 7939
rect 28316 7908 28733 7936
rect 28316 7896 28322 7908
rect 28721 7905 28733 7908
rect 28767 7936 28779 7939
rect 29362 7936 29368 7948
rect 28767 7908 29368 7936
rect 28767 7905 28779 7908
rect 28721 7899 28779 7905
rect 29362 7896 29368 7908
rect 29420 7896 29426 7948
rect 30466 7936 30472 7948
rect 30427 7908 30472 7936
rect 30466 7896 30472 7908
rect 30524 7896 30530 7948
rect 30576 7936 30604 7976
rect 30653 7973 30665 8007
rect 30699 8004 30711 8007
rect 31726 8004 31754 8044
rect 31846 8004 31852 8016
rect 30699 7976 31754 8004
rect 31807 7976 31852 8004
rect 30699 7973 30711 7976
rect 30653 7967 30711 7973
rect 31846 7964 31852 7976
rect 31904 7964 31910 8016
rect 32490 8004 32496 8016
rect 32451 7976 32496 8004
rect 32490 7964 32496 7976
rect 32548 7964 32554 8016
rect 32582 7964 32588 8016
rect 32640 8004 32646 8016
rect 32769 8007 32827 8013
rect 32769 8004 32781 8007
rect 32640 7976 32781 8004
rect 32640 7964 32646 7976
rect 32769 7973 32781 7976
rect 32815 7973 32827 8007
rect 32769 7967 32827 7973
rect 32950 7964 32956 8016
rect 33008 8004 33014 8016
rect 33229 8007 33287 8013
rect 33229 8004 33241 8007
rect 33008 7976 33241 8004
rect 33008 7964 33014 7976
rect 33229 7973 33241 7976
rect 33275 7973 33287 8007
rect 33428 8004 33456 8044
rect 33594 8032 33600 8044
rect 33652 8032 33658 8084
rect 33778 8072 33784 8084
rect 33739 8044 33784 8072
rect 33778 8032 33784 8044
rect 33836 8032 33842 8084
rect 33962 8032 33968 8084
rect 34020 8072 34026 8084
rect 39482 8072 39488 8084
rect 34020 8044 39488 8072
rect 34020 8032 34026 8044
rect 39482 8032 39488 8044
rect 39540 8032 39546 8084
rect 46014 8072 46020 8084
rect 39684 8044 46020 8072
rect 33428 7976 33732 8004
rect 33229 7967 33287 7973
rect 30745 7939 30803 7945
rect 30745 7936 30757 7939
rect 30576 7908 30757 7936
rect 30745 7905 30757 7908
rect 30791 7905 30803 7939
rect 30745 7899 30803 7905
rect 30837 7939 30895 7945
rect 30837 7905 30849 7939
rect 30883 7936 30895 7939
rect 31018 7936 31024 7948
rect 30883 7908 31024 7936
rect 30883 7905 30895 7908
rect 30837 7899 30895 7905
rect 31018 7896 31024 7908
rect 31076 7936 31082 7948
rect 31386 7936 31392 7948
rect 31076 7908 31392 7936
rect 31076 7896 31082 7908
rect 31386 7896 31392 7908
rect 31444 7896 31450 7948
rect 31662 7936 31668 7948
rect 31575 7908 31668 7936
rect 31662 7896 31668 7908
rect 31720 7896 31726 7948
rect 32858 7936 32864 7948
rect 32819 7908 32864 7936
rect 32858 7896 32864 7908
rect 32916 7896 32922 7948
rect 28810 7868 28816 7880
rect 25976 7840 28816 7868
rect 28810 7828 28816 7840
rect 28868 7868 28874 7880
rect 28905 7871 28963 7877
rect 28905 7868 28917 7871
rect 28868 7840 28917 7868
rect 28868 7828 28874 7840
rect 28905 7837 28917 7840
rect 28951 7837 28963 7871
rect 28905 7831 28963 7837
rect 29178 7828 29184 7880
rect 29236 7868 29242 7880
rect 31680 7868 31708 7896
rect 29236 7840 31708 7868
rect 29236 7828 29242 7840
rect 33318 7828 33324 7880
rect 33376 7828 33382 7880
rect 26234 7760 26240 7812
rect 26292 7800 26298 7812
rect 28258 7800 28264 7812
rect 26292 7772 28264 7800
rect 26292 7760 26298 7772
rect 28258 7760 28264 7772
rect 28316 7760 28322 7812
rect 20806 7692 20812 7744
rect 20864 7732 20870 7744
rect 21361 7735 21419 7741
rect 21361 7732 21373 7735
rect 20864 7704 21373 7732
rect 20864 7692 20870 7704
rect 21361 7701 21373 7704
rect 21407 7701 21419 7735
rect 21361 7695 21419 7701
rect 23474 7692 23480 7744
rect 23532 7732 23538 7744
rect 26145 7735 26203 7741
rect 26145 7732 26157 7735
rect 23532 7704 26157 7732
rect 23532 7692 23538 7704
rect 26145 7701 26157 7704
rect 26191 7701 26203 7735
rect 26145 7695 26203 7701
rect 26326 7692 26332 7744
rect 26384 7732 26390 7744
rect 28169 7735 28227 7741
rect 28169 7732 28181 7735
rect 26384 7704 28181 7732
rect 26384 7692 26390 7704
rect 28169 7701 28181 7704
rect 28215 7701 28227 7735
rect 28169 7695 28227 7701
rect 29270 7692 29276 7744
rect 29328 7732 29334 7744
rect 31021 7735 31079 7741
rect 31021 7732 31033 7735
rect 29328 7704 31033 7732
rect 29328 7692 29334 7704
rect 31021 7701 31033 7704
rect 31067 7701 31079 7735
rect 33704 7732 33732 7976
rect 34330 7964 34336 8016
rect 34388 8004 34394 8016
rect 36354 8004 36360 8016
rect 34388 7976 36360 8004
rect 34388 7964 34394 7976
rect 36354 7964 36360 7976
rect 36412 7964 36418 8016
rect 38286 8004 38292 8016
rect 38247 7976 38292 8004
rect 38286 7964 38292 7976
rect 38344 8004 38350 8016
rect 38562 8004 38568 8016
rect 38344 7976 38568 8004
rect 38344 7964 38350 7976
rect 38562 7964 38568 7976
rect 38620 7964 38626 8016
rect 39298 7964 39304 8016
rect 39356 8004 39362 8016
rect 39684 8013 39712 8044
rect 46014 8032 46020 8044
rect 46072 8032 46078 8084
rect 46842 8072 46848 8084
rect 46308 8044 46848 8072
rect 46308 8016 46336 8044
rect 46814 8032 46848 8044
rect 46900 8072 46906 8084
rect 55766 8072 55772 8084
rect 46900 8044 47808 8072
rect 46900 8032 46906 8044
rect 39669 8007 39727 8013
rect 39356 7976 39528 8004
rect 39356 7964 39362 7976
rect 35986 7896 35992 7948
rect 36044 7936 36050 7948
rect 36449 7939 36507 7945
rect 36449 7936 36461 7939
rect 36044 7908 36461 7936
rect 36044 7896 36050 7908
rect 36449 7905 36461 7908
rect 36495 7905 36507 7939
rect 36449 7899 36507 7905
rect 37458 7896 37464 7948
rect 37516 7936 37522 7948
rect 39500 7945 39528 7976
rect 39669 7973 39681 8007
rect 39715 7973 39727 8007
rect 39669 7967 39727 7973
rect 40862 7964 40868 8016
rect 40920 8004 40926 8016
rect 41874 8004 41880 8016
rect 40920 7976 41736 8004
rect 41835 7976 41880 8004
rect 40920 7964 40926 7976
rect 41708 7948 41736 7976
rect 41874 7964 41880 7976
rect 41932 7964 41938 8016
rect 41966 7964 41972 8016
rect 42024 8004 42030 8016
rect 42024 7976 42069 8004
rect 42024 7964 42030 7976
rect 43990 7964 43996 8016
rect 44048 8004 44054 8016
rect 46290 8004 46296 8016
rect 44048 7976 46296 8004
rect 44048 7964 44054 7976
rect 46290 7964 46296 7976
rect 46348 7964 46354 8016
rect 39485 7939 39543 7945
rect 37516 7908 39436 7936
rect 37516 7896 37522 7908
rect 33870 7828 33876 7880
rect 33928 7868 33934 7880
rect 36633 7871 36691 7877
rect 33928 7840 36492 7868
rect 33928 7828 33934 7840
rect 33778 7760 33784 7812
rect 33836 7800 33842 7812
rect 36354 7800 36360 7812
rect 33836 7772 36360 7800
rect 33836 7760 33842 7772
rect 36354 7760 36360 7772
rect 36412 7760 36418 7812
rect 36464 7800 36492 7840
rect 36633 7837 36645 7871
rect 36679 7868 36691 7871
rect 39114 7868 39120 7880
rect 36679 7840 39120 7868
rect 36679 7837 36691 7840
rect 36633 7831 36691 7837
rect 39114 7828 39120 7840
rect 39172 7828 39178 7880
rect 39408 7868 39436 7908
rect 39485 7905 39497 7939
rect 39531 7905 39543 7939
rect 39485 7899 39543 7905
rect 39761 7939 39819 7945
rect 39761 7905 39773 7939
rect 39807 7905 39819 7939
rect 39761 7899 39819 7905
rect 39853 7939 39911 7945
rect 39853 7905 39865 7939
rect 39899 7936 39911 7939
rect 39942 7936 39948 7948
rect 39899 7908 39948 7936
rect 39899 7905 39911 7908
rect 39853 7899 39911 7905
rect 39776 7868 39804 7899
rect 39942 7896 39948 7908
rect 40000 7896 40006 7948
rect 40126 7896 40132 7948
rect 40184 7936 40190 7948
rect 40957 7939 41015 7945
rect 40957 7936 40969 7939
rect 40184 7908 40969 7936
rect 40184 7896 40190 7908
rect 40957 7905 40969 7908
rect 41003 7905 41015 7939
rect 41598 7936 41604 7948
rect 40957 7899 41015 7905
rect 41064 7908 41604 7936
rect 39408 7840 39804 7868
rect 40034 7828 40040 7880
rect 40092 7868 40098 7880
rect 41064 7868 41092 7908
rect 41598 7896 41604 7908
rect 41656 7896 41662 7948
rect 41690 7896 41696 7948
rect 41748 7936 41754 7948
rect 42061 7939 42119 7945
rect 41748 7908 41793 7936
rect 41748 7896 41754 7908
rect 42061 7905 42073 7939
rect 42107 7905 42119 7939
rect 42061 7899 42119 7905
rect 40092 7840 41092 7868
rect 40092 7828 40098 7840
rect 41230 7828 41236 7880
rect 41288 7868 41294 7880
rect 42076 7868 42104 7899
rect 44174 7896 44180 7948
rect 44232 7936 44238 7948
rect 44545 7939 44603 7945
rect 44545 7936 44557 7939
rect 44232 7908 44557 7936
rect 44232 7896 44238 7908
rect 44545 7905 44557 7908
rect 44591 7905 44603 7939
rect 46382 7936 46388 7948
rect 46343 7908 46388 7936
rect 44545 7899 44603 7905
rect 46382 7896 46388 7908
rect 46440 7896 46446 7948
rect 46566 7936 46572 7948
rect 46527 7908 46572 7936
rect 46566 7896 46572 7908
rect 46624 7896 46630 7948
rect 46814 7945 46842 8032
rect 46661 7939 46719 7945
rect 46661 7905 46673 7939
rect 46707 7905 46719 7939
rect 46661 7899 46719 7905
rect 46799 7939 46857 7945
rect 46799 7905 46811 7939
rect 46845 7905 46857 7939
rect 46799 7899 46857 7905
rect 41288 7840 42104 7868
rect 41288 7828 41294 7840
rect 45094 7828 45100 7880
rect 45152 7868 45158 7880
rect 46676 7868 46704 7899
rect 47302 7896 47308 7948
rect 47360 7936 47366 7948
rect 47397 7939 47455 7945
rect 47397 7936 47409 7939
rect 47360 7908 47409 7936
rect 47360 7896 47366 7908
rect 47397 7905 47409 7908
rect 47443 7905 47455 7939
rect 47397 7899 47455 7905
rect 47486 7896 47492 7948
rect 47544 7945 47550 7948
rect 47544 7939 47593 7945
rect 47544 7905 47547 7939
rect 47581 7905 47593 7939
rect 47670 7936 47676 7948
rect 47631 7908 47676 7936
rect 47544 7899 47593 7905
rect 47544 7896 47550 7899
rect 47670 7896 47676 7908
rect 47728 7896 47734 7948
rect 47780 7945 47808 8044
rect 48608 8044 55772 8072
rect 47946 7964 47952 8016
rect 48004 8004 48010 8016
rect 48498 8004 48504 8016
rect 48004 7976 48504 8004
rect 48004 7964 48010 7976
rect 48498 7964 48504 7976
rect 48556 7964 48562 8016
rect 48608 8013 48636 8044
rect 55766 8032 55772 8044
rect 55824 8032 55830 8084
rect 55858 8032 55864 8084
rect 55916 8072 55922 8084
rect 60550 8072 60556 8084
rect 55916 8044 60556 8072
rect 55916 8032 55922 8044
rect 60550 8032 60556 8044
rect 60608 8032 60614 8084
rect 63126 8072 63132 8084
rect 62592 8044 63132 8072
rect 48593 8007 48651 8013
rect 48593 7973 48605 8007
rect 48639 7973 48651 8007
rect 48593 7967 48651 7973
rect 48682 7964 48688 8016
rect 48740 8004 48746 8016
rect 48740 7976 48785 8004
rect 48740 7964 48746 7976
rect 54754 7964 54760 8016
rect 54812 8004 54818 8016
rect 58066 8004 58072 8016
rect 54812 7976 58072 8004
rect 54812 7964 54818 7976
rect 58066 7964 58072 7976
rect 58124 8004 58130 8016
rect 59446 8004 59452 8016
rect 58124 7976 59452 8004
rect 58124 7964 58130 7976
rect 59446 7964 59452 7976
rect 59504 7964 59510 8016
rect 47765 7939 47823 7945
rect 47765 7905 47777 7939
rect 47811 7905 47823 7939
rect 48406 7936 48412 7948
rect 48367 7908 48412 7936
rect 47765 7899 47823 7905
rect 48406 7896 48412 7908
rect 48464 7896 48470 7948
rect 48777 7939 48835 7945
rect 48777 7905 48789 7939
rect 48823 7936 48835 7939
rect 49142 7936 49148 7948
rect 48823 7908 49148 7936
rect 48823 7905 48835 7908
rect 48777 7899 48835 7905
rect 49142 7896 49148 7908
rect 49200 7896 49206 7948
rect 49970 7896 49976 7948
rect 50028 7936 50034 7948
rect 62298 7936 62304 7948
rect 50028 7908 62304 7936
rect 50028 7896 50034 7908
rect 62298 7896 62304 7908
rect 62356 7896 62362 7948
rect 62592 7945 62620 8044
rect 63126 8032 63132 8044
rect 63184 8032 63190 8084
rect 64417 8075 64475 8081
rect 64417 8041 64429 8075
rect 64463 8072 64475 8075
rect 65334 8072 65340 8084
rect 64463 8044 65340 8072
rect 64463 8041 64475 8044
rect 64417 8035 64475 8041
rect 65334 8032 65340 8044
rect 65392 8032 65398 8084
rect 62577 7939 62635 7945
rect 62577 7905 62589 7939
rect 62623 7905 62635 7939
rect 62577 7899 62635 7905
rect 63494 7896 63500 7948
rect 63552 7945 63558 7948
rect 63552 7939 63573 7945
rect 63561 7905 63573 7939
rect 63614 7939 63672 7945
rect 63614 7936 63626 7939
rect 63552 7899 63573 7905
rect 63604 7905 63626 7936
rect 63660 7905 63672 7939
rect 63604 7899 63672 7905
rect 63552 7896 63558 7899
rect 45152 7840 46704 7868
rect 45152 7828 45158 7840
rect 46934 7828 46940 7880
rect 46992 7868 46998 7880
rect 56686 7868 56692 7880
rect 46992 7840 56692 7868
rect 46992 7828 46998 7840
rect 56686 7828 56692 7840
rect 56744 7828 56750 7880
rect 62390 7828 62396 7880
rect 62448 7868 62454 7880
rect 62666 7868 62672 7880
rect 62448 7840 62672 7868
rect 62448 7828 62454 7840
rect 62666 7828 62672 7840
rect 62724 7828 62730 7880
rect 62761 7871 62819 7877
rect 62761 7837 62773 7871
rect 62807 7868 62819 7871
rect 62942 7868 62948 7880
rect 62807 7840 62948 7868
rect 62807 7837 62819 7840
rect 62761 7831 62819 7837
rect 62942 7828 62948 7840
rect 63000 7828 63006 7880
rect 63126 7828 63132 7880
rect 63184 7868 63190 7880
rect 63604 7868 63632 7899
rect 64414 7896 64420 7948
rect 64472 7936 64478 7948
rect 68554 7936 68560 7948
rect 64472 7908 68560 7936
rect 64472 7896 64478 7908
rect 68554 7896 68560 7908
rect 68612 7936 68618 7948
rect 72602 7936 72608 7948
rect 68612 7908 72608 7936
rect 68612 7896 68618 7908
rect 72602 7896 72608 7908
rect 72660 7896 72666 7948
rect 63184 7840 63632 7868
rect 63773 7871 63831 7877
rect 63184 7828 63190 7840
rect 63773 7837 63785 7871
rect 63819 7868 63831 7871
rect 64138 7868 64144 7880
rect 63819 7840 64144 7868
rect 63819 7837 63831 7840
rect 63773 7831 63831 7837
rect 64138 7828 64144 7840
rect 64196 7868 64202 7880
rect 65518 7868 65524 7880
rect 64196 7840 65524 7868
rect 64196 7828 64202 7840
rect 65518 7828 65524 7840
rect 65576 7828 65582 7880
rect 36722 7800 36728 7812
rect 36464 7772 36728 7800
rect 36722 7760 36728 7772
rect 36780 7760 36786 7812
rect 38473 7803 38531 7809
rect 38473 7769 38485 7803
rect 38519 7800 38531 7803
rect 40862 7800 40868 7812
rect 38519 7772 40868 7800
rect 38519 7769 38531 7772
rect 38473 7763 38531 7769
rect 40862 7760 40868 7772
rect 40920 7760 40926 7812
rect 40954 7760 40960 7812
rect 41012 7800 41018 7812
rect 41141 7803 41199 7809
rect 41141 7800 41153 7803
rect 41012 7772 41153 7800
rect 41012 7760 41018 7772
rect 41141 7769 41153 7772
rect 41187 7769 41199 7803
rect 41141 7763 41199 7769
rect 41506 7760 41512 7812
rect 41564 7800 41570 7812
rect 46566 7800 46572 7812
rect 41564 7772 46572 7800
rect 41564 7760 41570 7772
rect 46566 7760 46572 7772
rect 46624 7760 46630 7812
rect 47486 7760 47492 7812
rect 47544 7800 47550 7812
rect 50982 7800 50988 7812
rect 47544 7772 50988 7800
rect 47544 7760 47550 7772
rect 50982 7760 50988 7772
rect 51040 7760 51046 7812
rect 55214 7760 55220 7812
rect 55272 7800 55278 7812
rect 56870 7800 56876 7812
rect 55272 7772 56876 7800
rect 55272 7760 55278 7772
rect 56870 7760 56876 7772
rect 56928 7760 56934 7812
rect 61102 7760 61108 7812
rect 61160 7800 61166 7812
rect 62574 7800 62580 7812
rect 61160 7772 62580 7800
rect 61160 7760 61166 7772
rect 62574 7760 62580 7772
rect 62632 7760 62638 7812
rect 62850 7760 62856 7812
rect 62908 7800 62914 7812
rect 63221 7803 63279 7809
rect 63221 7800 63233 7803
rect 62908 7772 63233 7800
rect 62908 7760 62914 7772
rect 63221 7769 63233 7772
rect 63267 7769 63279 7803
rect 63221 7763 63279 7769
rect 64230 7760 64236 7812
rect 64288 7800 64294 7812
rect 70118 7800 70124 7812
rect 64288 7772 70124 7800
rect 64288 7760 64294 7772
rect 70118 7760 70124 7772
rect 70176 7800 70182 7812
rect 70302 7800 70308 7812
rect 70176 7772 70308 7800
rect 70176 7760 70182 7772
rect 70302 7760 70308 7772
rect 70360 7760 70366 7812
rect 39942 7732 39948 7744
rect 33704 7704 39948 7732
rect 31021 7695 31079 7701
rect 39942 7692 39948 7704
rect 40000 7692 40006 7744
rect 40037 7735 40095 7741
rect 40037 7701 40049 7735
rect 40083 7732 40095 7735
rect 40126 7732 40132 7744
rect 40083 7704 40132 7732
rect 40083 7701 40095 7704
rect 40037 7695 40095 7701
rect 40126 7692 40132 7704
rect 40184 7692 40190 7744
rect 40218 7692 40224 7744
rect 40276 7732 40282 7744
rect 42245 7735 42303 7741
rect 42245 7732 42257 7735
rect 40276 7704 42257 7732
rect 40276 7692 40282 7704
rect 42245 7701 42257 7704
rect 42291 7701 42303 7735
rect 42245 7695 42303 7701
rect 44361 7735 44419 7741
rect 44361 7701 44373 7735
rect 44407 7732 44419 7735
rect 44726 7732 44732 7744
rect 44407 7704 44732 7732
rect 44407 7701 44419 7704
rect 44361 7695 44419 7701
rect 44726 7692 44732 7704
rect 44784 7692 44790 7744
rect 46937 7735 46995 7741
rect 46937 7701 46949 7735
rect 46983 7732 46995 7735
rect 47302 7732 47308 7744
rect 46983 7704 47308 7732
rect 46983 7701 46995 7704
rect 46937 7695 46995 7701
rect 47302 7692 47308 7704
rect 47360 7692 47366 7744
rect 47949 7735 48007 7741
rect 47949 7701 47961 7735
rect 47995 7732 48007 7735
rect 48130 7732 48136 7744
rect 47995 7704 48136 7732
rect 47995 7701 48007 7704
rect 47949 7695 48007 7701
rect 48130 7692 48136 7704
rect 48188 7692 48194 7744
rect 48774 7692 48780 7744
rect 48832 7732 48838 7744
rect 48961 7735 49019 7741
rect 48961 7732 48973 7735
rect 48832 7704 48973 7732
rect 48832 7692 48838 7704
rect 48961 7701 48973 7704
rect 49007 7701 49019 7735
rect 48961 7695 49019 7701
rect 49050 7692 49056 7744
rect 49108 7732 49114 7744
rect 65426 7732 65432 7744
rect 49108 7704 65432 7732
rect 49108 7692 49114 7704
rect 65426 7692 65432 7704
rect 65484 7692 65490 7744
rect 1104 7642 178848 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 34966 7642
rect 35018 7590 35030 7642
rect 35082 7590 35094 7642
rect 35146 7590 35158 7642
rect 35210 7590 65686 7642
rect 65738 7590 65750 7642
rect 65802 7590 65814 7642
rect 65866 7590 65878 7642
rect 65930 7590 96406 7642
rect 96458 7590 96470 7642
rect 96522 7590 96534 7642
rect 96586 7590 96598 7642
rect 96650 7590 127126 7642
rect 127178 7590 127190 7642
rect 127242 7590 127254 7642
rect 127306 7590 127318 7642
rect 127370 7590 157846 7642
rect 157898 7590 157910 7642
rect 157962 7590 157974 7642
rect 158026 7590 158038 7642
rect 158090 7590 178848 7642
rect 1104 7568 178848 7590
rect 22186 7528 22192 7540
rect 18892 7500 22192 7528
rect 18598 7324 18604 7336
rect 18559 7296 18604 7324
rect 18598 7284 18604 7296
rect 18656 7284 18662 7336
rect 18785 7327 18843 7333
rect 18785 7293 18797 7327
rect 18831 7324 18843 7327
rect 18892 7324 18920 7500
rect 22186 7488 22192 7500
rect 22244 7488 22250 7540
rect 29638 7528 29644 7540
rect 22296 7500 29500 7528
rect 29551 7500 29644 7528
rect 22296 7392 22324 7500
rect 29472 7460 29500 7500
rect 29638 7488 29644 7500
rect 29696 7528 29702 7540
rect 30466 7528 30472 7540
rect 29696 7500 30472 7528
rect 29696 7488 29702 7500
rect 30466 7488 30472 7500
rect 30524 7488 30530 7540
rect 32122 7528 32128 7540
rect 30559 7500 32128 7528
rect 30559 7460 30587 7500
rect 32122 7488 32128 7500
rect 32180 7488 32186 7540
rect 35802 7528 35808 7540
rect 35763 7500 35808 7528
rect 35802 7488 35808 7500
rect 35860 7488 35866 7540
rect 36170 7488 36176 7540
rect 36228 7528 36234 7540
rect 39390 7528 39396 7540
rect 36228 7500 39396 7528
rect 36228 7488 36234 7500
rect 39390 7488 39396 7500
rect 39448 7488 39454 7540
rect 40770 7488 40776 7540
rect 40828 7528 40834 7540
rect 40865 7531 40923 7537
rect 40865 7528 40877 7531
rect 40828 7500 40877 7528
rect 40828 7488 40834 7500
rect 40865 7497 40877 7500
rect 40911 7497 40923 7531
rect 40865 7491 40923 7497
rect 40954 7488 40960 7540
rect 41012 7528 41018 7540
rect 50890 7528 50896 7540
rect 41012 7500 50896 7528
rect 41012 7488 41018 7500
rect 50890 7488 50896 7500
rect 50948 7488 50954 7540
rect 50982 7488 50988 7540
rect 51040 7528 51046 7540
rect 56689 7531 56747 7537
rect 51040 7500 56456 7528
rect 51040 7488 51046 7500
rect 27586 7432 28856 7460
rect 29472 7432 30587 7460
rect 25958 7392 25964 7404
rect 20364 7364 22324 7392
rect 23400 7364 25964 7392
rect 18831 7296 18920 7324
rect 18831 7293 18843 7296
rect 18785 7287 18843 7293
rect 18966 7284 18972 7336
rect 19024 7324 19030 7336
rect 20162 7324 20168 7336
rect 19024 7296 19334 7324
rect 20123 7296 20168 7324
rect 19024 7284 19030 7296
rect 18046 7216 18052 7268
rect 18104 7256 18110 7268
rect 18877 7259 18935 7265
rect 18877 7256 18889 7259
rect 18104 7228 18889 7256
rect 18104 7216 18110 7228
rect 18877 7225 18889 7228
rect 18923 7225 18935 7259
rect 18877 7219 18935 7225
rect 17954 7148 17960 7200
rect 18012 7188 18018 7200
rect 19153 7191 19211 7197
rect 19153 7188 19165 7191
rect 18012 7160 19165 7188
rect 18012 7148 18018 7160
rect 19153 7157 19165 7160
rect 19199 7157 19211 7191
rect 19306 7188 19334 7296
rect 20162 7284 20168 7296
rect 20220 7284 20226 7336
rect 20364 7333 20392 7364
rect 20349 7327 20407 7333
rect 20349 7293 20361 7327
rect 20395 7293 20407 7327
rect 20349 7287 20407 7293
rect 20533 7327 20591 7333
rect 20533 7293 20545 7327
rect 20579 7324 20591 7327
rect 20898 7324 20904 7336
rect 20579 7296 20904 7324
rect 20579 7293 20591 7296
rect 20533 7287 20591 7293
rect 20438 7256 20444 7268
rect 20399 7228 20444 7256
rect 20438 7216 20444 7228
rect 20496 7216 20502 7268
rect 20548 7188 20576 7287
rect 20898 7284 20904 7296
rect 20956 7284 20962 7336
rect 23014 7324 23020 7336
rect 22975 7296 23020 7324
rect 23014 7284 23020 7296
rect 23072 7284 23078 7336
rect 23400 7333 23428 7364
rect 25958 7352 25964 7364
rect 26016 7392 26022 7404
rect 26016 7364 26740 7392
rect 26016 7352 26022 7364
rect 23293 7327 23351 7333
rect 23293 7324 23305 7327
rect 23124 7296 23305 7324
rect 22002 7216 22008 7268
rect 22060 7256 22066 7268
rect 23124 7256 23152 7296
rect 23293 7293 23305 7296
rect 23339 7293 23351 7327
rect 23293 7287 23351 7293
rect 23385 7327 23443 7333
rect 23385 7293 23397 7327
rect 23431 7293 23443 7327
rect 23385 7287 23443 7293
rect 25590 7284 25596 7336
rect 25648 7324 25654 7336
rect 26329 7327 26387 7333
rect 26329 7324 26341 7327
rect 25648 7296 26341 7324
rect 25648 7284 25654 7296
rect 26329 7293 26341 7296
rect 26375 7324 26387 7327
rect 26418 7324 26424 7336
rect 26375 7296 26424 7324
rect 26375 7293 26387 7296
rect 26329 7287 26387 7293
rect 26418 7284 26424 7296
rect 26476 7284 26482 7336
rect 26510 7284 26516 7336
rect 26568 7324 26574 7336
rect 26712 7333 26740 7364
rect 27430 7352 27436 7404
rect 27488 7392 27494 7404
rect 27586 7392 27614 7432
rect 27488 7364 27614 7392
rect 28828 7392 28856 7432
rect 30742 7420 30748 7472
rect 30800 7460 30806 7472
rect 31021 7463 31079 7469
rect 31021 7460 31033 7463
rect 30800 7432 31033 7460
rect 30800 7420 30806 7432
rect 31021 7429 31033 7432
rect 31067 7429 31079 7463
rect 31021 7423 31079 7429
rect 31570 7420 31576 7472
rect 31628 7460 31634 7472
rect 39482 7460 39488 7472
rect 31628 7432 32444 7460
rect 31628 7420 31634 7432
rect 32416 7392 32444 7432
rect 36648 7432 39488 7460
rect 32766 7392 32772 7404
rect 28828 7364 29040 7392
rect 32416 7364 32772 7392
rect 27488 7352 27494 7364
rect 26697 7327 26755 7333
rect 26568 7296 26613 7324
rect 26568 7284 26574 7296
rect 26697 7293 26709 7327
rect 26743 7293 26755 7327
rect 26697 7287 26755 7293
rect 27614 7284 27620 7336
rect 27672 7324 27678 7336
rect 28442 7324 28448 7336
rect 27672 7296 28448 7324
rect 27672 7284 27678 7296
rect 28442 7284 28448 7296
rect 28500 7284 28506 7336
rect 28534 7284 28540 7336
rect 28592 7333 28598 7336
rect 28902 7333 28908 7336
rect 28592 7327 28641 7333
rect 28592 7293 28595 7327
rect 28629 7293 28641 7327
rect 28592 7287 28641 7293
rect 28859 7327 28908 7333
rect 28859 7293 28871 7327
rect 28905 7293 28908 7327
rect 28859 7287 28908 7293
rect 28592 7284 28598 7287
rect 28902 7284 28908 7287
rect 28960 7284 28966 7336
rect 22060 7228 23152 7256
rect 22060 7216 22066 7228
rect 23198 7216 23204 7268
rect 23256 7256 23262 7268
rect 24857 7259 24915 7265
rect 23256 7228 23301 7256
rect 23256 7216 23262 7228
rect 24857 7225 24869 7259
rect 24903 7256 24915 7259
rect 26234 7256 26240 7268
rect 24903 7228 26240 7256
rect 24903 7225 24915 7228
rect 24857 7219 24915 7225
rect 26234 7216 26240 7228
rect 26292 7216 26298 7268
rect 26602 7216 26608 7268
rect 26660 7256 26666 7268
rect 28718 7256 28724 7268
rect 26660 7228 26705 7256
rect 28679 7228 28724 7256
rect 26660 7216 26666 7228
rect 28718 7216 28724 7228
rect 28776 7216 28782 7268
rect 20714 7188 20720 7200
rect 19306 7160 20576 7188
rect 20675 7160 20720 7188
rect 19153 7151 19211 7157
rect 20714 7148 20720 7160
rect 20772 7148 20778 7200
rect 22278 7148 22284 7200
rect 22336 7188 22342 7200
rect 23569 7191 23627 7197
rect 23569 7188 23581 7191
rect 22336 7160 23581 7188
rect 22336 7148 22342 7160
rect 23569 7157 23581 7160
rect 23615 7157 23627 7191
rect 24946 7188 24952 7200
rect 24907 7160 24952 7188
rect 23569 7151 23627 7157
rect 24946 7148 24952 7160
rect 25004 7148 25010 7200
rect 25038 7148 25044 7200
rect 25096 7188 25102 7200
rect 29012 7197 29040 7364
rect 32766 7352 32772 7364
rect 32824 7352 32830 7404
rect 33042 7352 33048 7404
rect 33100 7392 33106 7404
rect 33778 7392 33784 7404
rect 33100 7364 33784 7392
rect 33100 7352 33106 7364
rect 29914 7284 29920 7336
rect 29972 7324 29978 7336
rect 30650 7324 30656 7336
rect 29972 7296 30656 7324
rect 29972 7284 29978 7296
rect 30650 7284 30656 7296
rect 30708 7284 30714 7336
rect 30929 7327 30987 7333
rect 30929 7293 30941 7327
rect 30975 7293 30987 7327
rect 30929 7287 30987 7293
rect 31205 7327 31263 7333
rect 31205 7293 31217 7327
rect 31251 7324 31263 7327
rect 31294 7324 31300 7336
rect 31251 7296 31300 7324
rect 31251 7293 31263 7296
rect 31205 7287 31263 7293
rect 29178 7216 29184 7268
rect 29236 7256 29242 7268
rect 29549 7259 29607 7265
rect 29549 7256 29561 7259
rect 29236 7228 29561 7256
rect 29236 7216 29242 7228
rect 29549 7225 29561 7228
rect 29595 7225 29607 7259
rect 30944 7256 30972 7287
rect 31294 7284 31300 7296
rect 31352 7284 31358 7336
rect 33336 7333 33364 7364
rect 33778 7352 33784 7364
rect 33836 7352 33842 7404
rect 33980 7364 34362 7392
rect 33321 7327 33379 7333
rect 33321 7293 33333 7327
rect 33367 7293 33379 7327
rect 33502 7324 33508 7336
rect 33463 7296 33508 7324
rect 33321 7287 33379 7293
rect 33502 7284 33508 7296
rect 33560 7284 33566 7336
rect 33689 7327 33747 7333
rect 33689 7293 33701 7327
rect 33735 7324 33747 7327
rect 33870 7324 33876 7336
rect 33735 7296 33876 7324
rect 33735 7293 33747 7296
rect 33689 7287 33747 7293
rect 33870 7284 33876 7296
rect 33928 7284 33934 7336
rect 31110 7256 31116 7268
rect 30944 7228 31116 7256
rect 29549 7219 29607 7225
rect 31110 7216 31116 7228
rect 31168 7216 31174 7268
rect 33594 7256 33600 7268
rect 33555 7228 33600 7256
rect 33594 7216 33600 7228
rect 33652 7216 33658 7268
rect 33980 7256 34008 7364
rect 34054 7284 34060 7336
rect 34112 7324 34118 7336
rect 34885 7327 34943 7333
rect 34885 7324 34897 7327
rect 34112 7296 34897 7324
rect 34112 7284 34118 7296
rect 34885 7293 34897 7296
rect 34931 7293 34943 7327
rect 35250 7324 35256 7336
rect 35211 7296 35256 7324
rect 34885 7287 34943 7293
rect 35250 7284 35256 7296
rect 35308 7284 35314 7336
rect 36354 7324 36360 7336
rect 36267 7296 36360 7324
rect 36354 7284 36360 7296
rect 36412 7284 36418 7336
rect 36541 7327 36599 7333
rect 36541 7293 36553 7327
rect 36587 7324 36599 7327
rect 36648 7324 36676 7432
rect 39482 7420 39488 7432
rect 39540 7420 39546 7472
rect 43990 7460 43996 7472
rect 40880 7432 43996 7460
rect 40880 7404 40908 7432
rect 43990 7420 43996 7432
rect 44048 7420 44054 7472
rect 44174 7460 44180 7472
rect 44135 7432 44180 7460
rect 44174 7420 44180 7432
rect 44232 7420 44238 7472
rect 46290 7420 46296 7472
rect 46348 7460 46354 7472
rect 46385 7463 46443 7469
rect 46385 7460 46397 7463
rect 46348 7432 46397 7460
rect 46348 7420 46354 7432
rect 46385 7429 46397 7432
rect 46431 7429 46443 7463
rect 46385 7423 46443 7429
rect 46566 7420 46572 7472
rect 46624 7460 46630 7472
rect 46624 7432 49188 7460
rect 46624 7420 46630 7432
rect 37090 7352 37096 7404
rect 37148 7392 37154 7404
rect 37148 7364 38424 7392
rect 37148 7352 37154 7364
rect 36587 7296 36676 7324
rect 36587 7293 36599 7296
rect 36541 7287 36599 7293
rect 36722 7284 36728 7336
rect 36780 7324 36786 7336
rect 38289 7327 38347 7333
rect 36780 7296 36825 7324
rect 36780 7284 36786 7296
rect 38289 7293 38301 7327
rect 38335 7293 38347 7327
rect 38289 7287 38347 7293
rect 34471 7259 34529 7265
rect 34471 7256 34483 7259
rect 33704 7228 34008 7256
rect 34256 7228 34483 7256
rect 26881 7191 26939 7197
rect 26881 7188 26893 7191
rect 25096 7160 26893 7188
rect 25096 7148 25102 7160
rect 26881 7157 26893 7160
rect 26927 7157 26939 7191
rect 26881 7151 26939 7157
rect 28997 7191 29055 7197
rect 28997 7157 29009 7191
rect 29043 7157 29055 7191
rect 28997 7151 29055 7157
rect 29086 7148 29092 7200
rect 29144 7188 29150 7200
rect 29270 7188 29276 7200
rect 29144 7160 29276 7188
rect 29144 7148 29150 7160
rect 29270 7148 29276 7160
rect 29328 7148 29334 7200
rect 29362 7148 29368 7200
rect 29420 7188 29426 7200
rect 30558 7188 30564 7200
rect 29420 7160 30564 7188
rect 29420 7148 29426 7160
rect 30558 7148 30564 7160
rect 30616 7188 30622 7200
rect 31389 7191 31447 7197
rect 31389 7188 31401 7191
rect 30616 7160 31401 7188
rect 30616 7148 30622 7160
rect 31389 7157 31401 7160
rect 31435 7157 31447 7191
rect 31389 7151 31447 7157
rect 33042 7148 33048 7200
rect 33100 7188 33106 7200
rect 33318 7188 33324 7200
rect 33100 7160 33324 7188
rect 33100 7148 33106 7160
rect 33318 7148 33324 7160
rect 33376 7188 33382 7200
rect 33704 7188 33732 7228
rect 34256 7200 34284 7228
rect 34471 7225 34483 7228
rect 34517 7225 34529 7259
rect 34790 7256 34796 7268
rect 34751 7228 34796 7256
rect 34471 7219 34529 7225
rect 34790 7216 34796 7228
rect 34848 7216 34854 7268
rect 33870 7188 33876 7200
rect 33376 7160 33732 7188
rect 33831 7160 33876 7188
rect 33376 7148 33382 7160
rect 33870 7148 33876 7160
rect 33928 7148 33934 7200
rect 34146 7188 34152 7200
rect 34107 7160 34152 7188
rect 34146 7148 34152 7160
rect 34204 7148 34210 7200
rect 34238 7148 34244 7200
rect 34296 7148 34302 7200
rect 35618 7188 35624 7200
rect 35579 7160 35624 7188
rect 35618 7148 35624 7160
rect 35676 7148 35682 7200
rect 36372 7188 36400 7284
rect 36446 7216 36452 7268
rect 36504 7256 36510 7268
rect 36633 7259 36691 7265
rect 36633 7256 36645 7259
rect 36504 7228 36645 7256
rect 36504 7216 36510 7228
rect 36633 7225 36645 7228
rect 36679 7225 36691 7259
rect 38304 7256 38332 7287
rect 36633 7219 36691 7225
rect 36740 7228 38332 7256
rect 38396 7256 38424 7364
rect 38488 7364 39344 7392
rect 38488 7333 38516 7364
rect 38473 7327 38531 7333
rect 38473 7293 38485 7327
rect 38519 7293 38531 7327
rect 38473 7287 38531 7293
rect 38654 7284 38660 7336
rect 38712 7324 38718 7336
rect 38712 7296 38757 7324
rect 38712 7284 38718 7296
rect 38838 7284 38844 7336
rect 38896 7324 38902 7336
rect 39209 7327 39267 7333
rect 39209 7324 39221 7327
rect 38896 7296 39221 7324
rect 38896 7284 38902 7296
rect 39209 7293 39221 7296
rect 39255 7293 39267 7327
rect 39316 7324 39344 7364
rect 39758 7352 39764 7404
rect 39816 7352 39822 7404
rect 40862 7352 40868 7404
rect 40920 7352 40926 7404
rect 41230 7352 41236 7404
rect 41288 7392 41294 7404
rect 41288 7364 42012 7392
rect 41288 7352 41294 7364
rect 41690 7324 41696 7336
rect 39316 7296 40448 7324
rect 41651 7296 41696 7324
rect 39209 7287 39267 7293
rect 38565 7259 38623 7265
rect 38565 7256 38577 7259
rect 38396 7228 38577 7256
rect 36740 7188 36768 7228
rect 38565 7225 38577 7228
rect 38611 7225 38623 7259
rect 38565 7219 38623 7225
rect 36372 7160 36768 7188
rect 36814 7148 36820 7200
rect 36872 7188 36878 7200
rect 36909 7191 36967 7197
rect 36909 7188 36921 7191
rect 36872 7160 36921 7188
rect 36872 7148 36878 7160
rect 36909 7157 36921 7160
rect 36955 7157 36967 7191
rect 36909 7151 36967 7157
rect 37274 7148 37280 7200
rect 37332 7188 37338 7200
rect 38841 7191 38899 7197
rect 38841 7188 38853 7191
rect 37332 7160 38853 7188
rect 37332 7148 37338 7160
rect 38841 7157 38853 7160
rect 38887 7157 38899 7191
rect 39224 7188 39252 7287
rect 39574 7256 39580 7268
rect 39535 7228 39580 7256
rect 39574 7216 39580 7228
rect 39632 7216 39638 7268
rect 39666 7216 39672 7268
rect 39724 7256 39730 7268
rect 39853 7259 39911 7265
rect 39853 7256 39865 7259
rect 39724 7228 39865 7256
rect 39724 7216 39730 7228
rect 39853 7225 39865 7228
rect 39899 7225 39911 7259
rect 39853 7219 39911 7225
rect 39942 7216 39948 7268
rect 40000 7256 40006 7268
rect 40313 7259 40371 7265
rect 40000 7228 40045 7256
rect 40000 7216 40006 7228
rect 40313 7225 40325 7259
rect 40359 7225 40371 7259
rect 40313 7219 40371 7225
rect 39482 7188 39488 7200
rect 39224 7160 39488 7188
rect 38841 7151 38899 7157
rect 39482 7148 39488 7160
rect 39540 7148 39546 7200
rect 39592 7188 39620 7216
rect 40328 7188 40356 7219
rect 39592 7160 40356 7188
rect 40420 7188 40448 7296
rect 41690 7284 41696 7296
rect 41748 7284 41754 7336
rect 41874 7324 41880 7336
rect 41835 7296 41880 7324
rect 41874 7284 41880 7296
rect 41932 7284 41938 7336
rect 41984 7324 42012 7364
rect 42061 7327 42119 7333
rect 42061 7324 42073 7327
rect 41984 7296 42073 7324
rect 42061 7293 42073 7296
rect 42107 7293 42119 7327
rect 42061 7287 42119 7293
rect 42150 7284 42156 7336
rect 42208 7324 42214 7336
rect 43622 7324 43628 7336
rect 42208 7296 42564 7324
rect 43583 7296 43628 7324
rect 42208 7284 42214 7296
rect 40678 7256 40684 7268
rect 40639 7228 40684 7256
rect 40678 7216 40684 7228
rect 40736 7216 40742 7268
rect 40770 7216 40776 7268
rect 40828 7256 40834 7268
rect 41969 7259 42027 7265
rect 41969 7256 41981 7259
rect 40828 7228 41981 7256
rect 40828 7216 40834 7228
rect 41969 7225 41981 7228
rect 42015 7225 42027 7259
rect 42536 7256 42564 7296
rect 43622 7284 43628 7296
rect 43680 7284 43686 7336
rect 43999 7333 44027 7420
rect 44910 7352 44916 7404
rect 44968 7392 44974 7404
rect 45005 7395 45063 7401
rect 45005 7392 45017 7395
rect 44968 7364 45017 7392
rect 44968 7352 44974 7364
rect 45005 7361 45017 7364
rect 45051 7361 45063 7395
rect 48682 7392 48688 7404
rect 45005 7355 45063 7361
rect 46952 7364 48688 7392
rect 43901 7327 43959 7333
rect 43901 7324 43913 7327
rect 43732 7296 43913 7324
rect 43732 7256 43760 7296
rect 43901 7293 43913 7296
rect 43947 7293 43959 7327
rect 43901 7287 43959 7293
rect 43993 7327 44051 7333
rect 43993 7293 44005 7327
rect 44039 7293 44051 7327
rect 43993 7287 44051 7293
rect 45272 7327 45330 7333
rect 45272 7293 45284 7327
rect 45318 7324 45330 7327
rect 46952 7324 46980 7364
rect 48682 7352 48688 7364
rect 48740 7352 48746 7404
rect 49050 7392 49056 7404
rect 48976 7364 49056 7392
rect 45318 7296 46980 7324
rect 47029 7327 47087 7333
rect 45318 7293 45330 7296
rect 45272 7287 45330 7293
rect 47029 7293 47041 7327
rect 47075 7324 47087 7327
rect 47578 7324 47584 7336
rect 47075 7296 47584 7324
rect 47075 7293 47087 7296
rect 47029 7287 47087 7293
rect 47578 7284 47584 7296
rect 47636 7284 47642 7336
rect 48406 7284 48412 7336
rect 48464 7324 48470 7336
rect 48777 7327 48835 7333
rect 48777 7324 48789 7327
rect 48464 7296 48789 7324
rect 48464 7284 48470 7296
rect 48777 7293 48789 7296
rect 48823 7324 48835 7327
rect 48866 7324 48872 7336
rect 48823 7296 48872 7324
rect 48823 7293 48835 7296
rect 48777 7287 48835 7293
rect 48866 7284 48872 7296
rect 48924 7284 48930 7336
rect 48976 7333 49004 7364
rect 49050 7352 49056 7364
rect 49108 7352 49114 7404
rect 49160 7392 49188 7432
rect 49234 7420 49240 7472
rect 49292 7460 49298 7472
rect 54754 7460 54760 7472
rect 49292 7432 54760 7460
rect 49292 7420 49298 7432
rect 54754 7420 54760 7432
rect 54812 7420 54818 7472
rect 56428 7460 56456 7500
rect 56689 7497 56701 7531
rect 56735 7528 56747 7531
rect 57054 7528 57060 7540
rect 56735 7500 57060 7528
rect 56735 7497 56747 7500
rect 56689 7491 56747 7497
rect 57054 7488 57060 7500
rect 57112 7488 57118 7540
rect 59262 7488 59268 7540
rect 59320 7528 59326 7540
rect 60182 7528 60188 7540
rect 59320 7500 60188 7528
rect 59320 7488 59326 7500
rect 60182 7488 60188 7500
rect 60240 7528 60246 7540
rect 61286 7528 61292 7540
rect 60240 7500 61292 7528
rect 60240 7488 60246 7500
rect 61286 7488 61292 7500
rect 61344 7488 61350 7540
rect 61473 7531 61531 7537
rect 61473 7497 61485 7531
rect 61519 7528 61531 7531
rect 63310 7528 63316 7540
rect 61519 7500 63316 7528
rect 61519 7497 61531 7500
rect 61473 7491 61531 7497
rect 63310 7488 63316 7500
rect 63368 7488 63374 7540
rect 64598 7528 64604 7540
rect 64559 7500 64604 7528
rect 64598 7488 64604 7500
rect 64656 7488 64662 7540
rect 59906 7460 59912 7472
rect 54864 7432 55628 7460
rect 56428 7432 59912 7460
rect 54864 7401 54892 7432
rect 54849 7395 54907 7401
rect 49160 7364 51074 7392
rect 48961 7327 49019 7333
rect 48961 7293 48973 7327
rect 49007 7293 49019 7327
rect 49142 7324 49148 7336
rect 49103 7296 49148 7324
rect 48961 7287 49019 7293
rect 49142 7284 49148 7296
rect 49200 7284 49206 7336
rect 49326 7284 49332 7336
rect 49384 7324 49390 7336
rect 49789 7327 49847 7333
rect 49789 7324 49801 7327
rect 49384 7296 49801 7324
rect 49384 7284 49390 7296
rect 49789 7293 49801 7296
rect 49835 7293 49847 7327
rect 49970 7324 49976 7336
rect 49931 7296 49976 7324
rect 49789 7287 49847 7293
rect 49970 7284 49976 7296
rect 50028 7284 50034 7336
rect 50154 7324 50160 7336
rect 50115 7296 50160 7324
rect 50154 7284 50160 7296
rect 50212 7284 50218 7336
rect 51046 7324 51074 7364
rect 54849 7361 54861 7395
rect 54895 7361 54907 7395
rect 54849 7355 54907 7361
rect 55033 7395 55091 7401
rect 55033 7361 55045 7395
rect 55079 7392 55091 7395
rect 55122 7392 55128 7404
rect 55079 7364 55128 7392
rect 55079 7361 55091 7364
rect 55033 7355 55091 7361
rect 55122 7352 55128 7364
rect 55180 7352 55186 7404
rect 55490 7392 55496 7404
rect 55451 7364 55496 7392
rect 55490 7352 55496 7364
rect 55548 7352 55554 7404
rect 55600 7392 55628 7432
rect 59906 7420 59912 7432
rect 59964 7420 59970 7472
rect 55907 7395 55965 7401
rect 55907 7392 55919 7395
rect 55600 7364 55919 7392
rect 55907 7361 55919 7364
rect 55953 7392 55965 7395
rect 56594 7392 56600 7404
rect 55953 7364 56600 7392
rect 55953 7361 55965 7364
rect 55907 7355 55965 7361
rect 56594 7352 56600 7364
rect 56652 7352 56658 7404
rect 62273 7401 62279 7404
rect 62255 7395 62279 7401
rect 62255 7361 62267 7395
rect 62255 7355 62279 7361
rect 62273 7352 62279 7355
rect 62331 7352 62337 7404
rect 62669 7395 62727 7401
rect 62669 7361 62681 7395
rect 62715 7392 62727 7395
rect 62758 7392 62764 7404
rect 62715 7364 62764 7392
rect 62715 7361 62727 7364
rect 62669 7355 62727 7361
rect 62758 7352 62764 7364
rect 62816 7352 62822 7404
rect 63310 7392 63316 7404
rect 63223 7364 63316 7392
rect 63310 7352 63316 7364
rect 63368 7392 63374 7404
rect 64782 7392 64788 7404
rect 63368 7364 64788 7392
rect 63368 7352 63374 7364
rect 64782 7352 64788 7364
rect 64840 7352 64846 7404
rect 65058 7352 65064 7404
rect 65116 7352 65122 7404
rect 55214 7324 55220 7336
rect 51046 7296 55220 7324
rect 55214 7284 55220 7296
rect 55272 7284 55278 7336
rect 55766 7284 55772 7336
rect 55824 7333 55830 7336
rect 55824 7327 55845 7333
rect 55833 7293 55845 7327
rect 56042 7324 56048 7336
rect 56003 7296 56048 7324
rect 55824 7287 55845 7293
rect 55824 7284 55830 7287
rect 56042 7284 56048 7296
rect 56100 7284 56106 7336
rect 56686 7284 56692 7336
rect 56744 7324 56750 7336
rect 61378 7324 61384 7336
rect 56744 7296 61384 7324
rect 56744 7284 56750 7296
rect 61378 7284 61384 7296
rect 61436 7284 61442 7336
rect 62114 7284 62120 7336
rect 62172 7324 62178 7336
rect 62371 7324 62377 7336
rect 62172 7296 62217 7324
rect 62332 7296 62377 7324
rect 62172 7284 62178 7296
rect 62371 7284 62377 7296
rect 62429 7284 62435 7336
rect 63129 7327 63187 7333
rect 63129 7293 63141 7327
rect 63175 7293 63187 7327
rect 86586 7324 86592 7336
rect 63129 7287 63187 7293
rect 63420 7296 86592 7324
rect 41969 7219 42027 7225
rect 42168 7228 42472 7256
rect 42536 7228 43760 7256
rect 43809 7259 43867 7265
rect 42168 7188 42196 7228
rect 40420 7160 42196 7188
rect 42242 7148 42248 7200
rect 42300 7188 42306 7200
rect 42444 7188 42472 7228
rect 43809 7225 43821 7259
rect 43855 7256 43867 7259
rect 47670 7256 47676 7268
rect 43855 7228 47440 7256
rect 47631 7228 47676 7256
rect 43855 7225 43867 7228
rect 43809 7219 43867 7225
rect 46934 7188 46940 7200
rect 42300 7160 42345 7188
rect 42444 7160 46940 7188
rect 42300 7148 42306 7160
rect 46934 7148 46940 7160
rect 46992 7148 46998 7200
rect 47412 7188 47440 7228
rect 47670 7216 47676 7228
rect 47728 7216 47734 7268
rect 48222 7216 48228 7268
rect 48280 7256 48286 7268
rect 49053 7259 49111 7265
rect 49053 7256 49065 7259
rect 48280 7228 49065 7256
rect 48280 7216 48286 7228
rect 49053 7225 49065 7228
rect 49099 7225 49111 7259
rect 49053 7219 49111 7225
rect 49160 7228 49464 7256
rect 49160 7188 49188 7228
rect 49326 7188 49332 7200
rect 47412 7160 49188 7188
rect 49287 7160 49332 7188
rect 49326 7148 49332 7160
rect 49384 7148 49390 7200
rect 49436 7188 49464 7228
rect 49602 7216 49608 7268
rect 49660 7256 49666 7268
rect 50065 7259 50123 7265
rect 50065 7256 50077 7259
rect 49660 7228 50077 7256
rect 49660 7216 49666 7228
rect 50065 7225 50077 7228
rect 50111 7225 50123 7259
rect 50065 7219 50123 7225
rect 50264 7228 51074 7256
rect 50264 7188 50292 7228
rect 49436 7160 50292 7188
rect 50341 7191 50399 7197
rect 50341 7157 50353 7191
rect 50387 7188 50399 7191
rect 50614 7188 50620 7200
rect 50387 7160 50620 7188
rect 50387 7157 50399 7160
rect 50341 7151 50399 7157
rect 50614 7148 50620 7160
rect 50672 7148 50678 7200
rect 51046 7188 51074 7228
rect 56594 7216 56600 7268
rect 56652 7256 56658 7268
rect 61562 7256 61568 7268
rect 56652 7228 61568 7256
rect 56652 7216 56658 7228
rect 61562 7216 61568 7228
rect 61620 7216 61626 7268
rect 63144 7256 63172 7287
rect 63420 7256 63448 7296
rect 86586 7284 86592 7296
rect 86644 7284 86650 7336
rect 63144 7228 63448 7256
rect 65153 7259 65211 7265
rect 61194 7188 61200 7200
rect 51046 7160 61200 7188
rect 61194 7148 61200 7160
rect 61252 7148 61258 7200
rect 61381 7191 61439 7197
rect 61381 7157 61393 7191
rect 61427 7188 61439 7191
rect 63144 7188 63172 7228
rect 65153 7225 65165 7259
rect 65199 7225 65211 7259
rect 65518 7256 65524 7268
rect 65479 7228 65524 7256
rect 65153 7219 65211 7225
rect 61427 7160 63172 7188
rect 64417 7191 64475 7197
rect 61427 7157 61439 7160
rect 61381 7151 61439 7157
rect 64417 7157 64429 7191
rect 64463 7188 64475 7191
rect 64782 7188 64788 7200
rect 64463 7160 64788 7188
rect 64463 7157 64475 7160
rect 64417 7151 64475 7157
rect 64782 7148 64788 7160
rect 64840 7148 64846 7200
rect 65168 7188 65196 7219
rect 65518 7216 65524 7228
rect 65576 7216 65582 7268
rect 65613 7259 65671 7265
rect 65613 7225 65625 7259
rect 65659 7256 65671 7259
rect 66070 7256 66076 7268
rect 65659 7228 66076 7256
rect 65659 7225 65671 7228
rect 65613 7219 65671 7225
rect 66070 7216 66076 7228
rect 66128 7216 66134 7268
rect 66254 7216 66260 7268
rect 66312 7256 66318 7268
rect 68094 7256 68100 7268
rect 66312 7228 68100 7256
rect 66312 7216 66318 7228
rect 68094 7216 68100 7228
rect 68152 7216 68158 7268
rect 65889 7191 65947 7197
rect 65889 7188 65901 7191
rect 65168 7160 65901 7188
rect 65889 7157 65901 7160
rect 65935 7188 65947 7191
rect 68278 7188 68284 7200
rect 65935 7160 68284 7188
rect 65935 7157 65947 7160
rect 65889 7151 65947 7157
rect 68278 7148 68284 7160
rect 68336 7148 68342 7200
rect 1104 7098 178848 7120
rect 1104 7046 19606 7098
rect 19658 7046 19670 7098
rect 19722 7046 19734 7098
rect 19786 7046 19798 7098
rect 19850 7046 50326 7098
rect 50378 7046 50390 7098
rect 50442 7046 50454 7098
rect 50506 7046 50518 7098
rect 50570 7046 81046 7098
rect 81098 7046 81110 7098
rect 81162 7046 81174 7098
rect 81226 7046 81238 7098
rect 81290 7046 111766 7098
rect 111818 7046 111830 7098
rect 111882 7046 111894 7098
rect 111946 7046 111958 7098
rect 112010 7046 142486 7098
rect 142538 7046 142550 7098
rect 142602 7046 142614 7098
rect 142666 7046 142678 7098
rect 142730 7046 173206 7098
rect 173258 7046 173270 7098
rect 173322 7046 173334 7098
rect 173386 7046 173398 7098
rect 173450 7046 178848 7098
rect 1104 7024 178848 7046
rect 21082 6944 21088 6996
rect 21140 6984 21146 6996
rect 21140 6956 21185 6984
rect 21376 6956 21980 6984
rect 21140 6944 21146 6956
rect 18598 6916 18604 6928
rect 18511 6888 18604 6916
rect 16660 6851 16718 6857
rect 16660 6817 16672 6851
rect 16706 6848 16718 6851
rect 17954 6848 17960 6860
rect 16706 6820 17960 6848
rect 16706 6817 16718 6820
rect 16660 6811 16718 6817
rect 17954 6808 17960 6820
rect 18012 6808 18018 6860
rect 18524 6857 18552 6888
rect 18598 6876 18604 6888
rect 18656 6916 18662 6928
rect 18656 6888 19334 6916
rect 18656 6876 18662 6888
rect 18509 6851 18567 6857
rect 18509 6817 18521 6851
rect 18555 6817 18567 6851
rect 18690 6848 18696 6860
rect 18651 6820 18696 6848
rect 18509 6811 18567 6817
rect 18690 6808 18696 6820
rect 18748 6808 18754 6860
rect 18785 6851 18843 6857
rect 18785 6817 18797 6851
rect 18831 6817 18843 6851
rect 18785 6811 18843 6817
rect 18877 6851 18935 6857
rect 18877 6817 18889 6851
rect 18923 6848 18935 6851
rect 18966 6848 18972 6860
rect 18923 6820 18972 6848
rect 18923 6817 18935 6820
rect 18877 6811 18935 6817
rect 16393 6783 16451 6789
rect 16393 6749 16405 6783
rect 16439 6749 16451 6783
rect 16393 6743 16451 6749
rect 16408 6644 16436 6743
rect 18598 6740 18604 6792
rect 18656 6780 18662 6792
rect 18800 6780 18828 6811
rect 18966 6808 18972 6820
rect 19024 6808 19030 6860
rect 19306 6848 19334 6888
rect 20162 6848 20168 6860
rect 19306 6820 20168 6848
rect 20162 6808 20168 6820
rect 20220 6848 20226 6860
rect 20530 6848 20536 6860
rect 20220 6820 20536 6848
rect 20220 6808 20226 6820
rect 20530 6808 20536 6820
rect 20588 6808 20594 6860
rect 20622 6808 20628 6860
rect 20680 6848 20686 6860
rect 20717 6851 20775 6857
rect 20717 6848 20729 6851
rect 20680 6820 20729 6848
rect 20680 6808 20686 6820
rect 20717 6817 20729 6820
rect 20763 6817 20775 6851
rect 20717 6811 20775 6817
rect 20809 6851 20867 6857
rect 20809 6817 20821 6851
rect 20855 6817 20867 6851
rect 20809 6811 20867 6817
rect 18656 6752 18828 6780
rect 18656 6740 18662 6752
rect 17402 6672 17408 6724
rect 17460 6712 17466 6724
rect 17460 6684 19196 6712
rect 17460 6672 17466 6684
rect 17310 6644 17316 6656
rect 16408 6616 17316 6644
rect 17310 6604 17316 6616
rect 17368 6604 17374 6656
rect 17773 6647 17831 6653
rect 17773 6613 17785 6647
rect 17819 6644 17831 6647
rect 17954 6644 17960 6656
rect 17819 6616 17960 6644
rect 17819 6613 17831 6616
rect 17773 6607 17831 6613
rect 17954 6604 17960 6616
rect 18012 6604 18018 6656
rect 18046 6604 18052 6656
rect 18104 6644 18110 6656
rect 19061 6647 19119 6653
rect 19061 6644 19073 6647
rect 18104 6616 19073 6644
rect 18104 6604 18110 6616
rect 19061 6613 19073 6616
rect 19107 6613 19119 6647
rect 19168 6644 19196 6684
rect 20530 6672 20536 6724
rect 20588 6712 20594 6724
rect 20824 6712 20852 6811
rect 20898 6808 20904 6860
rect 20956 6848 20962 6860
rect 21376 6848 21404 6956
rect 21726 6916 21732 6928
rect 21687 6888 21732 6916
rect 21726 6876 21732 6888
rect 21784 6876 21790 6928
rect 21952 6916 21980 6956
rect 23198 6944 23204 6996
rect 23256 6984 23262 6996
rect 33318 6984 33324 6996
rect 23256 6956 33324 6984
rect 23256 6944 23262 6956
rect 33318 6944 33324 6956
rect 33376 6944 33382 6996
rect 33502 6944 33508 6996
rect 33560 6984 33566 6996
rect 40954 6984 40960 6996
rect 33560 6956 40960 6984
rect 33560 6944 33566 6956
rect 40954 6944 40960 6956
rect 41012 6944 41018 6996
rect 41138 6984 41144 6996
rect 41099 6956 41144 6984
rect 41138 6944 41144 6956
rect 41196 6944 41202 6996
rect 41230 6944 41236 6996
rect 41288 6984 41294 6996
rect 41288 6956 41460 6984
rect 41288 6944 41294 6956
rect 24946 6916 24952 6928
rect 21952 6888 24952 6916
rect 21542 6848 21548 6860
rect 20956 6820 21404 6848
rect 21503 6820 21548 6848
rect 20956 6808 20962 6820
rect 21542 6808 21548 6820
rect 21600 6808 21606 6860
rect 21952 6857 21980 6888
rect 24946 6876 24952 6888
rect 25004 6876 25010 6928
rect 29178 6916 29184 6928
rect 28828 6888 29184 6916
rect 21817 6851 21875 6857
rect 21817 6817 21829 6851
rect 21863 6817 21875 6851
rect 21817 6811 21875 6817
rect 21937 6851 21995 6857
rect 21937 6817 21949 6851
rect 21983 6817 21995 6851
rect 21937 6811 21995 6817
rect 25501 6851 25559 6857
rect 25501 6817 25513 6851
rect 25547 6848 25559 6851
rect 28537 6851 28595 6857
rect 28537 6848 28549 6851
rect 25547 6820 28549 6848
rect 25547 6817 25559 6820
rect 25501 6811 25559 6817
rect 28537 6817 28549 6820
rect 28583 6848 28595 6851
rect 28828 6848 28856 6888
rect 29178 6876 29184 6888
rect 29236 6876 29242 6928
rect 29288 6888 30972 6916
rect 28583 6820 28856 6848
rect 28583 6817 28595 6820
rect 28537 6811 28595 6817
rect 21836 6780 21864 6811
rect 28902 6808 28908 6860
rect 28960 6848 28966 6860
rect 29288 6848 29316 6888
rect 28960 6820 29316 6848
rect 28960 6808 28966 6820
rect 29362 6808 29368 6860
rect 29420 6848 29426 6860
rect 30558 6848 30564 6860
rect 29420 6820 29465 6848
rect 30519 6820 30564 6848
rect 29420 6808 29426 6820
rect 30558 6808 30564 6820
rect 30616 6808 30622 6860
rect 30944 6848 30972 6888
rect 31018 6876 31024 6928
rect 31076 6916 31082 6928
rect 31202 6916 31208 6928
rect 31076 6888 31208 6916
rect 31076 6876 31082 6888
rect 31202 6876 31208 6888
rect 31260 6876 31266 6928
rect 31389 6919 31447 6925
rect 31389 6885 31401 6919
rect 31435 6885 31447 6919
rect 31389 6879 31447 6885
rect 31404 6848 31432 6879
rect 31478 6876 31484 6928
rect 31536 6916 31542 6928
rect 31644 6919 31702 6925
rect 31644 6916 31656 6919
rect 31536 6888 31656 6916
rect 31536 6876 31542 6888
rect 31644 6885 31656 6888
rect 31690 6885 31702 6919
rect 31644 6879 31702 6885
rect 31754 6876 31760 6928
rect 31812 6916 31818 6928
rect 32493 6919 32551 6925
rect 31812 6888 31857 6916
rect 31812 6876 31818 6888
rect 32493 6885 32505 6919
rect 32539 6885 32551 6919
rect 32493 6879 32551 6885
rect 33413 6919 33471 6925
rect 33413 6885 33425 6919
rect 33459 6916 33471 6919
rect 34517 6919 34575 6925
rect 33459 6888 34192 6916
rect 33459 6885 33471 6888
rect 33413 6879 33471 6885
rect 32125 6851 32183 6857
rect 32125 6848 32137 6851
rect 30944 6820 32137 6848
rect 32125 6817 32137 6820
rect 32171 6817 32183 6851
rect 32508 6848 32536 6879
rect 32950 6848 32956 6860
rect 32508 6820 32956 6848
rect 32125 6811 32183 6817
rect 32950 6808 32956 6820
rect 33008 6808 33014 6860
rect 33134 6808 33140 6860
rect 33192 6848 33198 6860
rect 33428 6848 33456 6879
rect 33192 6820 33456 6848
rect 33192 6808 33198 6820
rect 33502 6808 33508 6860
rect 33560 6848 33566 6860
rect 33689 6851 33747 6857
rect 33689 6848 33701 6851
rect 33560 6820 33701 6848
rect 33560 6808 33566 6820
rect 33689 6817 33701 6820
rect 33735 6817 33747 6851
rect 33689 6811 33747 6817
rect 33778 6808 33784 6860
rect 33836 6848 33842 6860
rect 34054 6848 34060 6860
rect 33836 6820 34060 6848
rect 33836 6808 33842 6820
rect 34054 6808 34060 6820
rect 34112 6808 34118 6860
rect 34164 6857 34192 6888
rect 34517 6885 34529 6919
rect 34563 6885 34575 6919
rect 34517 6879 34575 6885
rect 34149 6851 34207 6857
rect 34149 6817 34161 6851
rect 34195 6817 34207 6851
rect 34532 6848 34560 6879
rect 34790 6876 34796 6928
rect 34848 6916 34854 6928
rect 36814 6916 36820 6928
rect 34848 6888 36820 6916
rect 34848 6876 34854 6888
rect 36814 6876 36820 6888
rect 36872 6876 36878 6928
rect 39761 6919 39819 6925
rect 39761 6885 39773 6919
rect 39807 6916 39819 6919
rect 40034 6916 40040 6928
rect 39807 6888 40040 6916
rect 39807 6885 39819 6888
rect 39761 6879 39819 6885
rect 40034 6876 40040 6888
rect 40092 6876 40098 6928
rect 35986 6848 35992 6860
rect 34532 6820 35296 6848
rect 35947 6820 35992 6848
rect 34149 6811 34207 6817
rect 30282 6780 30288 6792
rect 20588 6684 20852 6712
rect 20907 6752 21864 6780
rect 22020 6752 30288 6780
rect 20588 6672 20594 6684
rect 20907 6644 20935 6752
rect 21726 6672 21732 6724
rect 21784 6712 21790 6724
rect 22020 6712 22048 6752
rect 30282 6740 30288 6752
rect 30340 6740 30346 6792
rect 31018 6740 31024 6792
rect 31076 6780 31082 6792
rect 35268 6780 35296 6820
rect 35986 6808 35992 6820
rect 36044 6808 36050 6860
rect 36630 6848 36636 6860
rect 36591 6820 36636 6848
rect 36630 6808 36636 6820
rect 36688 6808 36694 6860
rect 37642 6808 37648 6860
rect 37700 6857 37706 6860
rect 37700 6851 37728 6857
rect 37716 6817 37728 6851
rect 37700 6811 37728 6817
rect 37700 6808 37706 6811
rect 38562 6808 38568 6860
rect 38620 6848 38626 6860
rect 41432 6857 41460 6956
rect 41874 6944 41880 6996
rect 41932 6984 41938 6996
rect 56594 6984 56600 6996
rect 41932 6956 56600 6984
rect 41932 6944 41938 6956
rect 56594 6944 56600 6956
rect 56652 6944 56658 6996
rect 62022 6984 62028 6996
rect 56704 6956 62028 6984
rect 42245 6919 42303 6925
rect 42245 6885 42257 6919
rect 42291 6916 42303 6919
rect 46753 6919 46811 6925
rect 42291 6888 42380 6916
rect 42291 6885 42303 6888
rect 42245 6879 42303 6885
rect 39577 6851 39635 6857
rect 39577 6848 39589 6851
rect 38620 6820 39589 6848
rect 38620 6808 38626 6820
rect 39577 6817 39589 6820
rect 39623 6817 39635 6851
rect 39577 6811 39635 6817
rect 41417 6851 41475 6857
rect 41417 6817 41429 6851
rect 41463 6817 41475 6851
rect 41417 6811 41475 6817
rect 41509 6851 41567 6857
rect 41509 6817 41521 6851
rect 41555 6848 41567 6851
rect 41690 6848 41696 6860
rect 41555 6820 41696 6848
rect 41555 6817 41567 6820
rect 41509 6811 41567 6817
rect 41690 6808 41696 6820
rect 41748 6808 41754 6860
rect 41874 6848 41880 6860
rect 41835 6820 41880 6848
rect 41874 6808 41880 6820
rect 41932 6808 41938 6860
rect 42352 6848 42380 6888
rect 46753 6885 46765 6919
rect 46799 6885 46811 6919
rect 46753 6879 46811 6885
rect 43530 6848 43536 6860
rect 42352 6820 43536 6848
rect 43530 6808 43536 6820
rect 43588 6808 43594 6860
rect 44450 6808 44456 6860
rect 44508 6857 44514 6860
rect 44508 6851 44536 6857
rect 44524 6817 44536 6851
rect 44634 6848 44640 6860
rect 44595 6820 44640 6848
rect 44508 6811 44536 6817
rect 44508 6808 44514 6811
rect 44634 6808 44640 6820
rect 44692 6808 44698 6860
rect 45278 6848 45284 6860
rect 45239 6820 45284 6848
rect 45278 6808 45284 6820
rect 45336 6808 45342 6860
rect 46382 6808 46388 6860
rect 46440 6848 46446 6860
rect 46477 6851 46535 6857
rect 46477 6848 46489 6851
rect 46440 6820 46489 6848
rect 46440 6808 46446 6820
rect 46477 6817 46489 6820
rect 46523 6817 46535 6851
rect 46658 6848 46664 6860
rect 46619 6820 46664 6848
rect 46477 6811 46535 6817
rect 46658 6808 46664 6820
rect 46716 6808 46722 6860
rect 31076 6752 31234 6780
rect 31076 6740 31082 6752
rect 21784 6684 22048 6712
rect 21784 6672 21790 6684
rect 22094 6672 22100 6724
rect 22152 6712 22158 6724
rect 22152 6684 22197 6712
rect 22152 6672 22158 6684
rect 23014 6672 23020 6724
rect 23072 6712 23078 6724
rect 25685 6715 25743 6721
rect 25685 6712 25697 6715
rect 23072 6684 25697 6712
rect 23072 6672 23078 6684
rect 25685 6681 25697 6684
rect 25731 6681 25743 6715
rect 31294 6712 31300 6724
rect 25685 6675 25743 6681
rect 28184 6684 29592 6712
rect 19168 6616 20935 6644
rect 19061 6607 19119 6613
rect 21174 6604 21180 6656
rect 21232 6644 21238 6656
rect 28184 6644 28212 6684
rect 21232 6616 28212 6644
rect 21232 6604 21238 6616
rect 28534 6604 28540 6656
rect 28592 6644 28598 6656
rect 28629 6647 28687 6653
rect 28629 6644 28641 6647
rect 28592 6616 28641 6644
rect 28592 6604 28598 6616
rect 28629 6613 28641 6616
rect 28675 6613 28687 6647
rect 28629 6607 28687 6613
rect 29178 6604 29184 6656
rect 29236 6644 29242 6656
rect 29457 6647 29515 6653
rect 29457 6644 29469 6647
rect 29236 6616 29469 6644
rect 29236 6604 29242 6616
rect 29457 6613 29469 6616
rect 29503 6613 29515 6647
rect 29564 6644 29592 6684
rect 30668 6684 31300 6712
rect 30668 6653 30696 6684
rect 31294 6672 31300 6684
rect 31352 6672 31358 6724
rect 32674 6712 32680 6724
rect 32635 6684 32680 6712
rect 32674 6672 32680 6684
rect 32732 6672 32738 6724
rect 33134 6672 33140 6724
rect 33192 6712 33198 6724
rect 33244 6712 33272 6766
rect 35268 6752 36676 6780
rect 33192 6684 33272 6712
rect 34701 6715 34759 6721
rect 33192 6672 33198 6684
rect 34701 6681 34713 6715
rect 34747 6712 34759 6715
rect 34882 6712 34888 6724
rect 34747 6684 34888 6712
rect 34747 6681 34759 6684
rect 34701 6675 34759 6681
rect 34882 6672 34888 6684
rect 34940 6672 34946 6724
rect 36173 6715 36231 6721
rect 36173 6681 36185 6715
rect 36219 6712 36231 6715
rect 36538 6712 36544 6724
rect 36219 6684 36544 6712
rect 36219 6681 36231 6684
rect 36173 6675 36231 6681
rect 36538 6672 36544 6684
rect 36596 6672 36602 6724
rect 36648 6712 36676 6752
rect 36722 6740 36728 6792
rect 36780 6780 36786 6792
rect 36817 6783 36875 6789
rect 36817 6780 36829 6783
rect 36780 6752 36829 6780
rect 36780 6740 36786 6752
rect 36817 6749 36829 6752
rect 36863 6749 36875 6783
rect 36817 6743 36875 6749
rect 36906 6740 36912 6792
rect 36964 6780 36970 6792
rect 36964 6752 37136 6780
rect 36964 6740 36970 6752
rect 37108 6712 37136 6752
rect 37182 6740 37188 6792
rect 37240 6780 37246 6792
rect 37277 6783 37335 6789
rect 37277 6780 37289 6783
rect 37240 6752 37289 6780
rect 37240 6740 37246 6752
rect 37277 6749 37289 6752
rect 37323 6749 37335 6783
rect 37553 6783 37611 6789
rect 37553 6780 37565 6783
rect 37277 6743 37335 6749
rect 37384 6752 37565 6780
rect 37384 6712 37412 6752
rect 37553 6749 37565 6752
rect 37599 6749 37611 6783
rect 37826 6780 37832 6792
rect 37787 6752 37832 6780
rect 37553 6743 37611 6749
rect 37826 6740 37832 6752
rect 37884 6740 37890 6792
rect 38378 6740 38384 6792
rect 38436 6780 38442 6792
rect 38473 6783 38531 6789
rect 38473 6780 38485 6783
rect 38436 6752 38485 6780
rect 38436 6740 38442 6752
rect 38473 6749 38485 6752
rect 38519 6749 38531 6783
rect 38473 6743 38531 6749
rect 39758 6740 39764 6792
rect 39816 6780 39822 6792
rect 40862 6780 40868 6792
rect 39816 6752 40868 6780
rect 39816 6740 39822 6752
rect 40862 6740 40868 6752
rect 40920 6780 40926 6792
rect 43349 6783 43407 6789
rect 40920 6752 40986 6780
rect 40920 6740 40926 6752
rect 43349 6749 43361 6783
rect 43395 6780 43407 6783
rect 43441 6783 43499 6789
rect 43441 6780 43453 6783
rect 43395 6752 43453 6780
rect 43395 6749 43407 6752
rect 43349 6743 43407 6749
rect 43441 6749 43453 6752
rect 43487 6749 43499 6783
rect 43622 6780 43628 6792
rect 43583 6752 43628 6780
rect 43441 6743 43499 6749
rect 43622 6740 43628 6752
rect 43680 6740 43686 6792
rect 44358 6740 44364 6792
rect 44416 6780 44422 6792
rect 44416 6752 44461 6780
rect 44416 6740 44422 6752
rect 42426 6712 42432 6724
rect 36648 6684 37044 6712
rect 37108 6684 37412 6712
rect 42387 6684 42432 6712
rect 30653 6647 30711 6653
rect 30653 6644 30665 6647
rect 29564 6616 30665 6644
rect 29457 6607 29515 6613
rect 30653 6613 30665 6616
rect 30699 6613 30711 6647
rect 30653 6607 30711 6613
rect 30834 6604 30840 6656
rect 30892 6644 30898 6656
rect 31021 6647 31079 6653
rect 31021 6644 31033 6647
rect 30892 6616 31033 6644
rect 30892 6604 30898 6616
rect 31021 6613 31033 6616
rect 31067 6644 31079 6647
rect 31386 6644 31392 6656
rect 31067 6616 31392 6644
rect 31067 6613 31079 6616
rect 31021 6607 31079 6613
rect 31386 6604 31392 6616
rect 31444 6604 31450 6656
rect 35894 6604 35900 6656
rect 35952 6644 35958 6656
rect 36449 6647 36507 6653
rect 36449 6644 36461 6647
rect 35952 6616 36461 6644
rect 35952 6604 35958 6616
rect 36449 6613 36461 6616
rect 36495 6644 36507 6647
rect 36814 6644 36820 6656
rect 36495 6616 36820 6644
rect 36495 6613 36507 6616
rect 36449 6607 36507 6613
rect 36814 6604 36820 6616
rect 36872 6604 36878 6656
rect 37016 6644 37044 6684
rect 42426 6672 42432 6684
rect 42484 6672 42490 6724
rect 44082 6712 44088 6724
rect 44043 6684 44088 6712
rect 44082 6672 44088 6684
rect 44140 6672 44146 6724
rect 45370 6672 45376 6724
rect 45428 6712 45434 6724
rect 46768 6712 46796 6879
rect 49970 6876 49976 6928
rect 50028 6916 50034 6928
rect 50157 6919 50215 6925
rect 50157 6916 50169 6919
rect 50028 6888 50169 6916
rect 50028 6876 50034 6888
rect 50157 6885 50169 6888
rect 50203 6885 50215 6919
rect 50157 6879 50215 6885
rect 55674 6876 55680 6928
rect 55732 6916 55738 6928
rect 56704 6916 56732 6956
rect 62022 6944 62028 6956
rect 62080 6944 62086 6996
rect 62574 6944 62580 6996
rect 62632 6984 62638 6996
rect 63497 6987 63555 6993
rect 63497 6984 63509 6987
rect 62632 6956 63509 6984
rect 62632 6944 62638 6956
rect 63497 6953 63509 6956
rect 63543 6984 63555 6987
rect 64598 6984 64604 6996
rect 63543 6956 64604 6984
rect 63543 6953 63555 6956
rect 63497 6947 63555 6953
rect 64598 6944 64604 6956
rect 64656 6944 64662 6996
rect 64782 6944 64788 6996
rect 64840 6984 64846 6996
rect 84838 6984 84844 6996
rect 64840 6956 84844 6984
rect 64840 6944 64846 6956
rect 84838 6944 84844 6956
rect 84896 6944 84902 6996
rect 55732 6888 56732 6916
rect 55732 6876 55738 6888
rect 59906 6876 59912 6928
rect 59964 6916 59970 6928
rect 61102 6916 61108 6928
rect 59964 6888 61108 6916
rect 59964 6876 59970 6888
rect 61102 6876 61108 6888
rect 61160 6876 61166 6928
rect 61378 6876 61384 6928
rect 61436 6916 61442 6928
rect 63586 6916 63592 6928
rect 61436 6888 62528 6916
rect 61436 6876 61442 6888
rect 62500 6860 62528 6888
rect 63512 6888 63592 6916
rect 46842 6808 46848 6860
rect 46900 6848 46906 6860
rect 46900 6820 46945 6848
rect 46900 6808 46906 6820
rect 47210 6808 47216 6860
rect 47268 6848 47274 6860
rect 47268 6820 47716 6848
rect 47268 6808 47274 6820
rect 47118 6780 47124 6792
rect 45428 6684 46796 6712
rect 47044 6752 47124 6780
rect 45428 6672 45434 6684
rect 41138 6644 41144 6656
rect 37016 6616 41144 6644
rect 41138 6604 41144 6616
rect 41196 6604 41202 6656
rect 43349 6647 43407 6653
rect 43349 6613 43361 6647
rect 43395 6644 43407 6647
rect 44450 6644 44456 6656
rect 43395 6616 44456 6644
rect 43395 6613 43407 6616
rect 43349 6607 43407 6613
rect 44450 6604 44456 6616
rect 44508 6604 44514 6656
rect 47044 6653 47072 6752
rect 47118 6740 47124 6752
rect 47176 6740 47182 6792
rect 47581 6783 47639 6789
rect 47581 6749 47593 6783
rect 47627 6749 47639 6783
rect 47581 6743 47639 6749
rect 47029 6647 47087 6653
rect 47029 6613 47041 6647
rect 47075 6613 47087 6647
rect 47596 6644 47624 6743
rect 47688 6712 47716 6820
rect 48590 6808 48596 6860
rect 48648 6857 48654 6860
rect 48648 6851 48676 6857
rect 48664 6817 48676 6851
rect 49418 6848 49424 6860
rect 49379 6820 49424 6848
rect 48648 6811 48676 6817
rect 48648 6808 48654 6811
rect 49418 6808 49424 6820
rect 49476 6808 49482 6860
rect 49881 6851 49939 6857
rect 49881 6817 49893 6851
rect 49927 6817 49939 6851
rect 49881 6811 49939 6817
rect 47765 6783 47823 6789
rect 47765 6749 47777 6783
rect 47811 6780 47823 6783
rect 47946 6780 47952 6792
rect 47811 6752 47952 6780
rect 47811 6749 47823 6752
rect 47765 6743 47823 6749
rect 47946 6740 47952 6752
rect 48004 6740 48010 6792
rect 48498 6780 48504 6792
rect 48459 6752 48504 6780
rect 48498 6740 48504 6752
rect 48556 6740 48562 6792
rect 48774 6780 48780 6792
rect 48735 6752 48780 6780
rect 48774 6740 48780 6752
rect 48832 6740 48838 6792
rect 48958 6740 48964 6792
rect 49016 6780 49022 6792
rect 49896 6780 49924 6811
rect 50062 6808 50068 6860
rect 50120 6848 50126 6860
rect 50246 6848 50252 6860
rect 50120 6820 50165 6848
rect 50207 6820 50252 6848
rect 50120 6808 50126 6820
rect 50246 6808 50252 6820
rect 50304 6808 50310 6860
rect 52822 6848 52828 6860
rect 52783 6820 52828 6848
rect 52822 6808 52828 6820
rect 52880 6808 52886 6860
rect 53466 6848 53472 6860
rect 53427 6820 53472 6848
rect 53466 6808 53472 6820
rect 53524 6808 53530 6860
rect 53576 6820 54248 6848
rect 49016 6752 49924 6780
rect 51629 6783 51687 6789
rect 49016 6740 49022 6752
rect 51629 6749 51641 6783
rect 51675 6749 51687 6783
rect 51810 6780 51816 6792
rect 51771 6752 51816 6780
rect 51629 6743 51687 6749
rect 48225 6715 48283 6721
rect 48225 6712 48237 6715
rect 47688 6684 48237 6712
rect 48225 6681 48237 6684
rect 48271 6681 48283 6715
rect 48225 6675 48283 6681
rect 48590 6644 48596 6656
rect 47596 6616 48596 6644
rect 47029 6607 47087 6613
rect 48590 6604 48596 6616
rect 48648 6604 48654 6656
rect 49510 6604 49516 6656
rect 49568 6644 49574 6656
rect 50433 6647 50491 6653
rect 50433 6644 50445 6647
rect 49568 6616 50445 6644
rect 49568 6604 49574 6616
rect 50433 6613 50445 6616
rect 50479 6613 50491 6647
rect 51644 6644 51672 6743
rect 51810 6740 51816 6752
rect 51868 6740 51874 6792
rect 52546 6740 52552 6792
rect 52604 6780 52610 6792
rect 52687 6783 52745 6789
rect 52604 6752 52649 6780
rect 52604 6740 52610 6752
rect 52687 6749 52699 6783
rect 52733 6780 52745 6783
rect 53576 6780 53604 6820
rect 52733 6752 53604 6780
rect 53929 6783 53987 6789
rect 52733 6749 52745 6752
rect 52687 6743 52745 6749
rect 52178 6672 52184 6724
rect 52236 6712 52242 6724
rect 52273 6715 52331 6721
rect 52273 6712 52285 6715
rect 52236 6684 52285 6712
rect 52236 6672 52242 6684
rect 52273 6681 52285 6684
rect 52319 6681 52331 6715
rect 52273 6675 52331 6681
rect 53208 6644 53236 6752
rect 53929 6749 53941 6783
rect 53975 6749 53987 6783
rect 53929 6743 53987 6749
rect 51644 6616 53236 6644
rect 53944 6644 53972 6743
rect 54018 6740 54024 6792
rect 54076 6780 54082 6792
rect 54113 6783 54171 6789
rect 54113 6780 54125 6783
rect 54076 6752 54125 6780
rect 54076 6740 54082 6752
rect 54113 6749 54125 6752
rect 54159 6749 54171 6783
rect 54220 6780 54248 6820
rect 54938 6808 54944 6860
rect 54996 6857 55002 6860
rect 54996 6851 55024 6857
rect 55012 6817 55024 6851
rect 54996 6811 55024 6817
rect 55769 6851 55827 6857
rect 55769 6817 55781 6851
rect 55815 6848 55827 6851
rect 56226 6848 56232 6860
rect 55815 6820 56232 6848
rect 55815 6817 55827 6820
rect 55769 6811 55827 6817
rect 54996 6808 55002 6811
rect 56226 6808 56232 6820
rect 56284 6808 56290 6860
rect 56870 6808 56876 6860
rect 56928 6848 56934 6860
rect 57057 6851 57115 6857
rect 57057 6848 57069 6851
rect 56928 6820 57069 6848
rect 56928 6808 56934 6820
rect 57057 6817 57069 6820
rect 57103 6817 57115 6851
rect 59170 6848 59176 6860
rect 59131 6820 59176 6848
rect 57057 6811 57115 6817
rect 59170 6808 59176 6820
rect 59228 6808 59234 6860
rect 59998 6848 60004 6860
rect 59740 6820 60004 6848
rect 54662 6780 54668 6792
rect 54220 6752 54668 6780
rect 54113 6743 54171 6749
rect 54662 6740 54668 6752
rect 54720 6740 54726 6792
rect 54846 6780 54852 6792
rect 54807 6752 54852 6780
rect 54846 6740 54852 6752
rect 54904 6740 54910 6792
rect 55125 6783 55183 6789
rect 55125 6749 55137 6783
rect 55171 6780 55183 6783
rect 55306 6780 55312 6792
rect 55171 6752 55312 6780
rect 55171 6749 55183 6752
rect 55125 6743 55183 6749
rect 55306 6740 55312 6752
rect 55364 6740 55370 6792
rect 58342 6780 58348 6792
rect 55784 6752 58348 6780
rect 54570 6712 54576 6724
rect 54531 6684 54576 6712
rect 54570 6672 54576 6684
rect 54628 6672 54634 6724
rect 54938 6644 54944 6656
rect 53944 6616 54944 6644
rect 50433 6607 50491 6613
rect 54938 6604 54944 6616
rect 54996 6604 55002 6656
rect 55122 6604 55128 6656
rect 55180 6644 55186 6656
rect 55784 6644 55812 6752
rect 58342 6740 58348 6752
rect 58400 6740 58406 6792
rect 58710 6780 58716 6792
rect 58544 6752 58716 6780
rect 56042 6672 56048 6724
rect 56100 6712 56106 6724
rect 57330 6712 57336 6724
rect 56100 6684 57336 6712
rect 56100 6672 56106 6684
rect 57330 6672 57336 6684
rect 57388 6712 57394 6724
rect 58544 6712 58572 6752
rect 58710 6740 58716 6752
rect 58768 6780 58774 6792
rect 58897 6783 58955 6789
rect 58897 6780 58909 6783
rect 58768 6752 58909 6780
rect 58768 6740 58774 6752
rect 58897 6749 58909 6752
rect 58943 6749 58955 6783
rect 58897 6743 58955 6749
rect 59035 6783 59093 6789
rect 59035 6749 59047 6783
rect 59081 6780 59093 6783
rect 59740 6780 59768 6820
rect 59998 6808 60004 6820
rect 60056 6848 60062 6860
rect 60093 6851 60151 6857
rect 60093 6848 60105 6851
rect 60056 6820 60105 6848
rect 60056 6808 60062 6820
rect 60093 6817 60105 6820
rect 60139 6817 60151 6851
rect 60093 6811 60151 6817
rect 61654 6808 61660 6860
rect 61712 6848 61718 6860
rect 62117 6851 62175 6857
rect 62117 6848 62129 6851
rect 61712 6820 62129 6848
rect 61712 6808 61718 6820
rect 62117 6817 62129 6820
rect 62163 6817 62175 6851
rect 62117 6811 62175 6817
rect 62482 6808 62488 6860
rect 62540 6848 62546 6860
rect 62945 6851 63003 6857
rect 62945 6848 62957 6851
rect 62540 6820 62957 6848
rect 62540 6808 62546 6820
rect 62945 6817 62957 6820
rect 62991 6817 63003 6851
rect 62945 6811 63003 6817
rect 59081 6752 59768 6780
rect 59909 6783 59967 6789
rect 59081 6749 59093 6752
rect 59035 6743 59093 6749
rect 59909 6749 59921 6783
rect 59955 6780 59967 6783
rect 60458 6780 60464 6792
rect 59955 6752 60464 6780
rect 59955 6749 59967 6752
rect 59909 6743 59967 6749
rect 60458 6740 60464 6752
rect 60516 6740 60522 6792
rect 61746 6740 61752 6792
rect 61804 6780 61810 6792
rect 63512 6780 63540 6888
rect 63586 6876 63592 6888
rect 63644 6876 63650 6928
rect 65426 6876 65432 6928
rect 65484 6916 65490 6928
rect 70946 6916 70952 6928
rect 65484 6888 70952 6916
rect 65484 6876 65490 6888
rect 70946 6876 70952 6888
rect 71004 6916 71010 6928
rect 74074 6916 74080 6928
rect 71004 6888 74080 6916
rect 71004 6876 71010 6888
rect 74074 6876 74080 6888
rect 74132 6876 74138 6928
rect 63678 6848 63684 6860
rect 63639 6820 63684 6848
rect 63678 6808 63684 6820
rect 63736 6808 63742 6860
rect 65521 6851 65579 6857
rect 65521 6848 65533 6851
rect 65260 6820 65533 6848
rect 61804 6752 63540 6780
rect 61804 6740 61810 6752
rect 64138 6740 64144 6792
rect 64196 6780 64202 6792
rect 64325 6783 64383 6789
rect 64325 6780 64337 6783
rect 64196 6752 64337 6780
rect 64196 6740 64202 6752
rect 64325 6749 64337 6752
rect 64371 6749 64383 6783
rect 64325 6743 64383 6749
rect 64414 6740 64420 6792
rect 64472 6789 64478 6792
rect 64472 6783 64521 6789
rect 64472 6749 64475 6783
rect 64509 6749 64521 6783
rect 64472 6743 64521 6749
rect 64472 6740 64478 6743
rect 64598 6740 64604 6792
rect 64656 6780 64662 6792
rect 64656 6752 64701 6780
rect 64656 6740 64662 6752
rect 64782 6740 64788 6792
rect 64840 6780 64846 6792
rect 65260 6780 65288 6820
rect 65521 6817 65533 6820
rect 65567 6848 65579 6851
rect 70670 6848 70676 6860
rect 65567 6820 70676 6848
rect 65567 6817 65579 6820
rect 65521 6811 65579 6817
rect 70670 6808 70676 6820
rect 70728 6808 70734 6860
rect 80514 6848 80520 6860
rect 80475 6820 80520 6848
rect 80514 6808 80520 6820
rect 80572 6808 80578 6860
rect 82906 6848 82912 6860
rect 82867 6820 82912 6848
rect 82906 6808 82912 6820
rect 82964 6808 82970 6860
rect 64840 6752 65288 6780
rect 65337 6783 65395 6789
rect 64840 6740 64846 6752
rect 65337 6749 65349 6783
rect 65383 6749 65395 6783
rect 65337 6743 65395 6749
rect 57388 6684 58572 6712
rect 57388 6672 57394 6684
rect 59354 6672 59360 6724
rect 59412 6712 59418 6724
rect 59449 6715 59507 6721
rect 59449 6712 59461 6715
rect 59412 6684 59461 6712
rect 59412 6672 59418 6684
rect 59449 6681 59461 6684
rect 59495 6681 59507 6715
rect 61470 6712 61476 6724
rect 59449 6675 59507 6681
rect 60706 6684 61476 6712
rect 55180 6616 55812 6644
rect 56873 6647 56931 6653
rect 55180 6604 55186 6616
rect 56873 6613 56885 6647
rect 56919 6644 56931 6647
rect 57698 6644 57704 6656
rect 56919 6616 57704 6644
rect 56919 6613 56931 6616
rect 56873 6607 56931 6613
rect 57698 6604 57704 6616
rect 57756 6604 57762 6656
rect 58066 6644 58072 6656
rect 58027 6616 58072 6644
rect 58066 6604 58072 6616
rect 58124 6604 58130 6656
rect 58253 6647 58311 6653
rect 58253 6613 58265 6647
rect 58299 6644 58311 6647
rect 60706 6644 60734 6684
rect 61470 6672 61476 6684
rect 61528 6672 61534 6724
rect 61654 6672 61660 6724
rect 61712 6712 61718 6724
rect 63310 6712 63316 6724
rect 61712 6684 63316 6712
rect 61712 6672 61718 6684
rect 63310 6672 63316 6684
rect 63368 6672 63374 6724
rect 64874 6712 64880 6724
rect 64835 6684 64880 6712
rect 64874 6672 64880 6684
rect 64932 6712 64938 6724
rect 65058 6712 65064 6724
rect 64932 6684 65064 6712
rect 64932 6672 64938 6684
rect 65058 6672 65064 6684
rect 65116 6672 65122 6724
rect 65150 6672 65156 6724
rect 65208 6712 65214 6724
rect 65352 6712 65380 6743
rect 65426 6740 65432 6792
rect 65484 6780 65490 6792
rect 87322 6780 87328 6792
rect 65484 6752 87328 6780
rect 65484 6740 65490 6752
rect 87322 6740 87328 6752
rect 87380 6740 87386 6792
rect 88886 6712 88892 6724
rect 65208 6684 65380 6712
rect 65444 6684 88892 6712
rect 65208 6672 65214 6684
rect 58299 6616 60734 6644
rect 58299 6613 58311 6616
rect 58253 6607 58311 6613
rect 60918 6604 60924 6656
rect 60976 6644 60982 6656
rect 61933 6647 61991 6653
rect 61933 6644 61945 6647
rect 60976 6616 61945 6644
rect 60976 6604 60982 6616
rect 61933 6613 61945 6616
rect 61979 6613 61991 6647
rect 62758 6644 62764 6656
rect 62719 6616 62764 6644
rect 61933 6607 61991 6613
rect 62758 6604 62764 6616
rect 62816 6604 62822 6656
rect 63402 6604 63408 6656
rect 63460 6644 63466 6656
rect 65444 6644 65472 6684
rect 88886 6672 88892 6684
rect 88944 6672 88950 6724
rect 63460 6616 65472 6644
rect 63460 6604 63466 6616
rect 65518 6604 65524 6656
rect 65576 6644 65582 6656
rect 67082 6644 67088 6656
rect 65576 6616 67088 6644
rect 65576 6604 65582 6616
rect 67082 6604 67088 6616
rect 67140 6644 67146 6656
rect 69750 6644 69756 6656
rect 67140 6616 69756 6644
rect 67140 6604 67146 6616
rect 69750 6604 69756 6616
rect 69808 6604 69814 6656
rect 69842 6604 69848 6656
rect 69900 6644 69906 6656
rect 80238 6644 80244 6656
rect 69900 6616 80244 6644
rect 69900 6604 69906 6616
rect 80238 6604 80244 6616
rect 80296 6604 80302 6656
rect 80330 6604 80336 6656
rect 80388 6644 80394 6656
rect 80701 6647 80759 6653
rect 80701 6644 80713 6647
rect 80388 6616 80713 6644
rect 80388 6604 80394 6616
rect 80701 6613 80713 6616
rect 80747 6613 80759 6647
rect 80701 6607 80759 6613
rect 83093 6647 83151 6653
rect 83093 6613 83105 6647
rect 83139 6644 83151 6647
rect 83182 6644 83188 6656
rect 83139 6616 83188 6644
rect 83139 6613 83151 6616
rect 83093 6607 83151 6613
rect 83182 6604 83188 6616
rect 83240 6604 83246 6656
rect 1104 6554 178848 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 34966 6554
rect 35018 6502 35030 6554
rect 35082 6502 35094 6554
rect 35146 6502 35158 6554
rect 35210 6502 65686 6554
rect 65738 6502 65750 6554
rect 65802 6502 65814 6554
rect 65866 6502 65878 6554
rect 65930 6502 96406 6554
rect 96458 6502 96470 6554
rect 96522 6502 96534 6554
rect 96586 6502 96598 6554
rect 96650 6502 127126 6554
rect 127178 6502 127190 6554
rect 127242 6502 127254 6554
rect 127306 6502 127318 6554
rect 127370 6502 157846 6554
rect 157898 6502 157910 6554
rect 157962 6502 157974 6554
rect 158026 6502 158038 6554
rect 158090 6502 178848 6554
rect 1104 6480 178848 6502
rect 21266 6440 21272 6452
rect 18524 6412 21272 6440
rect 17310 6236 17316 6248
rect 17271 6208 17316 6236
rect 17310 6196 17316 6208
rect 17368 6196 17374 6248
rect 17580 6239 17638 6245
rect 17580 6205 17592 6239
rect 17626 6236 17638 6239
rect 18046 6236 18052 6248
rect 17626 6208 18052 6236
rect 17626 6205 17638 6208
rect 17580 6199 17638 6205
rect 18046 6196 18052 6208
rect 18104 6196 18110 6248
rect 18524 6112 18552 6412
rect 21266 6400 21272 6412
rect 21324 6400 21330 6452
rect 30190 6440 30196 6452
rect 22066 6412 30196 6440
rect 20622 6332 20628 6384
rect 20680 6372 20686 6384
rect 22066 6372 22094 6412
rect 30190 6400 30196 6412
rect 30248 6400 30254 6452
rect 31754 6400 31760 6452
rect 31812 6440 31818 6452
rect 32306 6440 32312 6452
rect 31812 6412 32312 6440
rect 31812 6400 31818 6412
rect 32306 6400 32312 6412
rect 32364 6440 32370 6452
rect 33042 6440 33048 6452
rect 32364 6412 33048 6440
rect 32364 6400 32370 6412
rect 33042 6400 33048 6412
rect 33100 6400 33106 6452
rect 34422 6400 34428 6452
rect 34480 6440 34486 6452
rect 34517 6443 34575 6449
rect 34517 6440 34529 6443
rect 34480 6412 34529 6440
rect 34480 6400 34486 6412
rect 34517 6409 34529 6412
rect 34563 6409 34575 6443
rect 34517 6403 34575 6409
rect 35342 6400 35348 6452
rect 35400 6440 35406 6452
rect 36446 6440 36452 6452
rect 35400 6412 36452 6440
rect 35400 6400 35406 6412
rect 36446 6400 36452 6412
rect 36504 6400 36510 6452
rect 36538 6400 36544 6452
rect 36596 6440 36602 6452
rect 37366 6440 37372 6452
rect 36596 6412 37136 6440
rect 37327 6412 37372 6440
rect 36596 6400 36602 6412
rect 20680 6344 22094 6372
rect 29181 6375 29239 6381
rect 20680 6332 20686 6344
rect 29181 6341 29193 6375
rect 29227 6372 29239 6375
rect 30374 6372 30380 6384
rect 29227 6344 30380 6372
rect 29227 6341 29239 6344
rect 29181 6335 29239 6341
rect 30374 6332 30380 6344
rect 30432 6332 30438 6384
rect 31202 6332 31208 6384
rect 31260 6372 31266 6384
rect 31297 6375 31355 6381
rect 31297 6372 31309 6375
rect 31260 6344 31309 6372
rect 31260 6332 31266 6344
rect 31297 6341 31309 6344
rect 31343 6341 31355 6375
rect 37108 6372 37136 6412
rect 37366 6400 37372 6412
rect 37424 6400 37430 6452
rect 39761 6443 39819 6449
rect 39761 6409 39773 6443
rect 39807 6440 39819 6443
rect 40586 6440 40592 6452
rect 39807 6412 40592 6440
rect 39807 6409 39819 6412
rect 39761 6403 39819 6409
rect 40586 6400 40592 6412
rect 40644 6400 40650 6452
rect 42518 6440 42524 6452
rect 42479 6412 42524 6440
rect 42518 6400 42524 6412
rect 42576 6400 42582 6452
rect 45002 6440 45008 6452
rect 42628 6412 45008 6440
rect 37550 6372 37556 6384
rect 31297 6335 31355 6341
rect 35544 6344 36308 6372
rect 37108 6344 37556 6372
rect 35544 6316 35572 6344
rect 21174 6264 21180 6316
rect 21232 6304 21238 6316
rect 32674 6304 32680 6316
rect 21232 6276 21404 6304
rect 21232 6264 21238 6276
rect 19150 6236 19156 6248
rect 19111 6208 19156 6236
rect 19150 6196 19156 6208
rect 19208 6196 19214 6248
rect 19420 6239 19478 6245
rect 19420 6205 19432 6239
rect 19466 6236 19478 6239
rect 20714 6236 20720 6248
rect 19466 6208 20720 6236
rect 19466 6205 19478 6208
rect 19420 6199 19478 6205
rect 20714 6196 20720 6208
rect 20772 6196 20778 6248
rect 20990 6236 20996 6248
rect 20951 6208 20996 6236
rect 20990 6196 20996 6208
rect 21048 6196 21054 6248
rect 21376 6245 21404 6276
rect 28828 6276 32680 6304
rect 21269 6239 21327 6245
rect 21269 6236 21281 6239
rect 21100 6208 21281 6236
rect 18782 6128 18788 6180
rect 18840 6168 18846 6180
rect 21100 6168 21128 6208
rect 21269 6205 21281 6208
rect 21315 6205 21327 6239
rect 21269 6199 21327 6205
rect 21361 6239 21419 6245
rect 21361 6205 21373 6239
rect 21407 6205 21419 6239
rect 21361 6199 21419 6205
rect 23753 6239 23811 6245
rect 23753 6205 23765 6239
rect 23799 6236 23811 6239
rect 23842 6236 23848 6248
rect 23799 6208 23848 6236
rect 23799 6205 23811 6208
rect 23753 6199 23811 6205
rect 23842 6196 23848 6208
rect 23900 6196 23906 6248
rect 24020 6239 24078 6245
rect 24020 6205 24032 6239
rect 24066 6236 24078 6239
rect 25038 6236 25044 6248
rect 24066 6208 25044 6236
rect 24066 6205 24078 6208
rect 24020 6199 24078 6205
rect 25038 6196 25044 6208
rect 25096 6196 25102 6248
rect 27798 6236 27804 6248
rect 27759 6208 27804 6236
rect 27798 6196 27804 6208
rect 27856 6196 27862 6248
rect 28828 6236 28856 6276
rect 32674 6264 32680 6276
rect 32732 6264 32738 6316
rect 35526 6304 35532 6316
rect 27908 6208 28856 6236
rect 18840 6140 21128 6168
rect 21177 6171 21235 6177
rect 18840 6128 18846 6140
rect 21177 6137 21189 6171
rect 21223 6168 21235 6171
rect 27908 6168 27936 6208
rect 28902 6196 28908 6248
rect 28960 6236 28966 6248
rect 31018 6236 31024 6248
rect 28960 6208 31024 6236
rect 28960 6196 28966 6208
rect 31018 6196 31024 6208
rect 31076 6236 31082 6248
rect 33060 6236 33088 6290
rect 35487 6276 35532 6304
rect 35526 6264 35532 6276
rect 35584 6264 35590 6316
rect 36170 6304 36176 6316
rect 36131 6276 36176 6304
rect 36170 6264 36176 6276
rect 36228 6264 36234 6316
rect 36280 6304 36308 6344
rect 37550 6332 37556 6344
rect 37608 6332 37614 6384
rect 38292 6316 38344 6322
rect 36566 6307 36624 6313
rect 36566 6304 36578 6307
rect 36280 6276 36578 6304
rect 36566 6273 36578 6276
rect 36612 6273 36624 6307
rect 36566 6267 36624 6273
rect 36725 6307 36783 6313
rect 36725 6273 36737 6307
rect 36771 6304 36783 6307
rect 36906 6304 36912 6316
rect 36771 6276 36912 6304
rect 36771 6273 36783 6276
rect 36725 6267 36783 6273
rect 36906 6264 36912 6276
rect 36964 6304 36970 6316
rect 37826 6304 37832 6316
rect 36964 6276 37832 6304
rect 36964 6264 36970 6276
rect 37826 6264 37832 6276
rect 37884 6264 37890 6316
rect 40862 6264 40868 6316
rect 40920 6304 40926 6316
rect 40920 6276 41078 6304
rect 40920 6264 40926 6276
rect 38292 6258 38344 6264
rect 33134 6236 33140 6248
rect 31076 6208 33140 6236
rect 31076 6196 31082 6208
rect 33134 6196 33140 6208
rect 33192 6196 33198 6248
rect 33965 6239 34023 6245
rect 33965 6236 33977 6239
rect 33244 6208 33977 6236
rect 21223 6140 27936 6168
rect 28068 6171 28126 6177
rect 21223 6137 21235 6140
rect 21177 6131 21235 6137
rect 28068 6137 28080 6171
rect 28114 6168 28126 6171
rect 28994 6168 29000 6180
rect 28114 6140 29000 6168
rect 28114 6137 28126 6140
rect 28068 6131 28126 6137
rect 28994 6128 29000 6140
rect 29052 6128 29058 6180
rect 29104 6140 29316 6168
rect 16574 6060 16580 6112
rect 16632 6100 16638 6112
rect 18506 6100 18512 6112
rect 16632 6072 18512 6100
rect 16632 6060 16638 6072
rect 18506 6060 18512 6072
rect 18564 6060 18570 6112
rect 18598 6060 18604 6112
rect 18656 6100 18662 6112
rect 18693 6103 18751 6109
rect 18693 6100 18705 6103
rect 18656 6072 18705 6100
rect 18656 6060 18662 6072
rect 18693 6069 18705 6072
rect 18739 6069 18751 6103
rect 18693 6063 18751 6069
rect 19334 6060 19340 6112
rect 19392 6100 19398 6112
rect 20438 6100 20444 6112
rect 19392 6072 20444 6100
rect 19392 6060 19398 6072
rect 20438 6060 20444 6072
rect 20496 6100 20502 6112
rect 20533 6103 20591 6109
rect 20533 6100 20545 6103
rect 20496 6072 20545 6100
rect 20496 6060 20502 6072
rect 20533 6069 20545 6072
rect 20579 6069 20591 6103
rect 21542 6100 21548 6112
rect 21503 6072 21548 6100
rect 20533 6063 20591 6069
rect 21542 6060 21548 6072
rect 21600 6060 21606 6112
rect 21818 6060 21824 6112
rect 21876 6100 21882 6112
rect 25133 6103 25191 6109
rect 25133 6100 25145 6103
rect 21876 6072 25145 6100
rect 21876 6060 21882 6072
rect 25133 6069 25145 6072
rect 25179 6100 25191 6103
rect 26602 6100 26608 6112
rect 25179 6072 26608 6100
rect 25179 6069 25191 6072
rect 25133 6063 25191 6069
rect 26602 6060 26608 6072
rect 26660 6060 26666 6112
rect 28534 6060 28540 6112
rect 28592 6100 28598 6112
rect 29104 6100 29132 6140
rect 28592 6072 29132 6100
rect 29288 6100 29316 6140
rect 30558 6128 30564 6180
rect 30616 6168 30622 6180
rect 31113 6171 31171 6177
rect 31113 6168 31125 6171
rect 30616 6140 31125 6168
rect 30616 6128 30622 6140
rect 31113 6137 31125 6140
rect 31159 6137 31171 6171
rect 31113 6131 31171 6137
rect 31202 6128 31208 6180
rect 31260 6168 31266 6180
rect 33244 6177 33272 6208
rect 33965 6205 33977 6208
rect 34011 6205 34023 6239
rect 33965 6199 34023 6205
rect 35618 6196 35624 6248
rect 35676 6236 35682 6248
rect 35713 6239 35771 6245
rect 35713 6236 35725 6239
rect 35676 6208 35725 6236
rect 35676 6196 35682 6208
rect 35713 6205 35725 6208
rect 35759 6205 35771 6239
rect 35713 6199 35771 6205
rect 36446 6196 36452 6248
rect 36504 6236 36510 6248
rect 39209 6239 39267 6245
rect 39209 6236 39221 6239
rect 36504 6208 36549 6236
rect 38488 6208 39221 6236
rect 36504 6196 36510 6208
rect 33229 6171 33287 6177
rect 33229 6168 33241 6171
rect 31260 6140 33241 6168
rect 31260 6128 31266 6140
rect 33229 6137 33241 6140
rect 33275 6137 33287 6171
rect 33229 6131 33287 6137
rect 33318 6128 33324 6180
rect 33376 6168 33382 6180
rect 33505 6171 33563 6177
rect 33505 6168 33517 6171
rect 33376 6140 33517 6168
rect 33376 6128 33382 6140
rect 33505 6137 33517 6140
rect 33551 6137 33563 6171
rect 33505 6131 33563 6137
rect 33597 6171 33655 6177
rect 33597 6137 33609 6171
rect 33643 6168 33655 6171
rect 33778 6168 33784 6180
rect 33643 6140 33784 6168
rect 33643 6137 33655 6140
rect 33597 6131 33655 6137
rect 33778 6128 33784 6140
rect 33836 6128 33842 6180
rect 34256 6140 35756 6168
rect 34256 6100 34284 6140
rect 29288 6072 34284 6100
rect 34333 6103 34391 6109
rect 28592 6060 28598 6072
rect 34333 6069 34345 6103
rect 34379 6100 34391 6103
rect 34422 6100 34428 6112
rect 34379 6072 34428 6100
rect 34379 6069 34391 6072
rect 34333 6063 34391 6069
rect 34422 6060 34428 6072
rect 34480 6060 34486 6112
rect 35342 6100 35348 6112
rect 35303 6072 35348 6100
rect 35342 6060 35348 6072
rect 35400 6060 35406 6112
rect 35728 6100 35756 6140
rect 38194 6128 38200 6180
rect 38252 6168 38258 6180
rect 38488 6177 38516 6208
rect 39209 6205 39221 6208
rect 39255 6205 39267 6239
rect 41969 6239 42027 6245
rect 41969 6236 41981 6239
rect 39209 6199 39267 6205
rect 41248 6208 41981 6236
rect 38473 6171 38531 6177
rect 38473 6168 38485 6171
rect 38252 6140 38485 6168
rect 38252 6128 38258 6140
rect 38473 6137 38485 6140
rect 38519 6137 38531 6171
rect 38746 6168 38752 6180
rect 38707 6140 38752 6168
rect 38473 6131 38531 6137
rect 38746 6128 38752 6140
rect 38804 6128 38810 6180
rect 38841 6171 38899 6177
rect 38841 6137 38853 6171
rect 38887 6168 38899 6171
rect 39942 6168 39948 6180
rect 38887 6140 39948 6168
rect 38887 6137 38899 6140
rect 38841 6131 38899 6137
rect 35986 6100 35992 6112
rect 35728 6072 35992 6100
rect 35986 6060 35992 6072
rect 36044 6060 36050 6112
rect 37826 6060 37832 6112
rect 37884 6100 37890 6112
rect 38856 6100 38884 6131
rect 39942 6128 39948 6140
rect 40000 6128 40006 6180
rect 41248 6177 41276 6208
rect 41969 6205 41981 6208
rect 42015 6236 42027 6239
rect 42058 6236 42064 6248
rect 42015 6208 42064 6236
rect 42015 6205 42027 6208
rect 41969 6199 42027 6205
rect 42058 6196 42064 6208
rect 42116 6196 42122 6248
rect 42628 6236 42656 6412
rect 45002 6400 45008 6412
rect 45060 6400 45066 6452
rect 45557 6443 45615 6449
rect 45557 6409 45569 6443
rect 45603 6440 45615 6443
rect 46198 6440 46204 6452
rect 45603 6412 46204 6440
rect 45603 6409 45615 6412
rect 45557 6403 45615 6409
rect 46198 6400 46204 6412
rect 46256 6400 46262 6452
rect 46474 6440 46480 6452
rect 46308 6412 46480 6440
rect 46017 6375 46075 6381
rect 43732 6344 44496 6372
rect 43732 6313 43760 6344
rect 43717 6307 43775 6313
rect 43717 6273 43729 6307
rect 43763 6273 43775 6307
rect 43717 6267 43775 6273
rect 43806 6264 43812 6316
rect 43864 6304 43870 6316
rect 43901 6307 43959 6313
rect 43901 6304 43913 6307
rect 43864 6276 43913 6304
rect 43864 6264 43870 6276
rect 43901 6273 43913 6276
rect 43947 6273 43959 6307
rect 43901 6267 43959 6273
rect 44082 6264 44088 6316
rect 44140 6304 44146 6316
rect 44361 6307 44419 6313
rect 44361 6304 44373 6307
rect 44140 6276 44373 6304
rect 44140 6264 44146 6276
rect 44361 6273 44373 6276
rect 44407 6273 44419 6307
rect 44468 6304 44496 6344
rect 46017 6341 46029 6375
rect 46063 6372 46075 6375
rect 46308 6372 46336 6412
rect 46474 6400 46480 6412
rect 46532 6400 46538 6452
rect 46658 6400 46664 6452
rect 46716 6440 46722 6452
rect 46716 6412 47348 6440
rect 46716 6400 46722 6412
rect 47210 6372 47216 6384
rect 46063 6344 46336 6372
rect 47171 6344 47216 6372
rect 46063 6341 46075 6344
rect 46017 6335 46075 6341
rect 47210 6332 47216 6344
rect 47268 6332 47274 6384
rect 47320 6372 47348 6412
rect 47394 6400 47400 6452
rect 47452 6440 47458 6452
rect 48958 6440 48964 6452
rect 47452 6412 48964 6440
rect 47452 6400 47458 6412
rect 48958 6400 48964 6412
rect 49016 6400 49022 6452
rect 49050 6400 49056 6452
rect 49108 6440 49114 6452
rect 57974 6440 57980 6452
rect 49108 6412 57744 6440
rect 57935 6412 57980 6440
rect 49108 6400 49114 6412
rect 47578 6372 47584 6384
rect 47320 6344 47584 6372
rect 47578 6332 47584 6344
rect 47636 6372 47642 6384
rect 48774 6372 48780 6384
rect 47636 6344 48780 6372
rect 47636 6332 47642 6344
rect 48774 6332 48780 6344
rect 48832 6372 48838 6384
rect 51626 6372 51632 6384
rect 48832 6344 51632 6372
rect 48832 6332 48838 6344
rect 51626 6332 51632 6344
rect 51684 6372 51690 6384
rect 52822 6372 52828 6384
rect 51684 6344 52828 6372
rect 51684 6332 51690 6344
rect 52822 6332 52828 6344
rect 52880 6372 52886 6384
rect 54754 6372 54760 6384
rect 52880 6344 54760 6372
rect 52880 6332 52886 6344
rect 54754 6332 54760 6344
rect 54812 6372 54818 6384
rect 55306 6372 55312 6384
rect 54812 6344 55312 6372
rect 54812 6332 54818 6344
rect 55306 6332 55312 6344
rect 55364 6372 55370 6384
rect 56042 6372 56048 6384
rect 55364 6344 56048 6372
rect 55364 6332 55370 6344
rect 56042 6332 56048 6344
rect 56100 6332 56106 6384
rect 57716 6372 57744 6412
rect 57974 6400 57980 6412
rect 58032 6400 58038 6452
rect 61010 6440 61016 6452
rect 58084 6412 61016 6440
rect 58084 6372 58112 6412
rect 61010 6400 61016 6412
rect 61068 6400 61074 6452
rect 61105 6443 61163 6449
rect 61105 6409 61117 6443
rect 61151 6440 61163 6443
rect 61838 6440 61844 6452
rect 61151 6412 61844 6440
rect 61151 6409 61163 6412
rect 61105 6403 61163 6409
rect 61838 6400 61844 6412
rect 61896 6400 61902 6452
rect 62390 6400 62396 6452
rect 62448 6440 62454 6452
rect 62666 6440 62672 6452
rect 62448 6412 62672 6440
rect 62448 6400 62454 6412
rect 62666 6400 62672 6412
rect 62724 6400 62730 6452
rect 63126 6400 63132 6452
rect 63184 6440 63190 6452
rect 63184 6412 75224 6440
rect 63184 6400 63190 6412
rect 62942 6372 62948 6384
rect 56152 6344 56916 6372
rect 57716 6344 58112 6372
rect 62903 6344 62948 6372
rect 44775 6307 44833 6313
rect 44775 6304 44787 6307
rect 44468 6276 44787 6304
rect 44361 6267 44419 6273
rect 44775 6273 44787 6276
rect 44821 6304 44833 6307
rect 46106 6304 46112 6316
rect 44821 6276 46112 6304
rect 44821 6273 44833 6276
rect 44775 6267 44833 6273
rect 46106 6264 46112 6276
rect 46164 6264 46170 6316
rect 46658 6304 46664 6316
rect 46619 6276 46664 6304
rect 46658 6264 46664 6276
rect 46716 6264 46722 6316
rect 46842 6313 46848 6316
rect 46820 6307 46848 6313
rect 46820 6273 46832 6307
rect 46820 6267 46848 6273
rect 46842 6264 46848 6267
rect 46900 6264 46906 6316
rect 47854 6304 47860 6316
rect 47815 6276 47860 6304
rect 47854 6264 47860 6276
rect 47912 6264 47918 6316
rect 48590 6264 48596 6316
rect 48648 6304 48654 6316
rect 48648 6276 48912 6304
rect 48648 6264 48654 6276
rect 42260 6208 42656 6236
rect 41233 6171 41291 6177
rect 41233 6137 41245 6171
rect 41279 6137 41291 6171
rect 41233 6131 41291 6137
rect 41414 6128 41420 6180
rect 41472 6168 41478 6180
rect 41509 6171 41567 6177
rect 41509 6168 41521 6171
rect 41472 6140 41521 6168
rect 41472 6128 41478 6140
rect 41509 6137 41521 6140
rect 41555 6137 41567 6171
rect 41509 6131 41567 6137
rect 41601 6171 41659 6177
rect 41601 6137 41613 6171
rect 41647 6168 41659 6171
rect 41690 6168 41696 6180
rect 41647 6140 41696 6168
rect 41647 6137 41659 6140
rect 41601 6131 41659 6137
rect 41690 6128 41696 6140
rect 41748 6168 41754 6180
rect 42260 6168 42288 6208
rect 44634 6196 44640 6248
rect 44692 6236 44698 6248
rect 44910 6236 44916 6248
rect 44692 6208 44737 6236
rect 44871 6208 44916 6236
rect 44692 6196 44698 6208
rect 44910 6196 44916 6208
rect 44968 6196 44974 6248
rect 46934 6236 46940 6248
rect 46895 6208 46940 6236
rect 46934 6196 46940 6208
rect 46992 6196 46998 6248
rect 47670 6236 47676 6248
rect 47631 6208 47676 6236
rect 47670 6196 47676 6208
rect 47728 6196 47734 6248
rect 48774 6236 48780 6248
rect 48735 6208 48780 6236
rect 48774 6196 48780 6208
rect 48832 6196 48838 6248
rect 48884 6236 48912 6276
rect 49786 6264 49792 6316
rect 49844 6304 49850 6316
rect 49844 6276 50752 6304
rect 49844 6264 49850 6276
rect 49234 6245 49240 6248
rect 49049 6239 49107 6245
rect 49049 6236 49061 6239
rect 48884 6208 49061 6236
rect 49049 6205 49061 6208
rect 49095 6205 49107 6239
rect 49049 6199 49107 6205
rect 49191 6239 49240 6245
rect 49191 6205 49203 6239
rect 49237 6205 49240 6239
rect 49191 6199 49240 6205
rect 49234 6196 49240 6199
rect 49292 6196 49298 6248
rect 49418 6196 49424 6248
rect 49476 6236 49482 6248
rect 49973 6239 50031 6245
rect 49973 6236 49985 6239
rect 49476 6208 49985 6236
rect 49476 6196 49482 6208
rect 49973 6205 49985 6208
rect 50019 6205 50031 6239
rect 49973 6199 50031 6205
rect 50062 6196 50068 6248
rect 50120 6236 50126 6248
rect 50617 6239 50675 6245
rect 50617 6236 50629 6239
rect 50120 6208 50629 6236
rect 50120 6196 50126 6208
rect 50617 6205 50629 6208
rect 50663 6205 50675 6239
rect 50724 6236 50752 6276
rect 51074 6264 51080 6316
rect 51132 6304 51138 6316
rect 52270 6304 52276 6316
rect 51132 6276 52276 6304
rect 51132 6264 51138 6276
rect 52270 6264 52276 6276
rect 52328 6304 52334 6316
rect 55674 6304 55680 6316
rect 52328 6276 55680 6304
rect 52328 6264 52334 6276
rect 55674 6264 55680 6276
rect 55732 6264 55738 6316
rect 56152 6313 56180 6344
rect 56137 6307 56195 6313
rect 56137 6273 56149 6307
rect 56183 6273 56195 6307
rect 56686 6304 56692 6316
rect 56137 6267 56195 6273
rect 56244 6276 56692 6304
rect 51261 6239 51319 6245
rect 51261 6236 51273 6239
rect 50724 6208 51273 6236
rect 50617 6199 50675 6205
rect 51261 6205 51273 6208
rect 51307 6205 51319 6239
rect 51261 6199 51319 6205
rect 54213 6239 54271 6245
rect 54213 6205 54225 6239
rect 54259 6236 54271 6239
rect 54478 6236 54484 6248
rect 54259 6208 54484 6236
rect 54259 6205 54271 6208
rect 54213 6199 54271 6205
rect 54478 6196 54484 6208
rect 54536 6196 54542 6248
rect 56244 6236 56272 6276
rect 56686 6264 56692 6276
rect 56744 6304 56750 6316
rect 56781 6307 56839 6313
rect 56781 6304 56793 6307
rect 56744 6276 56793 6304
rect 56744 6264 56750 6276
rect 56781 6273 56793 6276
rect 56827 6273 56839 6307
rect 56888 6304 56916 6344
rect 62942 6332 62948 6344
rect 63000 6332 63006 6384
rect 64506 6372 64512 6384
rect 64467 6344 64512 6372
rect 64506 6332 64512 6344
rect 64564 6332 64570 6384
rect 65628 6344 66392 6372
rect 57238 6313 57244 6316
rect 57195 6307 57244 6313
rect 57195 6304 57207 6307
rect 56888 6276 57207 6304
rect 56781 6267 56839 6273
rect 57195 6273 57207 6276
rect 57241 6273 57244 6307
rect 57195 6267 57244 6273
rect 57238 6264 57244 6267
rect 57296 6264 57302 6316
rect 57330 6264 57336 6316
rect 57388 6304 57394 6316
rect 59262 6304 59268 6316
rect 57388 6276 57433 6304
rect 59223 6276 59268 6304
rect 57388 6264 57394 6276
rect 59262 6264 59268 6276
rect 59320 6264 59326 6316
rect 59909 6307 59967 6313
rect 59909 6304 59921 6307
rect 59372 6276 59921 6304
rect 59372 6248 59400 6276
rect 59909 6273 59921 6276
rect 59955 6273 59967 6307
rect 59909 6267 59967 6273
rect 59998 6264 60004 6316
rect 60056 6304 60062 6316
rect 60185 6307 60243 6313
rect 60185 6304 60197 6307
rect 60056 6276 60197 6304
rect 60056 6264 60062 6276
rect 60185 6273 60197 6276
rect 60231 6273 60243 6307
rect 60185 6267 60243 6273
rect 60461 6307 60519 6313
rect 60461 6273 60473 6307
rect 60507 6304 60519 6307
rect 60642 6304 60648 6316
rect 60507 6276 60648 6304
rect 60507 6273 60519 6276
rect 60461 6267 60519 6273
rect 60642 6264 60648 6276
rect 60700 6304 60706 6316
rect 62206 6304 62212 6316
rect 60700 6276 62212 6304
rect 60700 6264 60706 6276
rect 62206 6264 62212 6276
rect 62264 6304 62270 6316
rect 62393 6307 62451 6313
rect 62393 6304 62405 6307
rect 62264 6276 62405 6304
rect 62264 6264 62270 6276
rect 62393 6273 62405 6276
rect 62439 6273 62451 6307
rect 62393 6267 62451 6273
rect 62552 6307 62610 6313
rect 62552 6273 62564 6307
rect 62598 6304 62610 6307
rect 63402 6304 63408 6316
rect 62598 6276 63264 6304
rect 63363 6276 63408 6304
rect 62598 6273 62610 6276
rect 62552 6267 62610 6273
rect 55508 6208 56272 6236
rect 56321 6239 56379 6245
rect 55508 6180 55536 6208
rect 56321 6205 56333 6239
rect 56367 6205 56379 6239
rect 56321 6199 56379 6205
rect 41748 6140 42288 6168
rect 42337 6171 42395 6177
rect 41748 6128 41754 6140
rect 42337 6137 42349 6171
rect 42383 6168 42395 6171
rect 42383 6140 43852 6168
rect 42383 6137 42395 6140
rect 42337 6131 42395 6137
rect 37884 6072 38884 6100
rect 37884 6060 37890 6072
rect 39298 6060 39304 6112
rect 39356 6100 39362 6112
rect 39577 6103 39635 6109
rect 39577 6100 39589 6103
rect 39356 6072 39589 6100
rect 39356 6060 39362 6072
rect 39577 6069 39589 6072
rect 39623 6069 39635 6103
rect 39577 6063 39635 6069
rect 42426 6060 42432 6112
rect 42484 6100 42490 6112
rect 43714 6100 43720 6112
rect 42484 6072 43720 6100
rect 42484 6060 42490 6072
rect 43714 6060 43720 6072
rect 43772 6060 43778 6112
rect 43824 6100 43852 6140
rect 47854 6128 47860 6180
rect 47912 6168 47918 6180
rect 48682 6168 48688 6180
rect 47912 6140 48688 6168
rect 47912 6128 47918 6140
rect 48682 6128 48688 6140
rect 48740 6128 48746 6180
rect 48958 6128 48964 6180
rect 49016 6168 49022 6180
rect 49016 6140 49061 6168
rect 49016 6128 49022 6140
rect 53834 6128 53840 6180
rect 53892 6168 53898 6180
rect 54570 6168 54576 6180
rect 53892 6140 54576 6168
rect 53892 6128 53898 6140
rect 54570 6128 54576 6140
rect 54628 6168 54634 6180
rect 55490 6168 55496 6180
rect 54628 6140 55496 6168
rect 54628 6128 54634 6140
rect 55490 6128 55496 6140
rect 55548 6128 55554 6180
rect 56226 6128 56232 6180
rect 56284 6168 56290 6180
rect 56336 6168 56364 6199
rect 57054 6196 57060 6248
rect 57112 6236 57118 6248
rect 57112 6208 57157 6236
rect 57112 6196 57118 6208
rect 58158 6196 58164 6248
rect 58216 6236 58222 6248
rect 59354 6236 59360 6248
rect 58216 6208 59360 6236
rect 58216 6196 58222 6208
rect 59354 6196 59360 6208
rect 59412 6196 59418 6248
rect 59449 6239 59507 6245
rect 59449 6205 59461 6239
rect 59495 6236 59507 6239
rect 59630 6236 59636 6248
rect 59495 6208 59636 6236
rect 59495 6205 59507 6208
rect 59449 6199 59507 6205
rect 59630 6196 59636 6208
rect 59688 6196 59694 6248
rect 60320 6196 60326 6248
rect 60378 6236 60384 6248
rect 61746 6236 61752 6248
rect 60378 6208 60423 6236
rect 61707 6208 61752 6236
rect 60378 6196 60384 6208
rect 61746 6196 61752 6208
rect 61804 6196 61810 6248
rect 62666 6236 62672 6248
rect 62627 6208 62672 6236
rect 62666 6196 62672 6208
rect 62724 6196 62730 6248
rect 63236 6236 63264 6276
rect 63402 6264 63408 6276
rect 63460 6264 63466 6316
rect 64414 6304 64420 6316
rect 64375 6276 64420 6304
rect 64414 6264 64420 6276
rect 64472 6264 64478 6316
rect 65153 6307 65211 6313
rect 65153 6304 65165 6307
rect 64524 6276 65165 6304
rect 63589 6239 63647 6245
rect 63589 6236 63601 6239
rect 63236 6208 63601 6236
rect 63589 6205 63601 6208
rect 63635 6205 63647 6239
rect 63589 6199 63647 6205
rect 56284 6140 56364 6168
rect 56284 6128 56290 6140
rect 57882 6128 57888 6180
rect 57940 6168 57946 6180
rect 59262 6168 59268 6180
rect 57940 6140 59268 6168
rect 57940 6128 57946 6140
rect 59262 6128 59268 6140
rect 59320 6128 59326 6180
rect 63604 6168 63632 6199
rect 64046 6196 64052 6248
rect 64104 6236 64110 6248
rect 64524 6236 64552 6276
rect 65153 6273 65165 6276
rect 65199 6273 65211 6307
rect 65153 6267 65211 6273
rect 65312 6307 65370 6313
rect 65312 6273 65324 6307
rect 65358 6304 65370 6307
rect 65628 6304 65656 6344
rect 65358 6276 65656 6304
rect 65705 6307 65763 6313
rect 65358 6273 65370 6276
rect 65312 6267 65370 6273
rect 65705 6273 65717 6307
rect 65751 6304 65763 6307
rect 65794 6304 65800 6316
rect 65751 6276 65800 6304
rect 65751 6273 65763 6276
rect 65705 6267 65763 6273
rect 65794 6264 65800 6276
rect 65852 6264 65858 6316
rect 66364 6313 66392 6344
rect 69106 6332 69112 6384
rect 69164 6372 69170 6384
rect 75086 6372 75092 6384
rect 69164 6344 75092 6372
rect 69164 6332 69170 6344
rect 75086 6332 75092 6344
rect 75144 6332 75150 6384
rect 75196 6372 75224 6412
rect 75546 6400 75552 6452
rect 75604 6440 75610 6452
rect 83645 6443 83703 6449
rect 83645 6440 83657 6443
rect 75604 6412 83657 6440
rect 75604 6400 75610 6412
rect 83645 6409 83657 6412
rect 83691 6409 83703 6443
rect 83645 6403 83703 6409
rect 80606 6372 80612 6384
rect 75196 6344 80612 6372
rect 80606 6332 80612 6344
rect 80664 6332 80670 6384
rect 80885 6375 80943 6381
rect 80885 6341 80897 6375
rect 80931 6341 80943 6375
rect 80885 6335 80943 6341
rect 66349 6307 66407 6313
rect 66349 6273 66361 6307
rect 66395 6304 66407 6307
rect 69566 6304 69572 6316
rect 66395 6276 69572 6304
rect 66395 6273 66407 6276
rect 66349 6267 66407 6273
rect 69566 6264 69572 6276
rect 69624 6264 69630 6316
rect 69750 6264 69756 6316
rect 69808 6304 69814 6316
rect 69808 6276 75232 6304
rect 69808 6264 69814 6276
rect 65426 6236 65432 6248
rect 64104 6208 64552 6236
rect 65387 6208 65432 6236
rect 64104 6196 64110 6208
rect 65426 6196 65432 6208
rect 65484 6196 65490 6248
rect 65978 6196 65984 6248
rect 66036 6236 66042 6248
rect 66165 6239 66223 6245
rect 66165 6236 66177 6239
rect 66036 6208 66177 6236
rect 66036 6196 66042 6208
rect 66165 6205 66177 6208
rect 66211 6205 66223 6239
rect 66990 6236 66996 6248
rect 66951 6208 66996 6236
rect 66165 6199 66223 6205
rect 64598 6168 64604 6180
rect 63604 6140 64604 6168
rect 64598 6128 64604 6140
rect 64656 6128 64662 6180
rect 66180 6168 66208 6199
rect 66990 6196 66996 6208
rect 67048 6196 67054 6248
rect 68094 6236 68100 6248
rect 68055 6208 68100 6236
rect 68094 6196 68100 6208
rect 68152 6196 68158 6248
rect 70302 6236 70308 6248
rect 70263 6208 70308 6236
rect 70302 6196 70308 6208
rect 70360 6196 70366 6248
rect 71314 6236 71320 6248
rect 71275 6208 71320 6236
rect 71314 6196 71320 6208
rect 71372 6196 71378 6248
rect 75204 6245 75232 6276
rect 79134 6264 79140 6316
rect 79192 6304 79198 6316
rect 80900 6304 80928 6335
rect 79192 6276 80928 6304
rect 82357 6307 82415 6313
rect 79192 6264 79198 6276
rect 82357 6273 82369 6307
rect 82403 6304 82415 6307
rect 85298 6304 85304 6316
rect 82403 6276 85304 6304
rect 82403 6273 82415 6276
rect 82357 6267 82415 6273
rect 85298 6264 85304 6276
rect 85356 6264 85362 6316
rect 75181 6239 75239 6245
rect 75181 6205 75193 6239
rect 75227 6205 75239 6239
rect 77202 6236 77208 6248
rect 77163 6208 77208 6236
rect 75181 6199 75239 6205
rect 77202 6196 77208 6208
rect 77260 6196 77266 6248
rect 78306 6236 78312 6248
rect 78267 6208 78312 6236
rect 78306 6196 78312 6208
rect 78364 6196 78370 6248
rect 80054 6196 80060 6248
rect 80112 6236 80118 6248
rect 80241 6239 80299 6245
rect 80241 6236 80253 6239
rect 80112 6208 80253 6236
rect 80112 6196 80118 6208
rect 80241 6205 80253 6208
rect 80287 6205 80299 6239
rect 80241 6199 80299 6205
rect 80790 6196 80796 6248
rect 80848 6236 80854 6248
rect 81069 6239 81127 6245
rect 81069 6236 81081 6239
rect 80848 6208 81081 6236
rect 80848 6196 80854 6208
rect 81069 6205 81081 6208
rect 81115 6205 81127 6239
rect 81069 6199 81127 6205
rect 81529 6239 81587 6245
rect 81529 6205 81541 6239
rect 81575 6236 81587 6239
rect 81618 6236 81624 6248
rect 81575 6208 81624 6236
rect 81575 6205 81587 6208
rect 81529 6199 81587 6205
rect 81618 6196 81624 6208
rect 81676 6196 81682 6248
rect 81986 6196 81992 6248
rect 82044 6236 82050 6248
rect 83001 6239 83059 6245
rect 83001 6236 83013 6239
rect 82044 6208 83013 6236
rect 82044 6196 82050 6208
rect 83001 6205 83013 6208
rect 83047 6205 83059 6239
rect 83001 6199 83059 6205
rect 83090 6196 83096 6248
rect 83148 6236 83154 6248
rect 83461 6239 83519 6245
rect 83461 6236 83473 6239
rect 83148 6208 83473 6236
rect 83148 6196 83154 6208
rect 83461 6205 83473 6208
rect 83507 6205 83519 6239
rect 83461 6199 83519 6205
rect 83826 6196 83832 6248
rect 83884 6236 83890 6248
rect 84105 6239 84163 6245
rect 84105 6236 84117 6239
rect 83884 6208 84117 6236
rect 83884 6196 83890 6208
rect 84105 6205 84117 6208
rect 84151 6205 84163 6239
rect 84105 6199 84163 6205
rect 84838 6196 84844 6248
rect 84896 6236 84902 6248
rect 89806 6236 89812 6248
rect 84896 6208 89812 6236
rect 84896 6196 84902 6208
rect 89806 6196 89812 6208
rect 89864 6196 89870 6248
rect 88702 6168 88708 6180
rect 66180 6140 88708 6168
rect 88702 6128 88708 6140
rect 88760 6128 88766 6180
rect 44450 6100 44456 6112
rect 43824 6072 44456 6100
rect 44450 6060 44456 6072
rect 44508 6060 44514 6112
rect 45925 6103 45983 6109
rect 45925 6069 45937 6103
rect 45971 6100 45983 6103
rect 46566 6100 46572 6112
rect 45971 6072 46572 6100
rect 45971 6069 45983 6072
rect 45925 6063 45983 6069
rect 46566 6060 46572 6072
rect 46624 6060 46630 6112
rect 46934 6060 46940 6112
rect 46992 6100 46998 6112
rect 49329 6103 49387 6109
rect 49329 6100 49341 6103
rect 46992 6072 49341 6100
rect 46992 6060 46998 6072
rect 49329 6069 49341 6072
rect 49375 6069 49387 6103
rect 49786 6100 49792 6112
rect 49747 6072 49792 6100
rect 49329 6063 49387 6069
rect 49786 6060 49792 6072
rect 49844 6060 49850 6112
rect 50433 6103 50491 6109
rect 50433 6069 50445 6103
rect 50479 6100 50491 6103
rect 50982 6100 50988 6112
rect 50479 6072 50988 6100
rect 50479 6069 50491 6072
rect 50433 6063 50491 6069
rect 50982 6060 50988 6072
rect 51040 6060 51046 6112
rect 51077 6103 51135 6109
rect 51077 6069 51089 6103
rect 51123 6100 51135 6103
rect 53098 6100 53104 6112
rect 51123 6072 53104 6100
rect 51123 6069 51135 6072
rect 51077 6063 51135 6069
rect 53098 6060 53104 6072
rect 53156 6060 53162 6112
rect 54018 6100 54024 6112
rect 53979 6072 54024 6100
rect 54018 6060 54024 6072
rect 54076 6060 54082 6112
rect 54202 6060 54208 6112
rect 54260 6100 54266 6112
rect 61562 6100 61568 6112
rect 54260 6072 61568 6100
rect 54260 6060 54266 6072
rect 61562 6060 61568 6072
rect 61620 6060 61626 6112
rect 61657 6103 61715 6109
rect 61657 6069 61669 6103
rect 61703 6100 61715 6103
rect 63402 6100 63408 6112
rect 61703 6072 63408 6100
rect 61703 6069 61715 6072
rect 61657 6063 61715 6069
rect 63402 6060 63408 6072
rect 63460 6060 63466 6112
rect 63586 6060 63592 6112
rect 63644 6100 63650 6112
rect 65242 6100 65248 6112
rect 63644 6072 65248 6100
rect 63644 6060 63650 6072
rect 65242 6060 65248 6072
rect 65300 6060 65306 6112
rect 65426 6060 65432 6112
rect 65484 6100 65490 6112
rect 66441 6103 66499 6109
rect 66441 6100 66453 6103
rect 65484 6072 66453 6100
rect 65484 6060 65490 6072
rect 66441 6069 66453 6072
rect 66487 6069 66499 6103
rect 66806 6100 66812 6112
rect 66767 6072 66812 6100
rect 66441 6063 66499 6069
rect 66806 6060 66812 6072
rect 66864 6060 66870 6112
rect 67910 6100 67916 6112
rect 67871 6072 67916 6100
rect 67910 6060 67916 6072
rect 67968 6060 67974 6112
rect 69014 6060 69020 6112
rect 69072 6100 69078 6112
rect 70121 6103 70179 6109
rect 70121 6100 70133 6103
rect 69072 6072 70133 6100
rect 69072 6060 69078 6072
rect 70121 6069 70133 6072
rect 70167 6069 70179 6103
rect 71130 6100 71136 6112
rect 71091 6072 71136 6100
rect 70121 6063 70179 6069
rect 71130 6060 71136 6072
rect 71188 6060 71194 6112
rect 73614 6060 73620 6112
rect 73672 6100 73678 6112
rect 74997 6103 75055 6109
rect 74997 6100 75009 6103
rect 73672 6072 75009 6100
rect 73672 6060 73678 6072
rect 74997 6069 75009 6072
rect 75043 6069 75055 6103
rect 77386 6100 77392 6112
rect 77347 6072 77392 6100
rect 74997 6063 75055 6069
rect 77386 6060 77392 6072
rect 77444 6060 77450 6112
rect 78493 6103 78551 6109
rect 78493 6069 78505 6103
rect 78539 6100 78551 6103
rect 78582 6100 78588 6112
rect 78539 6072 78588 6100
rect 78539 6069 78551 6072
rect 78493 6063 78551 6069
rect 78582 6060 78588 6072
rect 78640 6060 78646 6112
rect 80422 6100 80428 6112
rect 80383 6072 80428 6100
rect 80422 6060 80428 6072
rect 80480 6060 80486 6112
rect 81713 6103 81771 6109
rect 81713 6069 81725 6103
rect 81759 6100 81771 6103
rect 82078 6100 82084 6112
rect 81759 6072 82084 6100
rect 81759 6069 81771 6072
rect 81713 6063 81771 6069
rect 82078 6060 82084 6072
rect 82136 6060 82142 6112
rect 82814 6100 82820 6112
rect 82775 6072 82820 6100
rect 82814 6060 82820 6072
rect 82872 6060 82878 6112
rect 84010 6060 84016 6112
rect 84068 6100 84074 6112
rect 84289 6103 84347 6109
rect 84289 6100 84301 6103
rect 84068 6072 84301 6100
rect 84068 6060 84074 6072
rect 84289 6069 84301 6072
rect 84335 6069 84347 6103
rect 84289 6063 84347 6069
rect 1104 6010 178848 6032
rect 1104 5958 19606 6010
rect 19658 5958 19670 6010
rect 19722 5958 19734 6010
rect 19786 5958 19798 6010
rect 19850 5958 50326 6010
rect 50378 5958 50390 6010
rect 50442 5958 50454 6010
rect 50506 5958 50518 6010
rect 50570 5958 81046 6010
rect 81098 5958 81110 6010
rect 81162 5958 81174 6010
rect 81226 5958 81238 6010
rect 81290 5958 111766 6010
rect 111818 5958 111830 6010
rect 111882 5958 111894 6010
rect 111946 5958 111958 6010
rect 112010 5958 142486 6010
rect 142538 5958 142550 6010
rect 142602 5958 142614 6010
rect 142666 5958 142678 6010
rect 142730 5958 173206 6010
rect 173258 5958 173270 6010
rect 173322 5958 173334 6010
rect 173386 5958 173398 6010
rect 173450 5958 178848 6010
rect 1104 5936 178848 5958
rect 15286 5856 15292 5908
rect 15344 5896 15350 5908
rect 17037 5899 17095 5905
rect 17037 5896 17049 5899
rect 15344 5868 17049 5896
rect 15344 5856 15350 5868
rect 17037 5865 17049 5868
rect 17083 5896 17095 5899
rect 17402 5896 17408 5908
rect 17083 5868 17408 5896
rect 17083 5865 17095 5868
rect 17037 5859 17095 5865
rect 17402 5856 17408 5868
rect 17460 5856 17466 5908
rect 18690 5856 18696 5908
rect 18748 5896 18754 5908
rect 31570 5896 31576 5908
rect 18748 5868 31576 5896
rect 18748 5856 18754 5868
rect 31570 5856 31576 5868
rect 31628 5856 31634 5908
rect 31849 5899 31907 5905
rect 31849 5865 31861 5899
rect 31895 5896 31907 5899
rect 31938 5896 31944 5908
rect 31895 5868 31944 5896
rect 31895 5865 31907 5868
rect 31849 5859 31907 5865
rect 31938 5856 31944 5868
rect 31996 5856 32002 5908
rect 33686 5896 33692 5908
rect 32140 5868 33692 5896
rect 15924 5831 15982 5837
rect 15924 5797 15936 5831
rect 15970 5828 15982 5831
rect 22094 5828 22100 5840
rect 15970 5800 22100 5828
rect 15970 5797 15982 5800
rect 15924 5791 15982 5797
rect 22094 5788 22100 5800
rect 22152 5788 22158 5840
rect 23100 5831 23158 5837
rect 23100 5797 23112 5831
rect 23146 5828 23158 5831
rect 23474 5828 23480 5840
rect 23146 5800 23480 5828
rect 23146 5797 23158 5800
rect 23100 5791 23158 5797
rect 23474 5788 23480 5800
rect 23532 5788 23538 5840
rect 25492 5831 25550 5837
rect 25492 5797 25504 5831
rect 25538 5828 25550 5831
rect 26326 5828 26332 5840
rect 25538 5800 26332 5828
rect 25538 5797 25550 5800
rect 25492 5791 25550 5797
rect 26326 5788 26332 5800
rect 26384 5788 26390 5840
rect 27332 5831 27390 5837
rect 27332 5797 27344 5831
rect 27378 5828 27390 5831
rect 27430 5828 27436 5840
rect 27378 5800 27436 5828
rect 27378 5797 27390 5800
rect 27332 5791 27390 5797
rect 27430 5788 27436 5800
rect 27488 5788 27494 5840
rect 32030 5828 32036 5840
rect 30484 5800 32036 5828
rect 15657 5763 15715 5769
rect 15657 5729 15669 5763
rect 15703 5760 15715 5763
rect 17310 5760 17316 5772
rect 15703 5732 17316 5760
rect 15703 5729 15715 5732
rect 15657 5723 15715 5729
rect 17310 5720 17316 5732
rect 17368 5720 17374 5772
rect 17764 5763 17822 5769
rect 17764 5729 17776 5763
rect 17810 5760 17822 5763
rect 20714 5760 20720 5772
rect 17810 5732 20720 5760
rect 17810 5729 17822 5732
rect 17764 5723 17822 5729
rect 20714 5720 20720 5732
rect 20772 5720 20778 5772
rect 20892 5763 20950 5769
rect 20892 5729 20904 5763
rect 20938 5760 20950 5763
rect 22278 5760 22284 5772
rect 20938 5732 22284 5760
rect 20938 5729 20950 5732
rect 20892 5723 20950 5729
rect 22278 5720 22284 5732
rect 22336 5720 22342 5772
rect 22833 5763 22891 5769
rect 22833 5729 22845 5763
rect 22879 5760 22891 5763
rect 23842 5760 23848 5772
rect 22879 5732 23848 5760
rect 22879 5729 22891 5732
rect 22833 5723 22891 5729
rect 17497 5695 17555 5701
rect 17497 5661 17509 5695
rect 17543 5661 17555 5695
rect 17497 5655 17555 5661
rect 17310 5516 17316 5568
rect 17368 5556 17374 5568
rect 17512 5556 17540 5655
rect 19150 5652 19156 5704
rect 19208 5692 19214 5704
rect 20622 5692 20628 5704
rect 19208 5664 20628 5692
rect 19208 5652 19214 5664
rect 20622 5652 20628 5664
rect 20680 5652 20686 5704
rect 21634 5652 21640 5704
rect 21692 5692 21698 5704
rect 22848 5692 22876 5723
rect 23842 5720 23848 5732
rect 23900 5760 23906 5772
rect 25225 5763 25283 5769
rect 25225 5760 25237 5763
rect 23900 5732 25237 5760
rect 23900 5720 23906 5732
rect 25225 5729 25237 5732
rect 25271 5760 25283 5763
rect 27065 5763 27123 5769
rect 27065 5760 27077 5763
rect 25271 5732 27077 5760
rect 25271 5729 25283 5732
rect 25225 5723 25283 5729
rect 27065 5729 27077 5732
rect 27111 5760 27123 5763
rect 27798 5760 27804 5772
rect 27111 5732 27804 5760
rect 27111 5729 27123 5732
rect 27065 5723 27123 5729
rect 27798 5720 27804 5732
rect 27856 5760 27862 5772
rect 29270 5760 29276 5772
rect 27856 5732 29276 5760
rect 27856 5720 27862 5732
rect 29270 5720 29276 5732
rect 29328 5760 29334 5772
rect 30484 5769 30512 5800
rect 32030 5788 32036 5800
rect 32088 5788 32094 5840
rect 30469 5763 30527 5769
rect 30469 5760 30481 5763
rect 29328 5732 30481 5760
rect 29328 5720 29334 5732
rect 30469 5729 30481 5732
rect 30515 5729 30527 5763
rect 30469 5723 30527 5729
rect 30736 5763 30794 5769
rect 30736 5729 30748 5763
rect 30782 5760 30794 5763
rect 32140 5760 32168 5868
rect 33686 5856 33692 5868
rect 33744 5856 33750 5908
rect 34793 5899 34851 5905
rect 34793 5865 34805 5899
rect 34839 5896 34851 5899
rect 40494 5896 40500 5908
rect 34839 5868 40500 5896
rect 34839 5865 34851 5868
rect 34793 5859 34851 5865
rect 40494 5856 40500 5868
rect 40552 5856 40558 5908
rect 43530 5856 43536 5908
rect 43588 5896 43594 5908
rect 45830 5896 45836 5908
rect 43588 5868 45836 5896
rect 43588 5856 43594 5868
rect 45830 5856 45836 5868
rect 45888 5856 45894 5908
rect 46201 5899 46259 5905
rect 46201 5865 46213 5899
rect 46247 5896 46259 5899
rect 46382 5896 46388 5908
rect 46247 5868 46388 5896
rect 46247 5865 46259 5868
rect 46201 5859 46259 5865
rect 46382 5856 46388 5868
rect 46440 5856 46446 5908
rect 47210 5856 47216 5908
rect 47268 5896 47274 5908
rect 47394 5896 47400 5908
rect 47268 5868 47400 5896
rect 47268 5856 47274 5868
rect 47394 5856 47400 5868
rect 47452 5856 47458 5908
rect 47486 5856 47492 5908
rect 47544 5896 47550 5908
rect 49418 5896 49424 5908
rect 47544 5868 49424 5896
rect 47544 5856 47550 5868
rect 49418 5856 49424 5868
rect 49476 5856 49482 5908
rect 55030 5896 55036 5908
rect 53392 5868 54892 5896
rect 54991 5868 55036 5896
rect 37182 5828 37188 5840
rect 30782 5732 32168 5760
rect 32232 5800 34652 5828
rect 30782 5729 30794 5732
rect 30736 5723 30794 5729
rect 21692 5664 22876 5692
rect 21692 5652 21698 5664
rect 31570 5652 31576 5704
rect 31628 5692 31634 5704
rect 31846 5692 31852 5704
rect 31628 5664 31852 5692
rect 31628 5652 31634 5664
rect 31846 5652 31852 5664
rect 31904 5652 31910 5704
rect 19168 5624 19196 5652
rect 18432 5596 19196 5624
rect 28445 5627 28503 5633
rect 18432 5556 18460 5596
rect 28445 5593 28457 5627
rect 28491 5624 28503 5627
rect 28718 5624 28724 5636
rect 28491 5596 28724 5624
rect 28491 5593 28503 5596
rect 28445 5587 28503 5593
rect 17368 5528 18460 5556
rect 17368 5516 17374 5528
rect 18506 5516 18512 5568
rect 18564 5556 18570 5568
rect 18877 5559 18935 5565
rect 18877 5556 18889 5559
rect 18564 5528 18889 5556
rect 18564 5516 18570 5528
rect 18877 5525 18889 5528
rect 18923 5525 18935 5559
rect 18877 5519 18935 5525
rect 21634 5516 21640 5568
rect 21692 5556 21698 5568
rect 22002 5556 22008 5568
rect 21692 5528 22008 5556
rect 21692 5516 21698 5528
rect 22002 5516 22008 5528
rect 22060 5516 22066 5568
rect 24210 5516 24216 5568
rect 24268 5556 24274 5568
rect 26602 5556 26608 5568
rect 24268 5528 24313 5556
rect 26563 5528 26608 5556
rect 24268 5516 24274 5528
rect 26602 5516 26608 5528
rect 26660 5556 26666 5568
rect 27798 5556 27804 5568
rect 26660 5528 27804 5556
rect 26660 5516 26666 5528
rect 27798 5516 27804 5528
rect 27856 5516 27862 5568
rect 27982 5516 27988 5568
rect 28040 5556 28046 5568
rect 28460 5556 28488 5587
rect 28718 5584 28724 5596
rect 28776 5584 28782 5636
rect 32232 5624 32260 5800
rect 32576 5763 32634 5769
rect 32576 5729 32588 5763
rect 32622 5760 32634 5763
rect 33870 5760 33876 5772
rect 32622 5732 33876 5760
rect 32622 5729 32634 5732
rect 32576 5723 32634 5729
rect 33870 5720 33876 5732
rect 33928 5720 33934 5772
rect 34624 5769 34652 5800
rect 37108 5800 37188 5828
rect 34609 5763 34667 5769
rect 34609 5729 34621 5763
rect 34655 5729 34667 5763
rect 34609 5723 34667 5729
rect 35434 5720 35440 5772
rect 35492 5760 35498 5772
rect 35897 5763 35955 5769
rect 35897 5760 35909 5763
rect 35492 5732 35909 5760
rect 35492 5720 35498 5732
rect 35897 5729 35909 5732
rect 35943 5729 35955 5763
rect 35897 5723 35955 5729
rect 36262 5720 36268 5772
rect 36320 5760 36326 5772
rect 37108 5769 37136 5800
rect 37182 5788 37188 5800
rect 37240 5788 37246 5840
rect 41230 5828 41236 5840
rect 38028 5800 41236 5828
rect 36449 5763 36507 5769
rect 36449 5760 36461 5763
rect 36320 5732 36461 5760
rect 36320 5720 36326 5732
rect 36449 5729 36461 5732
rect 36495 5729 36507 5763
rect 36449 5723 36507 5729
rect 37093 5763 37151 5769
rect 37093 5729 37105 5763
rect 37139 5729 37151 5763
rect 38028 5760 38056 5800
rect 41230 5788 41236 5800
rect 41288 5788 41294 5840
rect 42144 5831 42202 5837
rect 42144 5797 42156 5831
rect 42190 5828 42202 5831
rect 45922 5828 45928 5840
rect 42190 5800 45928 5828
rect 42190 5797 42202 5800
rect 42144 5791 42202 5797
rect 45922 5788 45928 5800
rect 45980 5788 45986 5840
rect 46109 5831 46167 5837
rect 46109 5797 46121 5831
rect 46155 5828 46167 5831
rect 48768 5831 48826 5837
rect 46155 5800 46336 5828
rect 46155 5797 46167 5800
rect 46109 5791 46167 5797
rect 37093 5723 37151 5729
rect 37200 5732 38056 5760
rect 32309 5695 32367 5701
rect 32309 5661 32321 5695
rect 32355 5661 32367 5695
rect 37200 5692 37228 5732
rect 38102 5720 38108 5772
rect 38160 5760 38166 5772
rect 39393 5763 39451 5769
rect 39393 5760 39405 5763
rect 38160 5732 39405 5760
rect 38160 5720 38166 5732
rect 39393 5729 39405 5732
rect 39439 5729 39451 5763
rect 39393 5723 39451 5729
rect 39482 5720 39488 5772
rect 39540 5760 39546 5772
rect 41417 5763 41475 5769
rect 41417 5760 41429 5763
rect 39540 5732 41429 5760
rect 39540 5720 39546 5732
rect 41417 5729 41429 5732
rect 41463 5729 41475 5763
rect 43806 5760 43812 5772
rect 41417 5723 41475 5729
rect 41800 5732 43812 5760
rect 32309 5655 32367 5661
rect 37016 5664 37228 5692
rect 37369 5695 37427 5701
rect 31726 5596 32260 5624
rect 28040 5528 28488 5556
rect 28040 5516 28046 5528
rect 30650 5516 30656 5568
rect 30708 5556 30714 5568
rect 31726 5556 31754 5596
rect 30708 5528 31754 5556
rect 30708 5516 30714 5528
rect 32030 5516 32036 5568
rect 32088 5556 32094 5568
rect 32324 5556 32352 5655
rect 33244 5596 33824 5624
rect 32088 5528 32352 5556
rect 32088 5516 32094 5528
rect 32674 5516 32680 5568
rect 32732 5556 32738 5568
rect 33244 5556 33272 5596
rect 33686 5556 33692 5568
rect 32732 5528 33272 5556
rect 33647 5528 33692 5556
rect 32732 5516 32738 5528
rect 33686 5516 33692 5528
rect 33744 5516 33750 5568
rect 33796 5556 33824 5596
rect 34054 5584 34060 5636
rect 34112 5624 34118 5636
rect 37016 5624 37044 5664
rect 37369 5661 37381 5695
rect 37415 5692 37427 5695
rect 37550 5692 37556 5704
rect 37415 5664 37556 5692
rect 37415 5661 37427 5664
rect 37369 5655 37427 5661
rect 37550 5652 37556 5664
rect 37608 5692 37614 5704
rect 41800 5692 41828 5732
rect 43806 5720 43812 5732
rect 43864 5720 43870 5772
rect 43984 5763 44042 5769
rect 43984 5729 43996 5763
rect 44030 5760 44042 5763
rect 44030 5732 46152 5760
rect 44030 5729 44042 5732
rect 43984 5723 44042 5729
rect 37608 5664 41828 5692
rect 37608 5652 37614 5664
rect 41874 5652 41880 5704
rect 41932 5692 41938 5704
rect 41932 5664 41977 5692
rect 41932 5652 41938 5664
rect 43438 5652 43444 5704
rect 43496 5692 43502 5704
rect 43717 5695 43775 5701
rect 43717 5692 43729 5695
rect 43496 5664 43729 5692
rect 43496 5652 43502 5664
rect 43717 5661 43729 5664
rect 43763 5661 43775 5695
rect 43717 5655 43775 5661
rect 41782 5624 41788 5636
rect 34112 5596 37044 5624
rect 38396 5596 41788 5624
rect 34112 5584 34118 5596
rect 35434 5556 35440 5568
rect 33796 5528 35440 5556
rect 35434 5516 35440 5528
rect 35492 5516 35498 5568
rect 35713 5559 35771 5565
rect 35713 5525 35725 5559
rect 35759 5556 35771 5559
rect 36538 5556 36544 5568
rect 35759 5528 36544 5556
rect 35759 5525 35771 5528
rect 35713 5519 35771 5525
rect 36538 5516 36544 5528
rect 36596 5516 36602 5568
rect 36633 5559 36691 5565
rect 36633 5525 36645 5559
rect 36679 5556 36691 5559
rect 38396 5556 38424 5596
rect 41782 5584 41788 5596
rect 41840 5584 41846 5636
rect 43254 5624 43260 5636
rect 43215 5596 43260 5624
rect 43254 5584 43260 5596
rect 43312 5584 43318 5636
rect 46014 5624 46020 5636
rect 44652 5596 46020 5624
rect 38654 5556 38660 5568
rect 36679 5528 38424 5556
rect 38615 5528 38660 5556
rect 36679 5525 36691 5528
rect 36633 5519 36691 5525
rect 38654 5516 38660 5528
rect 38712 5516 38718 5568
rect 39209 5559 39267 5565
rect 39209 5525 39221 5559
rect 39255 5556 39267 5559
rect 41138 5556 41144 5568
rect 39255 5528 41144 5556
rect 39255 5525 39267 5528
rect 39209 5519 39267 5525
rect 41138 5516 41144 5528
rect 41196 5516 41202 5568
rect 41233 5559 41291 5565
rect 41233 5525 41245 5559
rect 41279 5556 41291 5559
rect 42610 5556 42616 5568
rect 41279 5528 42616 5556
rect 41279 5525 41291 5528
rect 41233 5519 41291 5525
rect 42610 5516 42616 5528
rect 42668 5516 42674 5568
rect 42794 5516 42800 5568
rect 42852 5556 42858 5568
rect 44652 5556 44680 5596
rect 46014 5584 46020 5596
rect 46072 5584 46078 5636
rect 42852 5528 44680 5556
rect 42852 5516 42858 5528
rect 45002 5516 45008 5568
rect 45060 5556 45066 5568
rect 45097 5559 45155 5565
rect 45097 5556 45109 5559
rect 45060 5528 45109 5556
rect 45060 5516 45066 5528
rect 45097 5525 45109 5528
rect 45143 5525 45155 5559
rect 46124 5556 46152 5732
rect 46308 5692 46336 5800
rect 48768 5797 48780 5831
rect 48814 5828 48826 5831
rect 49510 5828 49516 5840
rect 48814 5800 49516 5828
rect 48814 5797 48826 5800
rect 48768 5791 48826 5797
rect 49510 5788 49516 5800
rect 49568 5788 49574 5840
rect 46842 5720 46848 5772
rect 46900 5760 46906 5772
rect 47118 5760 47124 5772
rect 46900 5732 46945 5760
rect 47079 5732 47124 5760
rect 46900 5720 46906 5732
rect 47118 5720 47124 5732
rect 47176 5720 47182 5772
rect 48038 5760 48044 5772
rect 47688 5732 48044 5760
rect 46658 5692 46664 5704
rect 46308 5664 46664 5692
rect 46658 5652 46664 5664
rect 46716 5652 46722 5704
rect 47004 5695 47062 5701
rect 47004 5661 47016 5695
rect 47050 5692 47062 5695
rect 47688 5692 47716 5732
rect 48038 5720 48044 5732
rect 48096 5720 48102 5772
rect 49050 5760 49056 5772
rect 48332 5732 49056 5760
rect 47050 5664 47716 5692
rect 47857 5695 47915 5701
rect 47050 5661 47062 5664
rect 47004 5655 47062 5661
rect 47857 5661 47869 5695
rect 47903 5692 47915 5695
rect 48332 5692 48360 5732
rect 49050 5720 49056 5732
rect 49108 5720 49114 5772
rect 52086 5760 52092 5772
rect 52047 5732 52092 5760
rect 52086 5720 52092 5732
rect 52144 5720 52150 5772
rect 53190 5760 53196 5772
rect 53151 5732 53196 5760
rect 53190 5720 53196 5732
rect 53248 5720 53254 5772
rect 53392 5769 53420 5868
rect 54864 5828 54892 5868
rect 55030 5856 55036 5868
rect 55088 5856 55094 5908
rect 56686 5856 56692 5908
rect 56744 5896 56750 5908
rect 58526 5896 58532 5908
rect 56744 5868 57192 5896
rect 56744 5856 56750 5868
rect 54864 5800 57100 5828
rect 54294 5769 54300 5772
rect 53377 5763 53435 5769
rect 53377 5729 53389 5763
rect 53423 5729 53435 5763
rect 53377 5723 53435 5729
rect 54251 5763 54300 5769
rect 54251 5729 54263 5763
rect 54297 5729 54300 5763
rect 54251 5723 54300 5729
rect 54294 5720 54300 5723
rect 54352 5720 54358 5772
rect 55674 5760 55680 5772
rect 55635 5732 55680 5760
rect 55674 5720 55680 5732
rect 55732 5720 55738 5772
rect 47903 5664 48360 5692
rect 48501 5695 48559 5701
rect 47903 5661 47915 5664
rect 47857 5655 47915 5661
rect 48501 5661 48513 5695
rect 48547 5661 48559 5695
rect 48501 5655 48559 5661
rect 47394 5624 47400 5636
rect 47355 5596 47400 5624
rect 47394 5584 47400 5596
rect 47452 5584 47458 5636
rect 47486 5584 47492 5636
rect 47544 5624 47550 5636
rect 47872 5624 47900 5655
rect 48516 5624 48544 5655
rect 52178 5652 52184 5704
rect 52236 5692 52242 5704
rect 53834 5692 53840 5704
rect 52236 5664 53840 5692
rect 52236 5652 52242 5664
rect 53834 5652 53840 5664
rect 53892 5652 53898 5704
rect 54113 5695 54171 5701
rect 54113 5692 54125 5695
rect 53944 5664 54125 5692
rect 53944 5624 53972 5664
rect 54113 5661 54125 5664
rect 54159 5661 54171 5695
rect 54113 5655 54171 5661
rect 54387 5695 54445 5701
rect 54387 5661 54399 5695
rect 54433 5692 54445 5695
rect 54754 5692 54760 5704
rect 54433 5664 54760 5692
rect 54433 5661 54445 5664
rect 54387 5655 54445 5661
rect 54754 5652 54760 5664
rect 54812 5652 54818 5704
rect 47544 5596 47900 5624
rect 47964 5596 48544 5624
rect 53760 5596 53972 5624
rect 47544 5584 47550 5596
rect 47302 5556 47308 5568
rect 46124 5528 47308 5556
rect 45097 5519 45155 5525
rect 47302 5516 47308 5528
rect 47360 5516 47366 5568
rect 47854 5516 47860 5568
rect 47912 5556 47918 5568
rect 47964 5556 47992 5596
rect 47912 5528 47992 5556
rect 47912 5516 47918 5528
rect 48038 5516 48044 5568
rect 48096 5556 48102 5568
rect 49881 5559 49939 5565
rect 49881 5556 49893 5559
rect 48096 5528 49893 5556
rect 48096 5516 48102 5528
rect 49881 5525 49893 5528
rect 49927 5556 49939 5559
rect 49970 5556 49976 5568
rect 49927 5528 49976 5556
rect 49927 5525 49939 5528
rect 49881 5519 49939 5525
rect 49970 5516 49976 5528
rect 50028 5516 50034 5568
rect 51905 5559 51963 5565
rect 51905 5525 51917 5559
rect 51951 5556 51963 5559
rect 52822 5556 52828 5568
rect 51951 5528 52828 5556
rect 51951 5525 51963 5528
rect 51905 5519 51963 5525
rect 52822 5516 52828 5528
rect 52880 5516 52886 5568
rect 52914 5516 52920 5568
rect 52972 5556 52978 5568
rect 53760 5556 53788 5596
rect 52972 5528 53788 5556
rect 55493 5559 55551 5565
rect 52972 5516 52978 5528
rect 55493 5525 55505 5559
rect 55539 5556 55551 5559
rect 56042 5556 56048 5568
rect 55539 5528 56048 5556
rect 55539 5525 55551 5528
rect 55493 5519 55551 5525
rect 56042 5516 56048 5528
rect 56100 5516 56106 5568
rect 57072 5556 57100 5800
rect 57164 5624 57192 5868
rect 57532 5868 58532 5896
rect 57532 5769 57560 5868
rect 58526 5856 58532 5868
rect 58584 5856 58590 5908
rect 59357 5899 59415 5905
rect 59357 5865 59369 5899
rect 59403 5896 59415 5899
rect 59538 5896 59544 5908
rect 59403 5868 59544 5896
rect 59403 5865 59415 5868
rect 59357 5859 59415 5865
rect 59538 5856 59544 5868
rect 59596 5856 59602 5908
rect 63126 5896 63132 5908
rect 60568 5868 63132 5896
rect 59262 5788 59268 5840
rect 59320 5828 59326 5840
rect 60568 5828 60596 5868
rect 63126 5856 63132 5868
rect 63184 5856 63190 5908
rect 63313 5899 63371 5905
rect 63313 5865 63325 5899
rect 63359 5896 63371 5899
rect 63359 5868 65104 5896
rect 63359 5865 63371 5868
rect 63313 5859 63371 5865
rect 59320 5800 60596 5828
rect 59320 5788 59326 5800
rect 57517 5763 57575 5769
rect 57517 5729 57529 5763
rect 57563 5729 57575 5763
rect 57517 5723 57575 5729
rect 58526 5720 58532 5772
rect 58584 5769 58590 5772
rect 58584 5763 58612 5769
rect 58600 5729 58612 5763
rect 58710 5760 58716 5772
rect 58671 5732 58716 5760
rect 58584 5723 58612 5729
rect 58584 5720 58590 5723
rect 58710 5720 58716 5732
rect 58768 5720 58774 5772
rect 59446 5720 59452 5772
rect 59504 5760 59510 5772
rect 60001 5763 60059 5769
rect 60001 5760 60013 5763
rect 59504 5732 60013 5760
rect 59504 5720 59510 5732
rect 60001 5729 60013 5732
rect 60047 5729 60059 5763
rect 60001 5723 60059 5729
rect 60642 5720 60648 5772
rect 60700 5769 60706 5772
rect 60700 5760 60711 5769
rect 60700 5732 60745 5760
rect 60700 5723 60711 5732
rect 60700 5720 60706 5723
rect 62114 5720 62120 5772
rect 62172 5760 62178 5772
rect 62942 5760 62948 5772
rect 62172 5732 62948 5760
rect 62172 5720 62178 5732
rect 62942 5720 62948 5732
rect 63000 5760 63006 5772
rect 63402 5760 63408 5772
rect 63000 5732 63408 5760
rect 63000 5720 63006 5732
rect 63402 5720 63408 5732
rect 63460 5720 63466 5772
rect 64230 5769 64236 5772
rect 64208 5763 64236 5769
rect 64208 5729 64220 5763
rect 64208 5723 64236 5729
rect 64230 5720 64236 5723
rect 64288 5720 64294 5772
rect 57606 5652 57612 5704
rect 57664 5692 57670 5704
rect 57701 5695 57759 5701
rect 57701 5692 57713 5695
rect 57664 5664 57713 5692
rect 57664 5652 57670 5664
rect 57701 5661 57713 5664
rect 57747 5661 57759 5695
rect 57701 5655 57759 5661
rect 58250 5652 58256 5704
rect 58308 5692 58314 5704
rect 58437 5695 58495 5701
rect 58437 5692 58449 5695
rect 58308 5664 58449 5692
rect 58308 5652 58314 5664
rect 58437 5661 58449 5664
rect 58483 5661 58495 5695
rect 58437 5655 58495 5661
rect 62298 5652 62304 5704
rect 62356 5692 62362 5704
rect 64046 5692 64052 5704
rect 62356 5664 64052 5692
rect 62356 5652 62362 5664
rect 64046 5652 64052 5664
rect 64104 5652 64110 5704
rect 64322 5692 64328 5704
rect 64283 5664 64328 5692
rect 64322 5652 64328 5664
rect 64380 5652 64386 5704
rect 65076 5701 65104 5868
rect 65242 5856 65248 5908
rect 65300 5896 65306 5908
rect 68002 5896 68008 5908
rect 65300 5868 68008 5896
rect 65300 5856 65306 5868
rect 68002 5856 68008 5868
rect 68060 5896 68066 5908
rect 68922 5896 68928 5908
rect 68060 5868 68928 5896
rect 68060 5856 68066 5868
rect 68922 5856 68928 5868
rect 68980 5856 68986 5908
rect 72421 5899 72479 5905
rect 72421 5865 72433 5899
rect 72467 5896 72479 5899
rect 73706 5896 73712 5908
rect 72467 5868 73712 5896
rect 72467 5865 72479 5868
rect 72421 5859 72479 5865
rect 73706 5856 73712 5868
rect 73764 5856 73770 5908
rect 75086 5856 75092 5908
rect 75144 5896 75150 5908
rect 77665 5899 77723 5905
rect 77665 5896 77677 5899
rect 75144 5868 77677 5896
rect 75144 5856 75150 5868
rect 77665 5865 77677 5868
rect 77711 5865 77723 5899
rect 77665 5859 77723 5865
rect 77754 5856 77760 5908
rect 77812 5896 77818 5908
rect 82814 5896 82820 5908
rect 77812 5868 82820 5896
rect 77812 5856 77818 5868
rect 82814 5856 82820 5868
rect 82872 5856 82878 5908
rect 83093 5899 83151 5905
rect 83093 5865 83105 5899
rect 83139 5896 83151 5899
rect 89070 5896 89076 5908
rect 83139 5868 89076 5896
rect 83139 5865 83151 5868
rect 83093 5859 83151 5865
rect 89070 5856 89076 5868
rect 89128 5856 89134 5908
rect 65518 5788 65524 5840
rect 65576 5828 65582 5840
rect 72050 5828 72056 5840
rect 65576 5800 72056 5828
rect 65576 5788 65582 5800
rect 72050 5788 72056 5800
rect 72108 5788 72114 5840
rect 72528 5800 79548 5828
rect 65334 5720 65340 5772
rect 65392 5760 65398 5772
rect 65889 5763 65947 5769
rect 65889 5760 65901 5763
rect 65392 5732 65901 5760
rect 65392 5720 65398 5732
rect 65889 5729 65901 5732
rect 65935 5729 65947 5763
rect 65889 5723 65947 5729
rect 68922 5720 68928 5772
rect 68980 5760 68986 5772
rect 69017 5763 69075 5769
rect 69017 5760 69029 5763
rect 68980 5732 69029 5760
rect 68980 5720 68986 5732
rect 69017 5729 69029 5732
rect 69063 5729 69075 5763
rect 69017 5723 69075 5729
rect 69658 5720 69664 5772
rect 69716 5760 69722 5772
rect 72528 5760 72556 5800
rect 69716 5732 72556 5760
rect 69716 5720 69722 5732
rect 72602 5720 72608 5772
rect 72660 5760 72666 5772
rect 73246 5760 73252 5772
rect 72660 5732 72705 5760
rect 73207 5732 73252 5760
rect 72660 5720 72666 5732
rect 73246 5720 73252 5732
rect 73304 5720 73310 5772
rect 74074 5760 74080 5772
rect 74035 5732 74080 5760
rect 74074 5720 74080 5732
rect 74132 5720 74138 5772
rect 74626 5720 74632 5772
rect 74684 5760 74690 5772
rect 77570 5760 77576 5772
rect 74684 5732 77576 5760
rect 74684 5720 74690 5732
rect 77570 5720 77576 5732
rect 77628 5720 77634 5772
rect 77662 5720 77668 5772
rect 77720 5760 77726 5772
rect 77849 5763 77907 5769
rect 77849 5760 77861 5763
rect 77720 5732 77861 5760
rect 77720 5720 77726 5732
rect 77849 5729 77861 5732
rect 77895 5729 77907 5763
rect 77849 5723 77907 5729
rect 78674 5720 78680 5772
rect 78732 5760 78738 5772
rect 79410 5760 79416 5772
rect 78732 5732 79416 5760
rect 78732 5720 78738 5732
rect 79410 5720 79416 5732
rect 79468 5720 79474 5772
rect 65061 5695 65119 5701
rect 65061 5661 65073 5695
rect 65107 5661 65119 5695
rect 65061 5655 65119 5661
rect 58158 5624 58164 5636
rect 57164 5596 58164 5624
rect 58158 5584 58164 5596
rect 58216 5584 58222 5636
rect 64598 5624 64604 5636
rect 59372 5596 63724 5624
rect 64559 5596 64604 5624
rect 59372 5556 59400 5596
rect 57072 5528 59400 5556
rect 59446 5516 59452 5568
rect 59504 5556 59510 5568
rect 59817 5559 59875 5565
rect 59817 5556 59829 5559
rect 59504 5528 59829 5556
rect 59504 5516 59510 5528
rect 59817 5525 59829 5528
rect 59863 5525 59875 5559
rect 59817 5519 59875 5525
rect 59906 5516 59912 5568
rect 59964 5556 59970 5568
rect 60461 5559 60519 5565
rect 60461 5556 60473 5559
rect 59964 5528 60473 5556
rect 59964 5516 59970 5528
rect 60461 5525 60473 5528
rect 60507 5525 60519 5559
rect 60461 5519 60519 5525
rect 63405 5559 63463 5565
rect 63405 5525 63417 5559
rect 63451 5556 63463 5559
rect 63586 5556 63592 5568
rect 63451 5528 63592 5556
rect 63451 5525 63463 5528
rect 63405 5519 63463 5525
rect 63586 5516 63592 5528
rect 63644 5516 63650 5568
rect 63696 5556 63724 5596
rect 64598 5584 64604 5596
rect 64656 5624 64662 5636
rect 64874 5624 64880 5636
rect 64656 5596 64880 5624
rect 64656 5584 64662 5596
rect 64874 5584 64880 5596
rect 64932 5584 64938 5636
rect 65076 5624 65104 5655
rect 65242 5652 65248 5704
rect 65300 5692 65306 5704
rect 68186 5692 68192 5704
rect 65300 5664 68192 5692
rect 65300 5652 65306 5664
rect 68186 5652 68192 5664
rect 68244 5652 68250 5704
rect 70210 5652 70216 5704
rect 70268 5692 70274 5704
rect 79134 5692 79140 5704
rect 70268 5664 79140 5692
rect 70268 5652 70274 5664
rect 79134 5652 79140 5664
rect 79192 5652 79198 5704
rect 79410 5624 79416 5636
rect 65076 5596 79416 5624
rect 79410 5584 79416 5596
rect 79468 5584 79474 5636
rect 79520 5633 79548 5800
rect 79870 5788 79876 5840
rect 79928 5828 79934 5840
rect 85945 5831 86003 5837
rect 85945 5828 85957 5831
rect 79928 5800 85957 5828
rect 79928 5788 79934 5800
rect 85945 5797 85957 5800
rect 85991 5797 86003 5831
rect 85945 5791 86003 5797
rect 79594 5720 79600 5772
rect 79652 5760 79658 5772
rect 79689 5763 79747 5769
rect 79689 5760 79701 5763
rect 79652 5732 79701 5760
rect 79652 5720 79658 5732
rect 79689 5729 79701 5732
rect 79735 5729 79747 5763
rect 79689 5723 79747 5729
rect 79778 5720 79784 5772
rect 79836 5760 79842 5772
rect 80333 5763 80391 5769
rect 80333 5760 80345 5763
rect 79836 5732 80345 5760
rect 79836 5720 79842 5732
rect 80333 5729 80345 5732
rect 80379 5729 80391 5763
rect 81710 5760 81716 5772
rect 81671 5732 81716 5760
rect 80333 5723 80391 5729
rect 81710 5720 81716 5732
rect 81768 5720 81774 5772
rect 82814 5720 82820 5772
rect 82872 5760 82878 5772
rect 83185 5763 83243 5769
rect 83185 5760 83197 5763
rect 82872 5732 83197 5760
rect 82872 5720 82878 5732
rect 83185 5729 83197 5732
rect 83231 5729 83243 5763
rect 84470 5760 84476 5772
rect 84431 5732 84476 5760
rect 83185 5723 83243 5729
rect 84470 5720 84476 5732
rect 84528 5720 84534 5772
rect 84930 5720 84936 5772
rect 84988 5760 84994 5772
rect 85117 5763 85175 5769
rect 85117 5760 85129 5763
rect 84988 5732 85129 5760
rect 84988 5720 84994 5732
rect 85117 5729 85129 5732
rect 85163 5729 85175 5763
rect 86034 5760 86040 5772
rect 85995 5732 86040 5760
rect 85117 5723 85175 5729
rect 86034 5720 86040 5732
rect 86092 5720 86098 5772
rect 177945 5763 178003 5769
rect 177945 5729 177957 5763
rect 177991 5760 178003 5763
rect 178678 5760 178684 5772
rect 177991 5732 178684 5760
rect 177991 5729 178003 5732
rect 177945 5723 178003 5729
rect 178678 5720 178684 5732
rect 178736 5720 178742 5772
rect 83093 5695 83151 5701
rect 83093 5692 83105 5695
rect 82096 5664 83105 5692
rect 79505 5627 79563 5633
rect 79505 5593 79517 5627
rect 79551 5593 79563 5627
rect 79505 5587 79563 5593
rect 79594 5584 79600 5636
rect 79652 5624 79658 5636
rect 80149 5627 80207 5633
rect 79652 5596 80100 5624
rect 79652 5584 79658 5596
rect 64782 5556 64788 5568
rect 63696 5528 64788 5556
rect 64782 5516 64788 5528
rect 64840 5516 64846 5568
rect 65242 5516 65248 5568
rect 65300 5556 65306 5568
rect 65705 5559 65763 5565
rect 65705 5556 65717 5559
rect 65300 5528 65717 5556
rect 65300 5516 65306 5528
rect 65705 5525 65717 5528
rect 65751 5525 65763 5559
rect 65705 5519 65763 5525
rect 67818 5516 67824 5568
rect 67876 5556 67882 5568
rect 68833 5559 68891 5565
rect 68833 5556 68845 5559
rect 67876 5528 68845 5556
rect 67876 5516 67882 5528
rect 68833 5525 68845 5528
rect 68879 5525 68891 5559
rect 68833 5519 68891 5525
rect 73065 5559 73123 5565
rect 73065 5525 73077 5559
rect 73111 5556 73123 5559
rect 73798 5556 73804 5568
rect 73111 5528 73804 5556
rect 73111 5525 73123 5528
rect 73065 5519 73123 5525
rect 73798 5516 73804 5528
rect 73856 5516 73862 5568
rect 73893 5559 73951 5565
rect 73893 5525 73905 5559
rect 73939 5556 73951 5559
rect 75178 5556 75184 5568
rect 73939 5528 75184 5556
rect 73939 5525 73951 5528
rect 73893 5519 73951 5525
rect 75178 5516 75184 5528
rect 75236 5516 75242 5568
rect 79045 5559 79103 5565
rect 79045 5525 79057 5559
rect 79091 5556 79103 5559
rect 79962 5556 79968 5568
rect 79091 5528 79968 5556
rect 79091 5525 79103 5528
rect 79045 5519 79103 5525
rect 79962 5516 79968 5528
rect 80020 5516 80026 5568
rect 80072 5556 80100 5596
rect 80149 5593 80161 5627
rect 80195 5624 80207 5627
rect 80238 5624 80244 5636
rect 80195 5596 80244 5624
rect 80195 5593 80207 5596
rect 80149 5587 80207 5593
rect 80238 5584 80244 5596
rect 80296 5584 80302 5636
rect 82096 5624 82124 5664
rect 83093 5661 83105 5664
rect 83139 5661 83151 5695
rect 83093 5655 83151 5661
rect 84013 5695 84071 5701
rect 84013 5661 84025 5695
rect 84059 5692 84071 5695
rect 89990 5692 89996 5704
rect 84059 5664 89996 5692
rect 84059 5661 84071 5664
rect 84013 5655 84071 5661
rect 89990 5652 89996 5664
rect 90048 5652 90054 5704
rect 80808 5596 82124 5624
rect 80808 5556 80836 5596
rect 82170 5584 82176 5636
rect 82228 5624 82234 5636
rect 85301 5627 85359 5633
rect 85301 5624 85313 5627
rect 82228 5596 85313 5624
rect 82228 5584 82234 5596
rect 85301 5593 85313 5596
rect 85347 5593 85359 5627
rect 85301 5587 85359 5593
rect 85945 5627 86003 5633
rect 85945 5593 85957 5627
rect 85991 5624 86003 5627
rect 86221 5627 86279 5633
rect 86221 5624 86233 5627
rect 85991 5596 86233 5624
rect 85991 5593 86003 5596
rect 85945 5587 86003 5593
rect 86221 5593 86233 5596
rect 86267 5593 86279 5627
rect 86221 5587 86279 5593
rect 80072 5528 80836 5556
rect 80882 5516 80888 5568
rect 80940 5556 80946 5568
rect 81253 5559 81311 5565
rect 81253 5556 81265 5559
rect 80940 5528 81265 5556
rect 80940 5516 80946 5528
rect 81253 5525 81265 5528
rect 81299 5525 81311 5559
rect 81253 5519 81311 5525
rect 81897 5559 81955 5565
rect 81897 5525 81909 5559
rect 81943 5556 81955 5559
rect 82446 5556 82452 5568
rect 81943 5528 82452 5556
rect 81943 5525 81955 5528
rect 81897 5519 81955 5525
rect 82446 5516 82452 5528
rect 82504 5516 82510 5568
rect 83369 5559 83427 5565
rect 83369 5525 83381 5559
rect 83415 5556 83427 5559
rect 83550 5556 83556 5568
rect 83415 5528 83556 5556
rect 83415 5525 83427 5528
rect 83369 5519 83427 5525
rect 83550 5516 83556 5528
rect 83608 5516 83614 5568
rect 84657 5559 84715 5565
rect 84657 5525 84669 5559
rect 84703 5556 84715 5559
rect 85114 5556 85120 5568
rect 84703 5528 85120 5556
rect 84703 5525 84715 5528
rect 84657 5519 84715 5525
rect 85114 5516 85120 5528
rect 85172 5516 85178 5568
rect 1104 5466 178848 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 34966 5466
rect 35018 5414 35030 5466
rect 35082 5414 35094 5466
rect 35146 5414 35158 5466
rect 35210 5414 65686 5466
rect 65738 5414 65750 5466
rect 65802 5414 65814 5466
rect 65866 5414 65878 5466
rect 65930 5414 96406 5466
rect 96458 5414 96470 5466
rect 96522 5414 96534 5466
rect 96586 5414 96598 5466
rect 96650 5414 127126 5466
rect 127178 5414 127190 5466
rect 127242 5414 127254 5466
rect 127306 5414 127318 5466
rect 127370 5414 157846 5466
rect 157898 5414 157910 5466
rect 157962 5414 157974 5466
rect 158026 5414 158038 5466
rect 158090 5414 178848 5466
rect 1104 5392 178848 5414
rect 1946 5312 1952 5364
rect 2004 5352 2010 5364
rect 23750 5352 23756 5364
rect 2004 5324 23756 5352
rect 2004 5312 2010 5324
rect 23750 5312 23756 5324
rect 23808 5312 23814 5364
rect 28810 5352 28816 5364
rect 23860 5324 28816 5352
rect 18690 5284 18696 5296
rect 18651 5256 18696 5284
rect 18690 5244 18696 5256
rect 18748 5244 18754 5296
rect 20530 5284 20536 5296
rect 20491 5256 20536 5284
rect 20530 5244 20536 5256
rect 20588 5244 20594 5296
rect 17310 5216 17316 5228
rect 17271 5188 17316 5216
rect 17310 5176 17316 5188
rect 17368 5176 17374 5228
rect 19150 5216 19156 5228
rect 19111 5188 19156 5216
rect 19150 5176 19156 5188
rect 19208 5176 19214 5228
rect 23860 5225 23888 5324
rect 28810 5312 28816 5324
rect 28868 5312 28874 5364
rect 28966 5324 30512 5352
rect 23845 5219 23903 5225
rect 23845 5185 23857 5219
rect 23891 5185 23903 5219
rect 28166 5216 28172 5228
rect 25622 5188 28172 5216
rect 23845 5179 23903 5185
rect 28166 5176 28172 5188
rect 28224 5216 28230 5228
rect 28966 5216 28994 5324
rect 30484 5284 30512 5324
rect 30558 5312 30564 5364
rect 30616 5352 30622 5364
rect 30926 5352 30932 5364
rect 30616 5324 30932 5352
rect 30616 5312 30622 5324
rect 30926 5312 30932 5324
rect 30984 5312 30990 5364
rect 34238 5352 34244 5364
rect 31726 5324 34244 5352
rect 31570 5284 31576 5296
rect 30484 5256 31576 5284
rect 31570 5244 31576 5256
rect 31628 5244 31634 5296
rect 29270 5216 29276 5228
rect 28224 5188 28994 5216
rect 29231 5188 29276 5216
rect 28224 5176 28230 5188
rect 29270 5176 29276 5188
rect 29328 5176 29334 5228
rect 19420 5151 19478 5157
rect 19420 5117 19432 5151
rect 19466 5148 19478 5151
rect 21082 5148 21088 5160
rect 19466 5120 21088 5148
rect 19466 5117 19478 5120
rect 19420 5111 19478 5117
rect 21082 5108 21088 5120
rect 21140 5108 21146 5160
rect 24946 5108 24952 5160
rect 25004 5108 25010 5160
rect 25406 5108 25412 5160
rect 25464 5148 25470 5160
rect 31726 5148 31754 5324
rect 34238 5312 34244 5324
rect 34296 5312 34302 5364
rect 34330 5312 34336 5364
rect 34388 5352 34394 5364
rect 34425 5355 34483 5361
rect 34425 5352 34437 5355
rect 34388 5324 34437 5352
rect 34388 5312 34394 5324
rect 34425 5321 34437 5324
rect 34471 5321 34483 5355
rect 35986 5352 35992 5364
rect 34425 5315 34483 5321
rect 34900 5324 35992 5352
rect 34790 5284 34796 5296
rect 34072 5256 34796 5284
rect 32030 5176 32036 5228
rect 32088 5216 32094 5228
rect 33045 5219 33103 5225
rect 33045 5216 33057 5219
rect 32088 5188 33057 5216
rect 32088 5176 32094 5188
rect 33045 5185 33057 5188
rect 33091 5185 33103 5219
rect 33045 5179 33103 5185
rect 25464 5120 31754 5148
rect 33060 5148 33088 5179
rect 33312 5151 33370 5157
rect 33060 5120 33272 5148
rect 25464 5108 25470 5120
rect 17580 5083 17638 5089
rect 17580 5049 17592 5083
rect 17626 5080 17638 5083
rect 21542 5080 21548 5092
rect 17626 5052 21548 5080
rect 17626 5049 17638 5052
rect 17580 5043 17638 5049
rect 21542 5040 21548 5052
rect 21600 5040 21606 5092
rect 27982 5040 27988 5092
rect 28040 5080 28046 5092
rect 29540 5083 29598 5089
rect 28040 5052 29500 5080
rect 28040 5040 28046 5052
rect 15654 4972 15660 5024
rect 15712 5012 15718 5024
rect 20530 5012 20536 5024
rect 15712 4984 20536 5012
rect 15712 4972 15718 4984
rect 20530 4972 20536 4984
rect 20588 4972 20594 5024
rect 24857 5015 24915 5021
rect 24857 4981 24869 5015
rect 24903 5012 24915 5015
rect 28350 5012 28356 5024
rect 24903 4984 28356 5012
rect 24903 4981 24915 4984
rect 24857 4975 24915 4981
rect 28350 4972 28356 4984
rect 28408 4972 28414 5024
rect 29472 5012 29500 5052
rect 29540 5049 29552 5083
rect 29586 5080 29598 5083
rect 33134 5080 33140 5092
rect 29586 5052 33140 5080
rect 29586 5049 29598 5052
rect 29540 5043 29598 5049
rect 33134 5040 33140 5052
rect 33192 5040 33198 5092
rect 33244 5080 33272 5120
rect 33312 5117 33324 5151
rect 33358 5148 33370 5151
rect 34072 5148 34100 5256
rect 34790 5244 34796 5256
rect 34848 5244 34854 5296
rect 34900 5225 34928 5324
rect 35986 5312 35992 5324
rect 36044 5312 36050 5364
rect 36078 5312 36084 5364
rect 36136 5352 36142 5364
rect 36136 5324 37504 5352
rect 36136 5312 36142 5324
rect 37274 5284 37280 5296
rect 35912 5256 37280 5284
rect 34885 5219 34943 5225
rect 34885 5216 34897 5219
rect 33358 5120 34100 5148
rect 34164 5188 34897 5216
rect 33358 5117 33370 5120
rect 33312 5111 33370 5117
rect 34164 5080 34192 5188
rect 34885 5185 34897 5188
rect 34931 5185 34943 5219
rect 34885 5179 34943 5185
rect 35152 5151 35210 5157
rect 35152 5117 35164 5151
rect 35198 5148 35210 5151
rect 35912 5148 35940 5256
rect 37274 5244 37280 5256
rect 37332 5244 37338 5296
rect 37476 5216 37504 5324
rect 38286 5312 38292 5364
rect 38344 5352 38350 5364
rect 38344 5324 41414 5352
rect 38344 5312 38350 5324
rect 39669 5287 39727 5293
rect 39669 5253 39681 5287
rect 39715 5284 39727 5287
rect 39850 5284 39856 5296
rect 39715 5256 39856 5284
rect 39715 5253 39727 5256
rect 39669 5247 39727 5253
rect 39850 5244 39856 5256
rect 39908 5244 39914 5296
rect 39960 5216 39988 5324
rect 41386 5284 41414 5324
rect 41506 5312 41512 5364
rect 41564 5352 41570 5364
rect 42150 5352 42156 5364
rect 41564 5324 42156 5352
rect 41564 5312 41570 5324
rect 42150 5312 42156 5324
rect 42208 5312 42214 5364
rect 42429 5355 42487 5361
rect 42429 5321 42441 5355
rect 42475 5352 42487 5355
rect 42475 5324 46704 5352
rect 42475 5321 42487 5324
rect 42429 5315 42487 5321
rect 41874 5284 41880 5296
rect 41386 5256 41880 5284
rect 41874 5244 41880 5256
rect 41932 5284 41938 5296
rect 43530 5284 43536 5296
rect 41932 5256 43536 5284
rect 41932 5244 41938 5256
rect 43530 5244 43536 5256
rect 43588 5244 43594 5296
rect 46676 5284 46704 5324
rect 46750 5312 46756 5364
rect 46808 5352 46814 5364
rect 47670 5352 47676 5364
rect 46808 5324 47676 5352
rect 46808 5312 46814 5324
rect 47670 5312 47676 5324
rect 47728 5352 47734 5364
rect 63129 5355 63187 5361
rect 47728 5324 63080 5352
rect 47728 5312 47734 5324
rect 47210 5284 47216 5296
rect 46676 5256 47216 5284
rect 47210 5244 47216 5256
rect 47268 5244 47274 5296
rect 63052 5284 63080 5324
rect 63129 5321 63141 5355
rect 63175 5352 63187 5355
rect 63218 5352 63224 5364
rect 63175 5324 63224 5352
rect 63175 5321 63187 5324
rect 63129 5315 63187 5321
rect 63218 5312 63224 5324
rect 63276 5312 63282 5364
rect 69201 5355 69259 5361
rect 69201 5352 69213 5355
rect 63328 5324 69213 5352
rect 63328 5284 63356 5324
rect 69201 5321 69213 5324
rect 69247 5321 69259 5355
rect 69201 5315 69259 5321
rect 72050 5312 72056 5364
rect 72108 5352 72114 5364
rect 76558 5352 76564 5364
rect 72108 5324 76564 5352
rect 72108 5312 72114 5324
rect 76558 5312 76564 5324
rect 76616 5312 76622 5364
rect 78217 5355 78275 5361
rect 78217 5321 78229 5355
rect 78263 5352 78275 5355
rect 78766 5352 78772 5364
rect 78263 5324 78772 5352
rect 78263 5321 78275 5324
rect 78217 5315 78275 5321
rect 78766 5312 78772 5324
rect 78824 5312 78830 5364
rect 78861 5355 78919 5361
rect 78861 5321 78873 5355
rect 78907 5352 78919 5355
rect 81802 5352 81808 5364
rect 78907 5324 81808 5352
rect 78907 5321 78919 5324
rect 78861 5315 78919 5321
rect 81802 5312 81808 5324
rect 81860 5312 81866 5364
rect 82265 5355 82323 5361
rect 82265 5321 82277 5355
rect 82311 5352 82323 5355
rect 82446 5352 82452 5364
rect 82311 5324 82452 5352
rect 82311 5321 82323 5324
rect 82265 5315 82323 5321
rect 82446 5312 82452 5324
rect 82504 5352 82510 5364
rect 84654 5352 84660 5364
rect 82504 5324 84660 5352
rect 82504 5312 82510 5324
rect 84654 5312 84660 5324
rect 84712 5312 84718 5364
rect 84746 5312 84752 5364
rect 84804 5352 84810 5364
rect 88978 5352 88984 5364
rect 84804 5324 88984 5352
rect 84804 5312 84810 5324
rect 88978 5312 88984 5324
rect 89036 5312 89042 5364
rect 94406 5352 94412 5364
rect 89686 5324 94412 5352
rect 82081 5287 82139 5293
rect 82081 5284 82093 5287
rect 61304 5256 62068 5284
rect 63052 5256 63356 5284
rect 63420 5256 82093 5284
rect 40129 5219 40187 5225
rect 40129 5216 40141 5219
rect 35198 5120 35940 5148
rect 36004 5188 37412 5216
rect 37476 5188 38424 5216
rect 39960 5188 40141 5216
rect 35198 5117 35210 5120
rect 35152 5111 35210 5117
rect 33244 5052 34192 5080
rect 34514 5040 34520 5092
rect 34572 5080 34578 5092
rect 36004 5080 36032 5188
rect 37384 5157 37412 5188
rect 37369 5151 37427 5157
rect 37369 5117 37381 5151
rect 37415 5117 37427 5151
rect 38286 5148 38292 5160
rect 38247 5120 38292 5148
rect 37369 5111 37427 5117
rect 38286 5108 38292 5120
rect 38344 5108 38350 5160
rect 38396 5148 38424 5188
rect 40129 5185 40141 5188
rect 40175 5185 40187 5219
rect 40129 5179 40187 5185
rect 44818 5176 44824 5228
rect 44876 5216 44882 5228
rect 45278 5216 45284 5228
rect 44876 5188 45284 5216
rect 44876 5176 44882 5188
rect 45278 5176 45284 5188
rect 45336 5216 45342 5228
rect 45373 5219 45431 5225
rect 45373 5216 45385 5219
rect 45336 5188 45385 5216
rect 45336 5176 45342 5188
rect 45373 5185 45385 5188
rect 45419 5185 45431 5219
rect 45373 5179 45431 5185
rect 46382 5176 46388 5228
rect 46440 5216 46446 5228
rect 47762 5216 47768 5228
rect 46440 5188 47768 5216
rect 46440 5176 46446 5188
rect 47762 5176 47768 5188
rect 47820 5176 47826 5228
rect 61304 5225 61332 5256
rect 61289 5219 61347 5225
rect 61289 5185 61301 5219
rect 61335 5185 61347 5219
rect 61289 5179 61347 5185
rect 61473 5219 61531 5225
rect 61473 5185 61485 5219
rect 61519 5216 61531 5219
rect 61654 5216 61660 5228
rect 61519 5188 61660 5216
rect 61519 5185 61531 5188
rect 61473 5179 61531 5185
rect 61654 5176 61660 5188
rect 61712 5176 61718 5228
rect 61930 5216 61936 5228
rect 61891 5188 61936 5216
rect 61930 5176 61936 5188
rect 61988 5176 61994 5228
rect 62040 5216 62068 5256
rect 62390 5225 62396 5228
rect 62347 5219 62396 5225
rect 62347 5216 62359 5219
rect 62040 5188 62359 5216
rect 62347 5185 62359 5188
rect 62393 5185 62396 5219
rect 62347 5179 62396 5185
rect 62390 5176 62396 5179
rect 62448 5176 62454 5228
rect 42613 5151 42671 5157
rect 42613 5148 42625 5151
rect 38396 5120 42625 5148
rect 42613 5117 42625 5120
rect 42659 5117 42671 5151
rect 43530 5148 43536 5160
rect 43491 5120 43536 5148
rect 42613 5111 42671 5117
rect 43530 5108 43536 5120
rect 43588 5108 43594 5160
rect 44174 5148 44180 5160
rect 43640 5120 44180 5148
rect 38378 5080 38384 5092
rect 34572 5052 36032 5080
rect 36096 5052 38384 5080
rect 34572 5040 34578 5052
rect 30466 5012 30472 5024
rect 29472 4984 30472 5012
rect 30466 4972 30472 4984
rect 30524 4972 30530 5024
rect 30558 4972 30564 5024
rect 30616 5012 30622 5024
rect 30653 5015 30711 5021
rect 30653 5012 30665 5015
rect 30616 4984 30665 5012
rect 30616 4972 30622 4984
rect 30653 4981 30665 4984
rect 30699 4981 30711 5015
rect 30653 4975 30711 4981
rect 30742 4972 30748 5024
rect 30800 5012 30806 5024
rect 31754 5012 31760 5024
rect 30800 4984 31760 5012
rect 30800 4972 30806 4984
rect 31754 4972 31760 4984
rect 31812 4972 31818 5024
rect 31846 4972 31852 5024
rect 31904 5012 31910 5024
rect 36096 5012 36124 5052
rect 38378 5040 38384 5052
rect 38436 5040 38442 5092
rect 38470 5040 38476 5092
rect 38528 5089 38534 5092
rect 38528 5083 38592 5089
rect 38528 5049 38546 5083
rect 38580 5049 38592 5083
rect 38528 5043 38592 5049
rect 38528 5040 38534 5043
rect 38654 5040 38660 5092
rect 38712 5080 38718 5092
rect 39206 5080 39212 5092
rect 38712 5052 39212 5080
rect 38712 5040 38718 5052
rect 39206 5040 39212 5052
rect 39264 5040 39270 5092
rect 39942 5080 39948 5092
rect 39592 5052 39948 5080
rect 36262 5012 36268 5024
rect 31904 4984 36124 5012
rect 36223 4984 36268 5012
rect 31904 4972 31910 4984
rect 36262 4972 36268 4984
rect 36320 5012 36326 5024
rect 37090 5012 37096 5024
rect 36320 4984 37096 5012
rect 36320 4972 36326 4984
rect 37090 4972 37096 4984
rect 37148 4972 37154 5024
rect 37185 5015 37243 5021
rect 37185 4981 37197 5015
rect 37231 5012 37243 5015
rect 39592 5012 39620 5052
rect 39942 5040 39948 5052
rect 40000 5040 40006 5092
rect 40396 5083 40454 5089
rect 40396 5049 40408 5083
rect 40442 5080 40454 5083
rect 43640 5080 43668 5120
rect 44174 5108 44180 5120
rect 44232 5108 44238 5160
rect 47026 5148 47032 5160
rect 45388 5120 47032 5148
rect 40442 5052 43668 5080
rect 43800 5083 43858 5089
rect 40442 5049 40454 5052
rect 40396 5043 40454 5049
rect 43800 5049 43812 5083
rect 43846 5080 43858 5083
rect 45388 5080 45416 5120
rect 47026 5108 47032 5120
rect 47084 5108 47090 5160
rect 47394 5108 47400 5160
rect 47452 5148 47458 5160
rect 47452 5120 47497 5148
rect 47452 5108 47458 5120
rect 62206 5108 62212 5160
rect 62264 5148 62270 5160
rect 62482 5148 62488 5160
rect 62264 5120 62309 5148
rect 62443 5120 62488 5148
rect 62264 5108 62270 5120
rect 62482 5108 62488 5120
rect 62540 5108 62546 5160
rect 43846 5052 45416 5080
rect 45640 5083 45698 5089
rect 43846 5049 43858 5052
rect 43800 5043 43858 5049
rect 45640 5049 45652 5083
rect 45686 5080 45698 5083
rect 50614 5080 50620 5092
rect 45686 5052 50620 5080
rect 45686 5049 45698 5052
rect 45640 5043 45698 5049
rect 50614 5040 50620 5052
rect 50672 5040 50678 5092
rect 37231 4984 39620 5012
rect 37231 4981 37243 4984
rect 37185 4975 37243 4981
rect 40034 4972 40040 5024
rect 40092 5012 40098 5024
rect 41506 5012 41512 5024
rect 40092 4984 41512 5012
rect 40092 4972 40098 4984
rect 41506 4972 41512 4984
rect 41564 4972 41570 5024
rect 43990 4972 43996 5024
rect 44048 5012 44054 5024
rect 44913 5015 44971 5021
rect 44913 5012 44925 5015
rect 44048 4984 44925 5012
rect 44048 4972 44054 4984
rect 44913 4981 44925 4984
rect 44959 5012 44971 5015
rect 45370 5012 45376 5024
rect 44959 4984 45376 5012
rect 44959 4981 44971 4984
rect 44913 4975 44971 4981
rect 45370 4972 45376 4984
rect 45428 4972 45434 5024
rect 45462 4972 45468 5024
rect 45520 5012 45526 5024
rect 46382 5012 46388 5024
rect 45520 4984 46388 5012
rect 45520 4972 45526 4984
rect 46382 4972 46388 4984
rect 46440 4972 46446 5024
rect 46474 4972 46480 5024
rect 46532 5012 46538 5024
rect 46753 5015 46811 5021
rect 46753 5012 46765 5015
rect 46532 4984 46765 5012
rect 46532 4972 46538 4984
rect 46753 4981 46765 4984
rect 46799 5012 46811 5015
rect 47026 5012 47032 5024
rect 46799 4984 47032 5012
rect 46799 4981 46811 4984
rect 46753 4975 46811 4981
rect 47026 4972 47032 4984
rect 47084 4972 47090 5024
rect 47213 5015 47271 5021
rect 47213 4981 47225 5015
rect 47259 5012 47271 5015
rect 49878 5012 49884 5024
rect 47259 4984 49884 5012
rect 47259 4981 47271 4984
rect 47213 4975 47271 4981
rect 49878 4972 49884 4984
rect 49936 4972 49942 5024
rect 60458 4972 60464 5024
rect 60516 5012 60522 5024
rect 63420 5012 63448 5256
rect 82081 5253 82093 5256
rect 82127 5253 82139 5287
rect 86957 5287 87015 5293
rect 86957 5284 86969 5287
rect 82081 5247 82139 5253
rect 82188 5256 86969 5284
rect 64782 5176 64788 5228
rect 64840 5216 64846 5228
rect 78214 5216 78220 5228
rect 64840 5188 77984 5216
rect 64840 5176 64846 5188
rect 63862 5108 63868 5160
rect 63920 5148 63926 5160
rect 64693 5151 64751 5157
rect 64693 5148 64705 5151
rect 63920 5120 64705 5148
rect 63920 5108 63926 5120
rect 64693 5117 64705 5120
rect 64739 5117 64751 5151
rect 64693 5111 64751 5117
rect 75825 5151 75883 5157
rect 75825 5117 75837 5151
rect 75871 5148 75883 5151
rect 76098 5148 76104 5160
rect 75871 5120 76104 5148
rect 75871 5117 75883 5120
rect 75825 5111 75883 5117
rect 76098 5108 76104 5120
rect 76156 5108 76162 5160
rect 76466 5108 76472 5160
rect 76524 5148 76530 5160
rect 76653 5151 76711 5157
rect 76653 5148 76665 5151
rect 76524 5120 76665 5148
rect 76524 5108 76530 5120
rect 76653 5117 76665 5120
rect 76699 5117 76711 5151
rect 77570 5148 77576 5160
rect 77531 5120 77576 5148
rect 76653 5111 76711 5117
rect 77570 5108 77576 5120
rect 77628 5108 77634 5160
rect 71958 5040 71964 5092
rect 72016 5080 72022 5092
rect 72016 5052 76512 5080
rect 72016 5040 72022 5052
rect 60516 4984 63448 5012
rect 60516 4972 60522 4984
rect 63494 4972 63500 5024
rect 63552 5012 63558 5024
rect 64509 5015 64567 5021
rect 64509 5012 64521 5015
rect 63552 4984 64521 5012
rect 63552 4972 63558 4984
rect 64509 4981 64521 4984
rect 64555 4981 64567 5015
rect 64509 4975 64567 4981
rect 69201 5015 69259 5021
rect 69201 4981 69213 5015
rect 69247 5012 69259 5015
rect 75914 5012 75920 5024
rect 69247 4984 75920 5012
rect 69247 4981 69259 4984
rect 69201 4975 69259 4981
rect 75914 4972 75920 4984
rect 75972 4972 75978 5024
rect 76009 5015 76067 5021
rect 76009 4981 76021 5015
rect 76055 5012 76067 5015
rect 76374 5012 76380 5024
rect 76055 4984 76380 5012
rect 76055 4981 76067 4984
rect 76009 4975 76067 4981
rect 76374 4972 76380 4984
rect 76432 4972 76438 5024
rect 76484 5021 76512 5052
rect 76469 5015 76527 5021
rect 76469 4981 76481 5015
rect 76515 4981 76527 5015
rect 77956 5012 77984 5188
rect 78048 5188 78220 5216
rect 78048 5157 78076 5188
rect 78214 5176 78220 5188
rect 78272 5176 78278 5228
rect 78766 5176 78772 5228
rect 78824 5216 78830 5228
rect 78824 5188 80652 5216
rect 78824 5176 78830 5188
rect 78033 5151 78091 5157
rect 78033 5117 78045 5151
rect 78079 5117 78091 5151
rect 78033 5111 78091 5117
rect 78122 5108 78128 5160
rect 78180 5148 78186 5160
rect 78677 5151 78735 5157
rect 78677 5148 78689 5151
rect 78180 5120 78689 5148
rect 78180 5108 78186 5120
rect 78677 5117 78689 5120
rect 78723 5117 78735 5151
rect 78677 5111 78735 5117
rect 80238 5108 80244 5160
rect 80296 5148 80302 5160
rect 80425 5151 80483 5157
rect 80425 5148 80437 5151
rect 80296 5120 80437 5148
rect 80296 5108 80302 5120
rect 80425 5117 80437 5120
rect 80471 5117 80483 5151
rect 80425 5111 80483 5117
rect 80624 5148 80652 5188
rect 80698 5176 80704 5228
rect 80756 5216 80762 5228
rect 82188 5216 82216 5256
rect 86957 5253 86969 5256
rect 87003 5253 87015 5287
rect 86957 5247 87015 5253
rect 82630 5216 82636 5228
rect 80756 5188 82216 5216
rect 82543 5188 82636 5216
rect 80756 5176 80762 5188
rect 82630 5176 82636 5188
rect 82688 5216 82694 5228
rect 85669 5219 85727 5225
rect 82688 5188 84240 5216
rect 82688 5176 82694 5188
rect 81437 5151 81495 5157
rect 81437 5148 81449 5151
rect 80624 5120 81449 5148
rect 79318 5012 79324 5024
rect 77956 4984 79324 5012
rect 76469 4975 76527 4981
rect 79318 4972 79324 4984
rect 79376 4972 79382 5024
rect 80330 4972 80336 5024
rect 80388 5012 80394 5024
rect 80624 5012 80652 5120
rect 81437 5117 81449 5120
rect 81483 5148 81495 5151
rect 82814 5148 82820 5160
rect 81483 5120 82820 5148
rect 81483 5117 81495 5120
rect 81437 5111 81495 5117
rect 82814 5108 82820 5120
rect 82872 5108 82878 5160
rect 83093 5151 83151 5157
rect 83093 5117 83105 5151
rect 83139 5148 83151 5151
rect 83366 5148 83372 5160
rect 83139 5120 83372 5148
rect 83139 5117 83151 5120
rect 83093 5111 83151 5117
rect 83366 5108 83372 5120
rect 83424 5108 83430 5160
rect 83458 5108 83464 5160
rect 83516 5148 83522 5160
rect 84105 5151 84163 5157
rect 83516 5120 83561 5148
rect 83516 5108 83522 5120
rect 84105 5117 84117 5151
rect 84151 5117 84163 5151
rect 84105 5111 84163 5117
rect 81989 5083 82047 5089
rect 81989 5049 82001 5083
rect 82035 5080 82047 5083
rect 82262 5080 82268 5092
rect 82035 5052 82268 5080
rect 82035 5049 82047 5052
rect 81989 5043 82047 5049
rect 82262 5040 82268 5052
rect 82320 5040 82326 5092
rect 82832 5080 82860 5108
rect 84120 5080 84148 5111
rect 82832 5052 84148 5080
rect 84212 5080 84240 5188
rect 85669 5185 85681 5219
rect 85715 5216 85727 5219
rect 86218 5216 86224 5228
rect 85715 5188 86224 5216
rect 85715 5185 85727 5188
rect 85669 5179 85727 5185
rect 86218 5176 86224 5188
rect 86276 5176 86282 5228
rect 89686 5216 89714 5324
rect 94406 5312 94412 5324
rect 94464 5312 94470 5364
rect 86328 5188 89714 5216
rect 85574 5108 85580 5160
rect 85632 5148 85638 5160
rect 86129 5151 86187 5157
rect 86129 5148 86141 5151
rect 85632 5120 86141 5148
rect 85632 5108 85638 5120
rect 86129 5117 86141 5120
rect 86175 5117 86187 5151
rect 86129 5111 86187 5117
rect 86328 5080 86356 5188
rect 86770 5148 86776 5160
rect 86731 5120 86776 5148
rect 86770 5108 86776 5120
rect 86828 5108 86834 5160
rect 87138 5108 87144 5160
rect 87196 5148 87202 5160
rect 87417 5151 87475 5157
rect 87417 5148 87429 5151
rect 87196 5120 87429 5148
rect 87196 5108 87202 5120
rect 87417 5117 87429 5120
rect 87463 5117 87475 5151
rect 87417 5111 87475 5117
rect 177301 5151 177359 5157
rect 177301 5117 177313 5151
rect 177347 5148 177359 5151
rect 177574 5148 177580 5160
rect 177347 5120 177580 5148
rect 177347 5117 177359 5120
rect 177301 5111 177359 5117
rect 177574 5108 177580 5120
rect 177632 5108 177638 5160
rect 177945 5151 178003 5157
rect 177945 5117 177957 5151
rect 177991 5148 178003 5151
rect 179046 5148 179052 5160
rect 177991 5120 179052 5148
rect 177991 5117 178003 5120
rect 177945 5111 178003 5117
rect 179046 5108 179052 5120
rect 179104 5108 179110 5160
rect 84212 5052 86356 5080
rect 86678 5040 86684 5092
rect 86736 5080 86742 5092
rect 86736 5052 89714 5080
rect 86736 5040 86742 5052
rect 80388 4984 80652 5012
rect 80388 4972 80394 4984
rect 81526 4972 81532 5024
rect 81584 5012 81590 5024
rect 81621 5015 81679 5021
rect 81621 5012 81633 5015
rect 81584 4984 81633 5012
rect 81584 4972 81590 4984
rect 81621 4981 81633 4984
rect 81667 4981 81679 5015
rect 83274 5012 83280 5024
rect 83235 4984 83280 5012
rect 81621 4975 81679 4981
rect 83274 4972 83280 4984
rect 83332 4972 83338 5024
rect 83366 4972 83372 5024
rect 83424 5012 83430 5024
rect 83642 5012 83648 5024
rect 83424 4984 83469 5012
rect 83603 4984 83648 5012
rect 83424 4972 83430 4984
rect 83642 4972 83648 4984
rect 83700 4972 83706 5024
rect 84286 5012 84292 5024
rect 84247 4984 84292 5012
rect 84286 4972 84292 4984
rect 84344 4972 84350 5024
rect 86218 4972 86224 5024
rect 86276 5012 86282 5024
rect 86313 5015 86371 5021
rect 86313 5012 86325 5015
rect 86276 4984 86325 5012
rect 86276 4972 86282 4984
rect 86313 4981 86325 4984
rect 86359 4981 86371 5015
rect 86313 4975 86371 4981
rect 86494 4972 86500 5024
rect 86552 5012 86558 5024
rect 87601 5015 87659 5021
rect 87601 5012 87613 5015
rect 86552 4984 87613 5012
rect 86552 4972 86558 4984
rect 87601 4981 87613 4984
rect 87647 4981 87659 5015
rect 89686 5012 89714 5052
rect 102778 5012 102784 5024
rect 89686 4984 102784 5012
rect 87601 4975 87659 4981
rect 102778 4972 102784 4984
rect 102836 4972 102842 5024
rect 1104 4922 178848 4944
rect 1104 4870 19606 4922
rect 19658 4870 19670 4922
rect 19722 4870 19734 4922
rect 19786 4870 19798 4922
rect 19850 4870 50326 4922
rect 50378 4870 50390 4922
rect 50442 4870 50454 4922
rect 50506 4870 50518 4922
rect 50570 4870 81046 4922
rect 81098 4870 81110 4922
rect 81162 4870 81174 4922
rect 81226 4870 81238 4922
rect 81290 4870 111766 4922
rect 111818 4870 111830 4922
rect 111882 4870 111894 4922
rect 111946 4870 111958 4922
rect 112010 4870 142486 4922
rect 142538 4870 142550 4922
rect 142602 4870 142614 4922
rect 142666 4870 142678 4922
rect 142730 4870 173206 4922
rect 173258 4870 173270 4922
rect 173322 4870 173334 4922
rect 173386 4870 173398 4922
rect 173450 4870 178848 4922
rect 1104 4848 178848 4870
rect 20070 4768 20076 4820
rect 20128 4808 20134 4820
rect 26602 4808 26608 4820
rect 20128 4780 26608 4808
rect 20128 4768 20134 4780
rect 26602 4768 26608 4780
rect 26660 4768 26666 4820
rect 28350 4808 28356 4820
rect 28311 4780 28356 4808
rect 28350 4768 28356 4780
rect 28408 4808 28414 4820
rect 33413 4811 33471 4817
rect 33413 4808 33425 4811
rect 28408 4780 33425 4808
rect 28408 4768 28414 4780
rect 33413 4777 33425 4780
rect 33459 4808 33471 4811
rect 36998 4808 37004 4820
rect 33459 4780 37004 4808
rect 33459 4777 33471 4780
rect 33413 4771 33471 4777
rect 36998 4768 37004 4780
rect 37056 4768 37062 4820
rect 37274 4768 37280 4820
rect 37332 4808 37338 4820
rect 37332 4780 38424 4808
rect 37332 4768 37338 4780
rect 23750 4700 23756 4752
rect 23808 4740 23814 4752
rect 27982 4740 27988 4752
rect 23808 4712 27988 4740
rect 23808 4700 23814 4712
rect 27982 4700 27988 4712
rect 28040 4700 28046 4752
rect 35989 4743 36047 4749
rect 35989 4709 36001 4743
rect 36035 4740 36047 4743
rect 36630 4740 36636 4752
rect 36035 4712 36636 4740
rect 36035 4709 36047 4712
rect 35989 4703 36047 4709
rect 36630 4700 36636 4712
rect 36688 4700 36694 4752
rect 11790 4672 11796 4684
rect 11751 4644 11796 4672
rect 11790 4632 11796 4644
rect 11848 4632 11854 4684
rect 21542 4632 21548 4684
rect 21600 4672 21606 4684
rect 27890 4672 27896 4684
rect 21600 4644 27896 4672
rect 21600 4632 21606 4644
rect 27890 4632 27896 4644
rect 27948 4632 27954 4684
rect 28074 4632 28080 4684
rect 28132 4632 28138 4684
rect 28902 4632 28908 4684
rect 28960 4672 28966 4684
rect 28960 4644 33166 4672
rect 28960 4632 28966 4644
rect 34238 4632 34244 4684
rect 34296 4672 34302 4684
rect 38197 4675 38255 4681
rect 38197 4672 38209 4675
rect 34296 4644 36754 4672
rect 38028 4644 38209 4672
rect 34296 4632 34302 4644
rect 27341 4607 27399 4613
rect 27341 4573 27353 4607
rect 27387 4604 27399 4607
rect 27387 4576 27660 4604
rect 27387 4573 27399 4576
rect 27341 4567 27399 4573
rect 14274 4496 14280 4548
rect 14332 4536 14338 4548
rect 21910 4536 21916 4548
rect 14332 4508 21916 4536
rect 14332 4496 14338 4508
rect 21910 4496 21916 4508
rect 21968 4496 21974 4548
rect 27632 4536 27660 4576
rect 28166 4564 28172 4616
rect 28224 4604 28230 4616
rect 28224 4576 28382 4604
rect 28224 4564 28230 4576
rect 30466 4564 30472 4616
rect 30524 4604 30530 4616
rect 31662 4604 31668 4616
rect 30524 4576 31668 4604
rect 30524 4564 30530 4576
rect 31662 4564 31668 4576
rect 31720 4564 31726 4616
rect 32398 4604 32404 4616
rect 32359 4576 32404 4604
rect 32398 4564 32404 4576
rect 32456 4564 32462 4616
rect 33778 4564 33784 4616
rect 33836 4564 33842 4616
rect 36633 4607 36691 4613
rect 36633 4604 36645 4607
rect 34440 4576 36645 4604
rect 30742 4536 30748 4548
rect 27632 4508 30748 4536
rect 30742 4496 30748 4508
rect 30800 4496 30806 4548
rect 33134 4496 33140 4548
rect 33192 4536 33198 4548
rect 33686 4536 33692 4548
rect 33192 4508 33692 4536
rect 33192 4496 33198 4508
rect 33686 4496 33692 4508
rect 33744 4496 33750 4548
rect 33796 4536 33824 4564
rect 34440 4536 34468 4576
rect 36633 4573 36645 4576
rect 36679 4604 36691 4607
rect 36906 4604 36912 4616
rect 36679 4576 36912 4604
rect 36679 4573 36691 4576
rect 36633 4567 36691 4573
rect 36906 4564 36912 4576
rect 36964 4564 36970 4616
rect 33796 4508 34468 4536
rect 36078 4496 36084 4548
rect 36136 4536 36142 4548
rect 37182 4536 37188 4548
rect 36136 4508 37188 4536
rect 36136 4496 36142 4508
rect 37182 4496 37188 4508
rect 37240 4536 37246 4548
rect 38028 4536 38056 4644
rect 38197 4641 38209 4644
rect 38243 4672 38255 4675
rect 38286 4672 38292 4684
rect 38243 4644 38292 4672
rect 38243 4641 38255 4644
rect 38197 4635 38255 4641
rect 38286 4632 38292 4644
rect 38344 4632 38350 4684
rect 38396 4672 38424 4780
rect 38654 4768 38660 4820
rect 38712 4808 38718 4820
rect 39577 4811 39635 4817
rect 39577 4808 39589 4811
rect 38712 4780 39589 4808
rect 38712 4768 38718 4780
rect 39577 4777 39589 4780
rect 39623 4808 39635 4811
rect 41966 4808 41972 4820
rect 39623 4780 41972 4808
rect 39623 4777 39635 4780
rect 39577 4771 39635 4777
rect 41966 4768 41972 4780
rect 42024 4768 42030 4820
rect 45189 4811 45247 4817
rect 45189 4777 45201 4811
rect 45235 4808 45247 4811
rect 45462 4808 45468 4820
rect 45235 4780 45468 4808
rect 45235 4777 45247 4780
rect 45189 4771 45247 4777
rect 45462 4768 45468 4780
rect 45520 4768 45526 4820
rect 48130 4808 48136 4820
rect 46032 4780 48136 4808
rect 38464 4743 38522 4749
rect 38464 4709 38476 4743
rect 38510 4740 38522 4743
rect 40218 4740 40224 4752
rect 38510 4712 40224 4740
rect 38510 4709 38522 4712
rect 38464 4703 38522 4709
rect 40218 4700 40224 4712
rect 40276 4700 40282 4752
rect 44076 4743 44134 4749
rect 44076 4709 44088 4743
rect 44122 4740 44134 4743
rect 46032 4740 46060 4780
rect 48130 4768 48136 4780
rect 48188 4768 48194 4820
rect 73890 4768 73896 4820
rect 73948 4808 73954 4820
rect 79321 4811 79379 4817
rect 79321 4808 79333 4811
rect 73948 4780 79333 4808
rect 73948 4768 73954 4780
rect 79321 4777 79333 4780
rect 79367 4777 79379 4811
rect 79321 4771 79379 4777
rect 81434 4768 81440 4820
rect 81492 4808 81498 4820
rect 83921 4811 83979 4817
rect 83921 4808 83933 4811
rect 81492 4780 83933 4808
rect 81492 4768 81498 4780
rect 83921 4777 83933 4780
rect 83967 4777 83979 4811
rect 83921 4771 83979 4777
rect 84102 4768 84108 4820
rect 84160 4808 84166 4820
rect 89625 4811 89683 4817
rect 89625 4808 89637 4811
rect 84160 4780 89637 4808
rect 84160 4768 84166 4780
rect 89625 4777 89637 4780
rect 89671 4777 89683 4811
rect 102778 4808 102784 4820
rect 102739 4780 102784 4808
rect 89625 4771 89683 4777
rect 102778 4768 102784 4780
rect 102836 4768 102842 4820
rect 44122 4712 46060 4740
rect 44122 4709 44134 4712
rect 44076 4703 44134 4709
rect 46106 4700 46112 4752
rect 46164 4740 46170 4752
rect 52178 4740 52184 4752
rect 46164 4712 52184 4740
rect 46164 4700 46170 4712
rect 52178 4700 52184 4712
rect 52236 4700 52242 4752
rect 53926 4700 53932 4752
rect 53984 4740 53990 4752
rect 53984 4712 77524 4740
rect 53984 4700 53990 4712
rect 39758 4672 39764 4684
rect 38396 4644 39764 4672
rect 39758 4632 39764 4644
rect 39816 4632 39822 4684
rect 43530 4632 43536 4684
rect 43588 4672 43594 4684
rect 43809 4675 43867 4681
rect 43809 4672 43821 4675
rect 43588 4644 43821 4672
rect 43588 4632 43594 4644
rect 43809 4641 43821 4644
rect 43855 4672 43867 4675
rect 43855 4644 45324 4672
rect 43855 4641 43867 4644
rect 43809 4635 43867 4641
rect 45296 4616 45324 4644
rect 45370 4632 45376 4684
rect 45428 4672 45434 4684
rect 46290 4672 46296 4684
rect 45428 4644 46296 4672
rect 45428 4632 45434 4644
rect 46290 4632 46296 4644
rect 46348 4632 46354 4684
rect 46468 4675 46526 4681
rect 46468 4641 46480 4675
rect 46514 4672 46526 4675
rect 46934 4672 46940 4684
rect 46514 4644 46940 4672
rect 46514 4641 46526 4644
rect 46468 4635 46526 4641
rect 46934 4632 46940 4644
rect 46992 4632 46998 4684
rect 47026 4632 47032 4684
rect 47084 4672 47090 4684
rect 49602 4672 49608 4684
rect 47084 4644 49608 4672
rect 47084 4632 47090 4644
rect 49602 4632 49608 4644
rect 49660 4632 49666 4684
rect 70578 4672 70584 4684
rect 70539 4644 70584 4672
rect 70578 4632 70584 4644
rect 70636 4632 70642 4684
rect 71774 4632 71780 4684
rect 71832 4672 71838 4684
rect 72421 4675 72479 4681
rect 72421 4672 72433 4675
rect 71832 4644 72433 4672
rect 71832 4632 71838 4644
rect 72421 4641 72433 4644
rect 72467 4641 72479 4675
rect 72421 4635 72479 4641
rect 72786 4632 72792 4684
rect 72844 4672 72850 4684
rect 73065 4675 73123 4681
rect 73065 4672 73077 4675
rect 72844 4644 73077 4672
rect 72844 4632 72850 4644
rect 73065 4641 73077 4644
rect 73111 4641 73123 4675
rect 73065 4635 73123 4641
rect 74721 4675 74779 4681
rect 74721 4641 74733 4675
rect 74767 4672 74779 4675
rect 74994 4672 75000 4684
rect 74767 4644 75000 4672
rect 74767 4641 74779 4644
rect 74721 4635 74779 4641
rect 74994 4632 75000 4644
rect 75052 4632 75058 4684
rect 75362 4632 75368 4684
rect 75420 4672 75426 4684
rect 75549 4675 75607 4681
rect 75549 4672 75561 4675
rect 75420 4644 75561 4672
rect 75420 4632 75426 4644
rect 75549 4641 75561 4644
rect 75595 4641 75607 4675
rect 75549 4635 75607 4641
rect 75914 4632 75920 4684
rect 75972 4672 75978 4684
rect 76650 4672 76656 4684
rect 75972 4644 76656 4672
rect 75972 4632 75978 4644
rect 76650 4632 76656 4644
rect 76708 4632 76714 4684
rect 77496 4672 77524 4712
rect 77570 4700 77576 4752
rect 77628 4740 77634 4752
rect 78033 4743 78091 4749
rect 78033 4740 78045 4743
rect 77628 4712 78045 4740
rect 77628 4700 77634 4712
rect 78033 4709 78045 4712
rect 78079 4709 78091 4743
rect 79226 4740 79232 4752
rect 78033 4703 78091 4709
rect 79060 4712 79232 4740
rect 79060 4672 79088 4712
rect 79226 4700 79232 4712
rect 79284 4700 79290 4752
rect 80238 4740 80244 4752
rect 80199 4712 80244 4740
rect 80238 4700 80244 4712
rect 80296 4700 80302 4752
rect 80882 4700 80888 4752
rect 80940 4740 80946 4752
rect 80977 4743 81035 4749
rect 80977 4740 80989 4743
rect 80940 4712 80989 4740
rect 80940 4700 80946 4712
rect 80977 4709 80989 4712
rect 81023 4709 81035 4743
rect 81989 4743 82047 4749
rect 81989 4740 82001 4743
rect 80977 4703 81035 4709
rect 81084 4712 82001 4740
rect 77496 4644 79088 4672
rect 79137 4675 79195 4681
rect 79137 4641 79149 4675
rect 79183 4672 79195 4675
rect 81084 4672 81112 4712
rect 81989 4709 82001 4712
rect 82035 4709 82047 4743
rect 83642 4740 83648 4752
rect 81989 4703 82047 4709
rect 82464 4712 83648 4740
rect 79183 4644 81112 4672
rect 81805 4675 81863 4681
rect 79183 4641 79195 4644
rect 79137 4635 79195 4641
rect 81805 4641 81817 4675
rect 81851 4672 81863 4675
rect 82464 4672 82492 4712
rect 83642 4700 83648 4712
rect 83700 4700 83706 4752
rect 84841 4743 84899 4749
rect 84841 4709 84853 4743
rect 84887 4740 84899 4743
rect 85117 4743 85175 4749
rect 85117 4740 85129 4743
rect 84887 4712 85129 4740
rect 84887 4709 84899 4712
rect 84841 4703 84899 4709
rect 85117 4709 85129 4712
rect 85163 4740 85175 4743
rect 98086 4740 98092 4752
rect 85163 4712 98092 4740
rect 85163 4709 85175 4712
rect 85117 4703 85175 4709
rect 98086 4700 98092 4712
rect 98144 4700 98150 4752
rect 81851 4644 82492 4672
rect 81851 4641 81863 4644
rect 81805 4635 81863 4641
rect 82814 4632 82820 4684
rect 82872 4672 82878 4684
rect 83093 4675 83151 4681
rect 83093 4672 83105 4675
rect 82872 4644 83105 4672
rect 82872 4632 82878 4644
rect 83093 4641 83105 4644
rect 83139 4641 83151 4675
rect 83093 4635 83151 4641
rect 83185 4675 83243 4681
rect 83185 4641 83197 4675
rect 83231 4672 83243 4675
rect 83461 4675 83519 4681
rect 83231 4644 83265 4672
rect 83231 4641 83243 4644
rect 83185 4635 83243 4641
rect 83461 4641 83473 4675
rect 83507 4672 83519 4675
rect 83918 4672 83924 4684
rect 83507 4644 83924 4672
rect 83507 4641 83519 4644
rect 83461 4635 83519 4641
rect 45278 4564 45284 4616
rect 45336 4604 45342 4616
rect 45738 4604 45744 4616
rect 45336 4576 45744 4604
rect 45336 4564 45342 4576
rect 45738 4564 45744 4576
rect 45796 4604 45802 4616
rect 46014 4604 46020 4616
rect 45796 4576 46020 4604
rect 45796 4564 45802 4576
rect 46014 4564 46020 4576
rect 46072 4604 46078 4616
rect 46201 4607 46259 4613
rect 46201 4604 46213 4607
rect 46072 4576 46213 4604
rect 46072 4564 46078 4576
rect 46201 4573 46213 4576
rect 46247 4573 46259 4607
rect 46201 4567 46259 4573
rect 59630 4564 59636 4616
rect 59688 4604 59694 4616
rect 81621 4607 81679 4613
rect 59688 4576 81480 4604
rect 59688 4564 59694 4576
rect 62114 4536 62120 4548
rect 37240 4508 38056 4536
rect 39132 4508 41414 4536
rect 37240 4496 37246 4508
rect 11977 4471 12035 4477
rect 11977 4437 11989 4471
rect 12023 4468 12035 4471
rect 35894 4468 35900 4480
rect 12023 4440 35900 4468
rect 12023 4437 12035 4440
rect 11977 4431 12035 4437
rect 35894 4428 35900 4440
rect 35952 4428 35958 4480
rect 36630 4428 36636 4480
rect 36688 4468 36694 4480
rect 39132 4468 39160 4508
rect 36688 4440 39160 4468
rect 36688 4428 36694 4440
rect 39206 4428 39212 4480
rect 39264 4468 39270 4480
rect 39758 4468 39764 4480
rect 39264 4440 39764 4468
rect 39264 4428 39270 4440
rect 39758 4428 39764 4440
rect 39816 4428 39822 4480
rect 41386 4468 41414 4508
rect 44744 4508 46244 4536
rect 44744 4468 44772 4508
rect 41386 4440 44772 4468
rect 46216 4468 46244 4508
rect 47136 4508 62120 4536
rect 47136 4468 47164 4508
rect 62114 4496 62120 4508
rect 62172 4496 62178 4548
rect 68002 4496 68008 4548
rect 68060 4536 68066 4548
rect 75365 4539 75423 4545
rect 75365 4536 75377 4539
rect 68060 4508 75377 4536
rect 68060 4496 68066 4508
rect 75365 4505 75377 4508
rect 75411 4505 75423 4539
rect 75365 4499 75423 4505
rect 75454 4496 75460 4548
rect 75512 4536 75518 4548
rect 80698 4536 80704 4548
rect 75512 4508 80704 4536
rect 75512 4496 75518 4508
rect 80698 4496 80704 4508
rect 80756 4496 80762 4548
rect 81161 4539 81219 4545
rect 81161 4505 81173 4539
rect 81207 4536 81219 4539
rect 81342 4536 81348 4548
rect 81207 4508 81348 4536
rect 81207 4505 81219 4508
rect 81161 4499 81219 4505
rect 81342 4496 81348 4508
rect 81400 4496 81406 4548
rect 81452 4536 81480 4576
rect 81621 4573 81633 4607
rect 81667 4604 81679 4607
rect 82538 4604 82544 4616
rect 81667 4576 82544 4604
rect 81667 4573 81679 4576
rect 81621 4567 81679 4573
rect 82538 4564 82544 4576
rect 82596 4564 82602 4616
rect 82998 4564 83004 4616
rect 83056 4604 83062 4616
rect 83200 4604 83228 4635
rect 83918 4632 83924 4644
rect 83976 4632 83982 4684
rect 84010 4632 84016 4684
rect 84068 4672 84074 4684
rect 84105 4675 84163 4681
rect 84105 4672 84117 4675
rect 84068 4644 84117 4672
rect 84068 4632 84074 4644
rect 84105 4641 84117 4644
rect 84151 4641 84163 4675
rect 84105 4635 84163 4641
rect 84197 4675 84255 4681
rect 84197 4641 84209 4675
rect 84243 4641 84255 4675
rect 84197 4635 84255 4641
rect 84473 4675 84531 4681
rect 84473 4641 84485 4675
rect 84519 4672 84531 4675
rect 84519 4644 86448 4672
rect 84519 4641 84531 4644
rect 84473 4635 84531 4641
rect 83369 4607 83427 4613
rect 83369 4604 83381 4607
rect 83056 4576 83381 4604
rect 83056 4564 83062 4576
rect 83369 4573 83381 4576
rect 83415 4604 83427 4607
rect 83642 4604 83648 4616
rect 83415 4576 83648 4604
rect 83415 4573 83427 4576
rect 83369 4567 83427 4573
rect 83642 4564 83648 4576
rect 83700 4604 83706 4616
rect 84212 4604 84240 4635
rect 84381 4607 84439 4613
rect 84381 4604 84393 4607
rect 83700 4576 84393 4604
rect 83700 4564 83706 4576
rect 84381 4573 84393 4576
rect 84427 4573 84439 4607
rect 84381 4567 84439 4573
rect 84933 4539 84991 4545
rect 84933 4536 84945 4539
rect 81452 4508 84945 4536
rect 84933 4505 84945 4508
rect 84979 4505 84991 4539
rect 85482 4536 85488 4548
rect 85443 4508 85488 4536
rect 84933 4499 84991 4505
rect 85482 4496 85488 4508
rect 85540 4496 85546 4548
rect 86420 4536 86448 4644
rect 87506 4632 87512 4684
rect 87564 4672 87570 4684
rect 88153 4675 88211 4681
rect 88153 4672 88165 4675
rect 87564 4644 88165 4672
rect 87564 4632 87570 4644
rect 88153 4641 88165 4644
rect 88199 4641 88211 4675
rect 88153 4635 88211 4641
rect 88334 4632 88340 4684
rect 88392 4672 88398 4684
rect 88797 4675 88855 4681
rect 88797 4672 88809 4675
rect 88392 4644 88809 4672
rect 88392 4632 88398 4644
rect 88797 4641 88809 4644
rect 88843 4641 88855 4675
rect 88797 4635 88855 4641
rect 89346 4632 89352 4684
rect 89404 4672 89410 4684
rect 89441 4675 89499 4681
rect 89441 4672 89453 4675
rect 89404 4644 89453 4672
rect 89404 4632 89410 4644
rect 89441 4641 89453 4644
rect 89487 4641 89499 4675
rect 93762 4672 93768 4684
rect 93723 4644 93768 4672
rect 89441 4635 89499 4641
rect 93762 4632 93768 4644
rect 93820 4632 93826 4684
rect 102594 4672 102600 4684
rect 102555 4644 102600 4672
rect 102594 4632 102600 4644
rect 102652 4632 102658 4684
rect 175366 4672 175372 4684
rect 175327 4644 175372 4672
rect 175366 4632 175372 4644
rect 175424 4632 175430 4684
rect 176197 4675 176255 4681
rect 176197 4641 176209 4675
rect 176243 4641 176255 4675
rect 176197 4635 176255 4641
rect 86494 4564 86500 4616
rect 86552 4604 86558 4616
rect 176212 4604 176240 4635
rect 176654 4632 176660 4684
rect 176712 4672 176718 4684
rect 177301 4675 177359 4681
rect 177301 4672 177313 4675
rect 176712 4644 177313 4672
rect 176712 4632 176718 4644
rect 177301 4641 177313 4644
rect 177347 4641 177359 4675
rect 177942 4672 177948 4684
rect 177903 4644 177948 4672
rect 177301 4635 177359 4641
rect 177942 4632 177948 4644
rect 178000 4632 178006 4684
rect 179782 4604 179788 4616
rect 86552 4576 93992 4604
rect 176212 4576 179788 4604
rect 86552 4564 86558 4576
rect 88150 4536 88156 4548
rect 86420 4508 88156 4536
rect 88150 4496 88156 4508
rect 88208 4496 88214 4548
rect 88337 4539 88395 4545
rect 88337 4505 88349 4539
rect 88383 4536 88395 4539
rect 88426 4536 88432 4548
rect 88383 4508 88432 4536
rect 88383 4505 88395 4508
rect 88337 4499 88395 4505
rect 88426 4496 88432 4508
rect 88484 4496 88490 4548
rect 88978 4536 88984 4548
rect 88939 4508 88984 4536
rect 88978 4496 88984 4508
rect 89036 4496 89042 4548
rect 93964 4545 93992 4576
rect 179782 4564 179788 4576
rect 179840 4564 179846 4616
rect 93949 4539 94007 4545
rect 93949 4505 93961 4539
rect 93995 4505 94007 4539
rect 93949 4499 94007 4505
rect 46216 4440 47164 4468
rect 47581 4471 47639 4477
rect 47581 4437 47593 4471
rect 47627 4468 47639 4471
rect 48314 4468 48320 4480
rect 47627 4440 48320 4468
rect 47627 4437 47639 4440
rect 47581 4431 47639 4437
rect 48314 4428 48320 4440
rect 48372 4468 48378 4480
rect 48590 4468 48596 4480
rect 48372 4440 48596 4468
rect 48372 4428 48378 4440
rect 48590 4428 48596 4440
rect 48648 4428 48654 4480
rect 74718 4428 74724 4480
rect 74776 4468 74782 4480
rect 74905 4471 74963 4477
rect 74905 4468 74917 4471
rect 74776 4440 74917 4468
rect 74776 4428 74782 4440
rect 74905 4437 74917 4440
rect 74951 4468 74963 4471
rect 75638 4468 75644 4480
rect 74951 4440 75644 4468
rect 74951 4437 74963 4440
rect 74905 4431 74963 4437
rect 75638 4428 75644 4440
rect 75696 4428 75702 4480
rect 76742 4468 76748 4480
rect 76703 4440 76748 4468
rect 76742 4428 76748 4440
rect 76800 4428 76806 4480
rect 77938 4428 77944 4480
rect 77996 4468 78002 4480
rect 78125 4471 78183 4477
rect 78125 4468 78137 4471
rect 77996 4440 78137 4468
rect 77996 4428 78002 4440
rect 78125 4437 78137 4440
rect 78171 4437 78183 4471
rect 78125 4431 78183 4437
rect 80146 4428 80152 4480
rect 80204 4468 80210 4480
rect 80333 4471 80391 4477
rect 80333 4468 80345 4471
rect 80204 4440 80345 4468
rect 80204 4428 80210 4440
rect 80333 4437 80345 4440
rect 80379 4437 80391 4471
rect 80333 4431 80391 4437
rect 80882 4428 80888 4480
rect 80940 4468 80946 4480
rect 81710 4468 81716 4480
rect 80940 4440 81716 4468
rect 80940 4428 80946 4440
rect 81710 4428 81716 4440
rect 81768 4428 81774 4480
rect 82262 4428 82268 4480
rect 82320 4468 82326 4480
rect 82909 4471 82967 4477
rect 82909 4468 82921 4471
rect 82320 4440 82921 4468
rect 82320 4428 82326 4440
rect 82909 4437 82921 4440
rect 82955 4437 82967 4471
rect 82909 4431 82967 4437
rect 84654 4428 84660 4480
rect 84712 4468 84718 4480
rect 85117 4471 85175 4477
rect 85117 4468 85129 4471
rect 84712 4440 85129 4468
rect 84712 4428 84718 4440
rect 85117 4437 85129 4440
rect 85163 4437 85175 4471
rect 86126 4468 86132 4480
rect 86087 4440 86132 4468
rect 85117 4431 85175 4437
rect 86126 4428 86132 4440
rect 86184 4428 86190 4480
rect 86773 4471 86831 4477
rect 86773 4437 86785 4471
rect 86819 4468 86831 4471
rect 86954 4468 86960 4480
rect 86819 4440 86960 4468
rect 86819 4437 86831 4440
rect 86773 4431 86831 4437
rect 86954 4428 86960 4440
rect 87012 4428 87018 4480
rect 89162 4428 89168 4480
rect 89220 4468 89226 4480
rect 94498 4468 94504 4480
rect 89220 4440 94504 4468
rect 89220 4428 89226 4440
rect 94498 4428 94504 4440
rect 94556 4428 94562 4480
rect 1104 4378 178848 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 34966 4378
rect 35018 4326 35030 4378
rect 35082 4326 35094 4378
rect 35146 4326 35158 4378
rect 35210 4326 65686 4378
rect 65738 4326 65750 4378
rect 65802 4326 65814 4378
rect 65866 4326 65878 4378
rect 65930 4326 96406 4378
rect 96458 4326 96470 4378
rect 96522 4326 96534 4378
rect 96586 4326 96598 4378
rect 96650 4326 127126 4378
rect 127178 4326 127190 4378
rect 127242 4326 127254 4378
rect 127306 4326 127318 4378
rect 127370 4326 157846 4378
rect 157898 4326 157910 4378
rect 157962 4326 157974 4378
rect 158026 4326 158038 4378
rect 158090 4326 178848 4378
rect 1104 4304 178848 4326
rect 5810 4224 5816 4276
rect 5868 4264 5874 4276
rect 32306 4264 32312 4276
rect 5868 4236 32312 4264
rect 5868 4224 5874 4236
rect 32306 4224 32312 4236
rect 32364 4224 32370 4276
rect 32398 4224 32404 4276
rect 32456 4264 32462 4276
rect 46106 4264 46112 4276
rect 32456 4236 46112 4264
rect 32456 4224 32462 4236
rect 46106 4224 46112 4236
rect 46164 4224 46170 4276
rect 51810 4224 51816 4276
rect 51868 4264 51874 4276
rect 78030 4264 78036 4276
rect 51868 4236 78036 4264
rect 51868 4224 51874 4236
rect 78030 4224 78036 4236
rect 78088 4224 78094 4276
rect 78309 4267 78367 4273
rect 78309 4233 78321 4267
rect 78355 4264 78367 4267
rect 78398 4264 78404 4276
rect 78355 4236 78404 4264
rect 78355 4233 78367 4236
rect 78309 4227 78367 4233
rect 78398 4224 78404 4236
rect 78456 4224 78462 4276
rect 78490 4224 78496 4276
rect 78548 4264 78554 4276
rect 80882 4264 80888 4276
rect 78548 4236 80888 4264
rect 78548 4224 78554 4236
rect 80882 4224 80888 4236
rect 80940 4224 80946 4276
rect 81713 4267 81771 4273
rect 81713 4233 81725 4267
rect 81759 4264 81771 4267
rect 82446 4264 82452 4276
rect 81759 4236 82452 4264
rect 81759 4233 81771 4236
rect 81713 4227 81771 4233
rect 82446 4224 82452 4236
rect 82504 4224 82510 4276
rect 82909 4267 82967 4273
rect 82909 4233 82921 4267
rect 82955 4264 82967 4267
rect 83918 4264 83924 4276
rect 82955 4236 83924 4264
rect 82955 4233 82967 4236
rect 82909 4227 82967 4233
rect 83918 4224 83924 4236
rect 83976 4224 83982 4276
rect 84010 4224 84016 4276
rect 84068 4264 84074 4276
rect 85206 4264 85212 4276
rect 84068 4236 85212 4264
rect 84068 4224 84074 4236
rect 85206 4224 85212 4236
rect 85264 4224 85270 4276
rect 86221 4267 86279 4273
rect 86221 4233 86233 4267
rect 86267 4233 86279 4267
rect 86221 4227 86279 4233
rect 13541 4199 13599 4205
rect 13541 4165 13553 4199
rect 13587 4196 13599 4199
rect 19334 4196 19340 4208
rect 13587 4168 19340 4196
rect 13587 4165 13599 4168
rect 13541 4159 13599 4165
rect 19334 4156 19340 4168
rect 19392 4156 19398 4208
rect 21910 4156 21916 4208
rect 21968 4196 21974 4208
rect 34054 4196 34060 4208
rect 21968 4168 34060 4196
rect 21968 4156 21974 4168
rect 34054 4156 34060 4168
rect 34112 4156 34118 4208
rect 39669 4199 39727 4205
rect 39669 4165 39681 4199
rect 39715 4165 39727 4199
rect 39669 4159 39727 4165
rect 3142 4088 3148 4140
rect 3200 4128 3206 4140
rect 12342 4128 12348 4140
rect 3200 4100 12348 4128
rect 3200 4088 3206 4100
rect 12342 4088 12348 4100
rect 12400 4088 12406 4140
rect 12452 4100 14412 4128
rect 1118 4020 1124 4072
rect 1176 4060 1182 4072
rect 1397 4063 1455 4069
rect 1397 4060 1409 4063
rect 1176 4032 1409 4060
rect 1176 4020 1182 4032
rect 1397 4029 1409 4032
rect 1443 4029 1455 4063
rect 1397 4023 1455 4029
rect 1854 4020 1860 4072
rect 1912 4060 1918 4072
rect 2041 4063 2099 4069
rect 2041 4060 2053 4063
rect 1912 4032 2053 4060
rect 1912 4020 1918 4032
rect 2041 4029 2053 4032
rect 2087 4029 2099 4063
rect 2041 4023 2099 4029
rect 10962 4020 10968 4072
rect 11020 4060 11026 4072
rect 12452 4060 12480 4100
rect 11020 4032 12480 4060
rect 12555 4063 12613 4069
rect 11020 4020 11026 4032
rect 12555 4029 12567 4063
rect 12601 4060 12613 4063
rect 12710 4060 12716 4072
rect 12601 4032 12716 4060
rect 12601 4029 12613 4032
rect 12555 4023 12613 4029
rect 12710 4020 12716 4032
rect 12768 4020 12774 4072
rect 13630 4060 13636 4072
rect 13591 4032 13636 4060
rect 13630 4020 13636 4032
rect 13688 4020 13694 4072
rect 14384 4060 14412 4100
rect 14826 4088 14832 4140
rect 14884 4128 14890 4140
rect 21818 4128 21824 4140
rect 14884 4100 21824 4128
rect 14884 4088 14890 4100
rect 21818 4088 21824 4100
rect 21876 4088 21882 4140
rect 24946 4128 24952 4140
rect 21928 4100 24952 4128
rect 15654 4060 15660 4072
rect 14384 4032 15660 4060
rect 15654 4020 15660 4032
rect 15712 4020 15718 4072
rect 15838 4060 15844 4072
rect 15799 4032 15844 4060
rect 15838 4020 15844 4032
rect 15896 4020 15902 4072
rect 16206 4020 16212 4072
rect 16264 4060 16270 4072
rect 20070 4060 20076 4072
rect 16264 4032 20076 4060
rect 16264 4020 16270 4032
rect 20070 4020 20076 4032
rect 20128 4020 20134 4072
rect 20254 4060 20260 4072
rect 20215 4032 20260 4060
rect 20254 4020 20260 4032
rect 20312 4020 20318 4072
rect 21928 4060 21956 4100
rect 24946 4088 24952 4100
rect 25004 4088 25010 4140
rect 25498 4088 25504 4140
rect 25556 4128 25562 4140
rect 35986 4128 35992 4140
rect 25556 4100 33088 4128
rect 35947 4100 35992 4128
rect 25556 4088 25562 4100
rect 20364 4032 21956 4060
rect 12066 3992 12072 4004
rect 1596 3964 12072 3992
rect 1596 3933 1624 3964
rect 12066 3952 12072 3964
rect 12124 3952 12130 4004
rect 12250 3952 12256 4004
rect 12308 3992 12314 4004
rect 12434 3992 12440 4004
rect 12308 3964 12440 3992
rect 12308 3952 12314 3964
rect 12434 3952 12440 3964
rect 12492 3952 12498 4004
rect 13541 3995 13599 4001
rect 13541 3992 13553 3995
rect 12544 3964 13553 3992
rect 1581 3927 1639 3933
rect 1581 3893 1593 3927
rect 1627 3893 1639 3927
rect 1581 3887 1639 3893
rect 2225 3927 2283 3933
rect 2225 3893 2237 3927
rect 2271 3924 2283 3927
rect 9950 3924 9956 3936
rect 2271 3896 9956 3924
rect 2271 3893 2283 3896
rect 2225 3887 2283 3893
rect 9950 3884 9956 3896
rect 10008 3884 10014 3936
rect 10042 3884 10048 3936
rect 10100 3924 10106 3936
rect 12544 3924 12572 3964
rect 13541 3961 13553 3964
rect 13587 3961 13599 3995
rect 13541 3955 13599 3961
rect 13722 3952 13728 4004
rect 13780 3992 13786 4004
rect 20364 3992 20392 4032
rect 22370 4020 22376 4072
rect 22428 4060 22434 4072
rect 31938 4060 31944 4072
rect 22428 4032 31944 4060
rect 22428 4020 22434 4032
rect 31938 4020 31944 4032
rect 31996 4020 32002 4072
rect 33060 4060 33088 4100
rect 35986 4088 35992 4100
rect 36044 4088 36050 4140
rect 38286 4128 38292 4140
rect 38247 4100 38292 4128
rect 38286 4088 38292 4100
rect 38344 4088 38350 4140
rect 39574 4088 39580 4140
rect 39632 4128 39638 4140
rect 39684 4128 39712 4159
rect 39758 4156 39764 4208
rect 39816 4196 39822 4208
rect 51626 4196 51632 4208
rect 39816 4168 44128 4196
rect 51587 4168 51632 4196
rect 39816 4156 39822 4168
rect 40770 4128 40776 4140
rect 39632 4100 40776 4128
rect 39632 4088 39638 4100
rect 40770 4088 40776 4100
rect 40828 4088 40834 4140
rect 40954 4088 40960 4140
rect 41012 4128 41018 4140
rect 43990 4128 43996 4140
rect 41012 4100 43996 4128
rect 41012 4088 41018 4100
rect 43990 4088 43996 4100
rect 44048 4088 44054 4140
rect 44100 4128 44128 4168
rect 51626 4156 51632 4168
rect 51684 4156 51690 4208
rect 56226 4156 56232 4208
rect 56284 4196 56290 4208
rect 56284 4168 80376 4196
rect 56284 4156 56290 4168
rect 71038 4128 71044 4140
rect 44100 4100 45876 4128
rect 36078 4060 36084 4072
rect 33060 4032 36084 4060
rect 36078 4020 36084 4032
rect 36136 4020 36142 4072
rect 38194 4060 38200 4072
rect 36188 4032 38200 4060
rect 34146 3992 34152 4004
rect 13780 3964 20392 3992
rect 22480 3964 34152 3992
rect 13780 3952 13786 3964
rect 10100 3896 12572 3924
rect 10100 3884 10106 3896
rect 12618 3884 12624 3936
rect 12676 3924 12682 3936
rect 18782 3924 18788 3936
rect 12676 3896 18788 3924
rect 12676 3884 12682 3896
rect 18782 3884 18788 3896
rect 18840 3884 18846 3936
rect 18874 3884 18880 3936
rect 18932 3924 18938 3936
rect 22094 3924 22100 3936
rect 18932 3896 22100 3924
rect 18932 3884 18938 3896
rect 22094 3884 22100 3896
rect 22152 3884 22158 3936
rect 22186 3884 22192 3936
rect 22244 3924 22250 3936
rect 22480 3924 22508 3964
rect 34146 3952 34152 3964
rect 34204 3952 34210 4004
rect 22244 3896 22508 3924
rect 22244 3884 22250 3896
rect 27890 3884 27896 3936
rect 27948 3924 27954 3936
rect 36188 3924 36216 4032
rect 38194 4020 38200 4032
rect 38252 4020 38258 4072
rect 38556 4063 38614 4069
rect 38556 4029 38568 4063
rect 38602 4060 38614 4063
rect 42242 4060 42248 4072
rect 38602 4032 42248 4060
rect 38602 4029 38614 4032
rect 38556 4023 38614 4029
rect 42242 4020 42248 4032
rect 42300 4020 42306 4072
rect 45738 4060 45744 4072
rect 45699 4032 45744 4060
rect 45738 4020 45744 4032
rect 45796 4020 45802 4072
rect 45848 4060 45876 4100
rect 51736 4100 71044 4128
rect 51736 4069 51764 4100
rect 71038 4088 71044 4100
rect 71096 4088 71102 4140
rect 73430 4128 73436 4140
rect 71240 4100 73436 4128
rect 71240 4072 71268 4100
rect 73430 4088 73436 4100
rect 73488 4128 73494 4140
rect 73488 4100 77524 4128
rect 73488 4088 73494 4100
rect 50617 4063 50675 4069
rect 50617 4060 50629 4063
rect 45848 4032 50629 4060
rect 50617 4029 50629 4032
rect 50663 4029 50675 4063
rect 50617 4023 50675 4029
rect 51721 4063 51779 4069
rect 51721 4029 51733 4063
rect 51767 4029 51779 4063
rect 56962 4060 56968 4072
rect 56875 4032 56968 4060
rect 51721 4023 51779 4029
rect 56962 4020 56968 4032
rect 57020 4060 57026 4072
rect 59265 4063 59323 4069
rect 59265 4060 59277 4063
rect 57020 4032 59277 4060
rect 57020 4020 57026 4032
rect 59265 4029 59277 4032
rect 59311 4029 59323 4063
rect 66162 4060 66168 4072
rect 66123 4032 66168 4060
rect 59265 4023 59323 4029
rect 66162 4020 66168 4032
rect 66220 4020 66226 4072
rect 67266 4060 67272 4072
rect 67227 4032 67272 4060
rect 67266 4020 67272 4032
rect 67324 4020 67330 4072
rect 68370 4060 68376 4072
rect 68331 4032 68376 4060
rect 68370 4020 68376 4032
rect 68428 4020 68434 4072
rect 69474 4020 69480 4072
rect 69532 4060 69538 4072
rect 69753 4063 69811 4069
rect 69753 4060 69765 4063
rect 69532 4032 69765 4060
rect 69532 4020 69538 4032
rect 69753 4029 69765 4032
rect 69799 4029 69811 4063
rect 69753 4023 69811 4029
rect 70489 4063 70547 4069
rect 70489 4029 70501 4063
rect 70535 4060 70547 4063
rect 70946 4060 70952 4072
rect 70535 4032 70952 4060
rect 70535 4029 70547 4032
rect 70489 4023 70547 4029
rect 70946 4020 70952 4032
rect 71004 4020 71010 4072
rect 71222 4060 71228 4072
rect 71135 4032 71228 4060
rect 71222 4020 71228 4032
rect 71280 4020 71286 4072
rect 72050 4060 72056 4072
rect 72011 4032 72056 4060
rect 72050 4020 72056 4032
rect 72108 4020 72114 4072
rect 73154 4060 73160 4072
rect 73115 4032 73160 4060
rect 73154 4020 73160 4032
rect 73212 4020 73218 4072
rect 73890 4060 73896 4072
rect 73851 4032 73896 4060
rect 73890 4020 73896 4032
rect 73948 4020 73954 4072
rect 74258 4020 74264 4072
rect 74316 4060 74322 4072
rect 75181 4063 75239 4069
rect 75181 4060 75193 4063
rect 74316 4032 75193 4060
rect 74316 4020 74322 4032
rect 75181 4029 75193 4032
rect 75227 4029 75239 4063
rect 75181 4023 75239 4029
rect 76009 4063 76067 4069
rect 76009 4029 76021 4063
rect 76055 4029 76067 4063
rect 76742 4060 76748 4072
rect 76703 4032 76748 4060
rect 76009 4023 76067 4029
rect 36256 3995 36314 4001
rect 36256 3961 36268 3995
rect 36302 3992 36314 3995
rect 36302 3964 38148 3992
rect 36302 3961 36314 3964
rect 36256 3955 36314 3961
rect 27948 3896 36216 3924
rect 37369 3927 37427 3933
rect 27948 3884 27954 3896
rect 37369 3893 37381 3927
rect 37415 3924 37427 3927
rect 37458 3924 37464 3936
rect 37415 3896 37464 3924
rect 37415 3893 37427 3896
rect 37369 3887 37427 3893
rect 37458 3884 37464 3896
rect 37516 3884 37522 3936
rect 38120 3924 38148 3964
rect 38378 3952 38384 4004
rect 38436 3992 38442 4004
rect 46008 3995 46066 4001
rect 38436 3964 41414 3992
rect 38436 3952 38442 3964
rect 40126 3924 40132 3936
rect 38120 3896 40132 3924
rect 40126 3884 40132 3896
rect 40184 3884 40190 3936
rect 41386 3924 41414 3964
rect 46008 3961 46020 3995
rect 46054 3992 46066 3995
rect 49326 3992 49332 4004
rect 46054 3964 49332 3992
rect 46054 3961 46066 3964
rect 46008 3955 46066 3961
rect 49326 3952 49332 3964
rect 49384 3952 49390 4004
rect 57149 3995 57207 4001
rect 57149 3961 57161 3995
rect 57195 3992 57207 3995
rect 70854 3992 70860 4004
rect 57195 3964 70860 3992
rect 57195 3961 57207 3964
rect 57149 3955 57207 3961
rect 70854 3952 70860 3964
rect 70912 3952 70918 4004
rect 71406 3952 71412 4004
rect 71464 3992 71470 4004
rect 76024 3992 76052 4023
rect 76742 4020 76748 4032
rect 76800 4020 76806 4072
rect 77496 4069 77524 4100
rect 77570 4088 77576 4140
rect 77628 4128 77634 4140
rect 77665 4131 77723 4137
rect 77665 4128 77677 4131
rect 77628 4100 77677 4128
rect 77628 4088 77634 4100
rect 77665 4097 77677 4100
rect 77711 4128 77723 4131
rect 78490 4128 78496 4140
rect 77711 4100 78496 4128
rect 77711 4097 77723 4100
rect 77665 4091 77723 4097
rect 78490 4088 78496 4100
rect 78548 4088 78554 4140
rect 79137 4131 79195 4137
rect 79137 4097 79149 4131
rect 79183 4128 79195 4131
rect 80238 4128 80244 4140
rect 79183 4100 80244 4128
rect 79183 4097 79195 4100
rect 79137 4091 79195 4097
rect 80238 4088 80244 4100
rect 80296 4088 80302 4140
rect 80348 4128 80376 4168
rect 80422 4156 80428 4208
rect 80480 4196 80486 4208
rect 82354 4196 82360 4208
rect 80480 4168 82360 4196
rect 80480 4156 80486 4168
rect 82354 4156 82360 4168
rect 82412 4156 82418 4208
rect 84102 4196 84108 4208
rect 82924 4168 84108 4196
rect 81894 4128 81900 4140
rect 80348 4100 81900 4128
rect 81894 4088 81900 4100
rect 81952 4088 81958 4140
rect 77481 4063 77539 4069
rect 77481 4029 77493 4063
rect 77527 4060 77539 4063
rect 78122 4060 78128 4072
rect 77527 4032 78128 4060
rect 77527 4029 77539 4032
rect 77481 4023 77539 4029
rect 78122 4020 78128 4032
rect 78180 4020 78186 4072
rect 79962 4020 79968 4072
rect 80020 4060 80026 4072
rect 80333 4063 80391 4069
rect 80333 4060 80345 4063
rect 80020 4032 80345 4060
rect 80020 4020 80026 4032
rect 80333 4029 80345 4032
rect 80379 4029 80391 4063
rect 80333 4023 80391 4029
rect 80422 4020 80428 4072
rect 80480 4060 80486 4072
rect 80698 4060 80704 4072
rect 80480 4032 80704 4060
rect 80480 4020 80486 4032
rect 80698 4020 80704 4032
rect 80756 4020 80762 4072
rect 81345 4063 81403 4069
rect 81345 4060 81357 4063
rect 80808 4032 81357 4060
rect 78214 3992 78220 4004
rect 71464 3964 75040 3992
rect 76024 3964 76972 3992
rect 78175 3964 78220 3992
rect 71464 3952 71470 3964
rect 47121 3927 47179 3933
rect 47121 3924 47133 3927
rect 41386 3896 47133 3924
rect 47121 3893 47133 3896
rect 47167 3924 47179 3927
rect 48222 3924 48228 3936
rect 47167 3896 48228 3924
rect 47167 3893 47179 3896
rect 47121 3887 47179 3893
rect 48222 3884 48228 3896
rect 48280 3884 48286 3936
rect 59357 3927 59415 3933
rect 59357 3893 59369 3927
rect 59403 3924 59415 3927
rect 70394 3924 70400 3936
rect 59403 3896 70400 3924
rect 59403 3893 59415 3896
rect 59357 3887 59415 3893
rect 70394 3884 70400 3896
rect 70452 3884 70458 3936
rect 71038 3884 71044 3936
rect 71096 3924 71102 3936
rect 71498 3924 71504 3936
rect 71096 3896 71504 3924
rect 71096 3884 71102 3896
rect 71498 3884 71504 3896
rect 71556 3884 71562 3936
rect 75012 3933 75040 3964
rect 74997 3927 75055 3933
rect 74997 3893 75009 3927
rect 75043 3893 75055 3927
rect 74997 3887 75055 3893
rect 75086 3884 75092 3936
rect 75144 3924 75150 3936
rect 76193 3927 76251 3933
rect 76193 3924 76205 3927
rect 75144 3896 76205 3924
rect 75144 3884 75150 3896
rect 76193 3893 76205 3896
rect 76239 3893 76251 3927
rect 76834 3924 76840 3936
rect 76795 3896 76840 3924
rect 76193 3887 76251 3893
rect 76834 3884 76840 3896
rect 76892 3884 76898 3936
rect 76944 3924 76972 3964
rect 78214 3952 78220 3964
rect 78272 3992 78278 4004
rect 78953 3995 79011 4001
rect 78953 3992 78965 3995
rect 78272 3964 78965 3992
rect 78272 3952 78278 3964
rect 78953 3961 78965 3964
rect 78999 3961 79011 3995
rect 78953 3955 79011 3961
rect 79134 3952 79140 4004
rect 79192 3992 79198 4004
rect 80517 3995 80575 4001
rect 80517 3992 80529 3995
rect 79192 3964 80529 3992
rect 79192 3952 79198 3964
rect 80517 3961 80529 3964
rect 80563 3961 80575 3995
rect 80517 3955 80575 3961
rect 77570 3924 77576 3936
rect 76944 3896 77576 3924
rect 77570 3884 77576 3896
rect 77628 3884 77634 3936
rect 79594 3884 79600 3936
rect 79652 3924 79658 3936
rect 80054 3924 80060 3936
rect 79652 3896 80060 3924
rect 79652 3884 79658 3896
rect 80054 3884 80060 3896
rect 80112 3884 80118 3936
rect 80330 3884 80336 3936
rect 80388 3924 80394 3936
rect 80808 3924 80836 4032
rect 81345 4029 81357 4032
rect 81391 4029 81403 4063
rect 82924 4060 82952 4168
rect 84102 4156 84108 4168
rect 84160 4156 84166 4208
rect 84562 4196 84568 4208
rect 84523 4168 84568 4196
rect 84562 4156 84568 4168
rect 84620 4156 84626 4208
rect 85022 4156 85028 4208
rect 85080 4196 85086 4208
rect 86236 4196 86264 4227
rect 86862 4224 86868 4276
rect 86920 4264 86926 4276
rect 86920 4236 87736 4264
rect 86920 4224 86926 4236
rect 87046 4196 87052 4208
rect 85080 4168 87052 4196
rect 85080 4156 85086 4168
rect 87046 4156 87052 4168
rect 87104 4156 87110 4208
rect 82998 4088 83004 4140
rect 83056 4128 83062 4140
rect 83369 4131 83427 4137
rect 83369 4128 83381 4131
rect 83056 4100 83381 4128
rect 83056 4088 83062 4100
rect 83200 4069 83228 4100
rect 83369 4097 83381 4100
rect 83415 4097 83427 4131
rect 87598 4128 87604 4140
rect 83369 4091 83427 4097
rect 83844 4100 87604 4128
rect 83093 4063 83151 4069
rect 83093 4060 83105 4063
rect 81345 4023 81403 4029
rect 81728 4032 83105 4060
rect 80882 3952 80888 4004
rect 80940 3992 80946 4004
rect 81728 3992 81756 4032
rect 83093 4029 83105 4032
rect 83139 4029 83151 4063
rect 83093 4023 83151 4029
rect 83185 4063 83243 4069
rect 83185 4029 83197 4063
rect 83231 4060 83243 4063
rect 83461 4063 83519 4069
rect 83231 4032 83265 4060
rect 83231 4029 83243 4032
rect 83185 4023 83243 4029
rect 83461 4029 83473 4063
rect 83507 4060 83519 4063
rect 83734 4060 83740 4072
rect 83507 4032 83740 4060
rect 83507 4029 83519 4032
rect 83461 4023 83519 4029
rect 83734 4020 83740 4032
rect 83792 4020 83798 4072
rect 80940 3964 81756 3992
rect 80940 3952 80946 3964
rect 81802 3952 81808 4004
rect 81860 3992 81866 4004
rect 82814 3992 82820 4004
rect 81860 3964 82820 3992
rect 81860 3952 81866 3964
rect 82814 3952 82820 3964
rect 82872 3992 82878 4004
rect 83844 3992 83872 4100
rect 87598 4088 87604 4100
rect 87656 4088 87662 4140
rect 87708 4128 87736 4236
rect 88518 4224 88524 4276
rect 88576 4264 88582 4276
rect 88613 4267 88671 4273
rect 88613 4264 88625 4267
rect 88576 4236 88625 4264
rect 88576 4224 88582 4236
rect 88613 4233 88625 4236
rect 88659 4233 88671 4267
rect 88613 4227 88671 4233
rect 88702 4224 88708 4276
rect 88760 4264 88766 4276
rect 88797 4267 88855 4273
rect 88797 4264 88809 4267
rect 88760 4236 88809 4264
rect 88760 4224 88766 4236
rect 88797 4233 88809 4236
rect 88843 4233 88855 4267
rect 89438 4264 89444 4276
rect 89399 4236 89444 4264
rect 88797 4227 88855 4233
rect 89438 4224 89444 4236
rect 89496 4224 89502 4276
rect 89530 4224 89536 4276
rect 89588 4264 89594 4276
rect 109310 4264 109316 4276
rect 89588 4236 109316 4264
rect 89588 4224 89594 4236
rect 109310 4224 109316 4236
rect 109368 4224 109374 4276
rect 87785 4199 87843 4205
rect 87785 4165 87797 4199
rect 87831 4196 87843 4199
rect 90818 4196 90824 4208
rect 87831 4168 90824 4196
rect 87831 4165 87843 4168
rect 87785 4159 87843 4165
rect 90818 4156 90824 4168
rect 90876 4156 90882 4208
rect 90913 4199 90971 4205
rect 90913 4165 90925 4199
rect 90959 4165 90971 4199
rect 90913 4159 90971 4165
rect 87708 4100 89208 4128
rect 84194 4060 84200 4072
rect 84155 4032 84200 4060
rect 84194 4020 84200 4032
rect 84252 4020 84258 4072
rect 84381 4063 84439 4069
rect 84381 4029 84393 4063
rect 84427 4060 84439 4063
rect 85853 4063 85911 4069
rect 84427 4032 84516 4060
rect 84427 4029 84439 4032
rect 84381 4023 84439 4029
rect 82872 3964 83872 3992
rect 82872 3952 82878 3964
rect 83918 3952 83924 4004
rect 83976 3992 83982 4004
rect 84013 3995 84071 4001
rect 84013 3992 84025 3995
rect 83976 3964 84025 3992
rect 83976 3952 83982 3964
rect 84013 3961 84025 3964
rect 84059 3961 84071 3995
rect 84488 3992 84516 4032
rect 85853 4029 85865 4063
rect 85899 4060 85911 4063
rect 86678 4060 86684 4072
rect 85899 4032 86684 4060
rect 85899 4029 85911 4032
rect 85853 4023 85911 4029
rect 84562 3992 84568 4004
rect 84488 3964 84568 3992
rect 84013 3955 84071 3961
rect 84562 3952 84568 3964
rect 84620 3952 84626 4004
rect 85390 3952 85396 4004
rect 85448 3992 85454 4004
rect 85868 3992 85896 4023
rect 86678 4020 86684 4032
rect 86736 4020 86742 4072
rect 86954 4060 86960 4072
rect 86915 4032 86960 4060
rect 86954 4020 86960 4032
rect 87012 4020 87018 4072
rect 87782 4020 87788 4072
rect 87840 4060 87846 4072
rect 88245 4063 88303 4069
rect 88245 4060 88257 4063
rect 87840 4032 88257 4060
rect 87840 4020 87846 4032
rect 88245 4029 88257 4032
rect 88291 4029 88303 4063
rect 88245 4023 88303 4029
rect 88444 4032 89116 4060
rect 85448 3964 85896 3992
rect 85960 3964 87184 3992
rect 85448 3952 85454 3964
rect 81710 3924 81716 3936
rect 80388 3896 80836 3924
rect 81671 3896 81716 3924
rect 80388 3884 80394 3896
rect 81710 3884 81716 3896
rect 81768 3884 81774 3936
rect 81894 3924 81900 3936
rect 81855 3896 81900 3924
rect 81894 3884 81900 3896
rect 81952 3884 81958 3936
rect 84289 3927 84347 3933
rect 84289 3893 84301 3927
rect 84335 3924 84347 3927
rect 85022 3924 85028 3936
rect 84335 3896 85028 3924
rect 84335 3893 84347 3896
rect 84289 3887 84347 3893
rect 85022 3884 85028 3896
rect 85080 3884 85086 3936
rect 85666 3884 85672 3936
rect 85724 3924 85730 3936
rect 85960 3924 85988 3964
rect 86218 3924 86224 3936
rect 85724 3896 85988 3924
rect 86179 3896 86224 3924
rect 85724 3884 85730 3896
rect 86218 3884 86224 3896
rect 86276 3884 86282 3936
rect 86405 3927 86463 3933
rect 86405 3893 86417 3927
rect 86451 3924 86463 3927
rect 86586 3924 86592 3936
rect 86451 3896 86592 3924
rect 86451 3893 86463 3896
rect 86405 3887 86463 3893
rect 86586 3884 86592 3896
rect 86644 3884 86650 3936
rect 86770 3884 86776 3936
rect 86828 3924 86834 3936
rect 87049 3927 87107 3933
rect 87049 3924 87061 3927
rect 86828 3896 87061 3924
rect 86828 3884 86834 3896
rect 87049 3893 87061 3896
rect 87095 3893 87107 3927
rect 87156 3924 87184 3964
rect 88444 3924 88472 4032
rect 88610 3992 88616 4004
rect 88571 3964 88616 3992
rect 88610 3952 88616 3964
rect 88668 3952 88674 4004
rect 87156 3896 88472 3924
rect 89088 3924 89116 4032
rect 89180 3992 89208 4100
rect 89714 4088 89720 4140
rect 89772 4128 89778 4140
rect 90928 4128 90956 4159
rect 91094 4156 91100 4208
rect 91152 4196 91158 4208
rect 92382 4196 92388 4208
rect 91152 4168 92388 4196
rect 91152 4156 91158 4168
rect 92382 4156 92388 4168
rect 92440 4156 92446 4208
rect 94317 4199 94375 4205
rect 94317 4165 94329 4199
rect 94363 4165 94375 4199
rect 94317 4159 94375 4165
rect 89772 4100 90956 4128
rect 89772 4088 89778 4100
rect 91002 4088 91008 4140
rect 91060 4128 91066 4140
rect 94332 4128 94360 4159
rect 94498 4156 94504 4208
rect 94556 4196 94562 4208
rect 109954 4196 109960 4208
rect 94556 4168 109960 4196
rect 94556 4156 94562 4168
rect 109954 4156 109960 4168
rect 110012 4156 110018 4208
rect 91060 4100 94360 4128
rect 91060 4088 91066 4100
rect 94406 4088 94412 4140
rect 94464 4128 94470 4140
rect 94464 4100 96292 4128
rect 94464 4088 94470 4100
rect 90450 4020 90456 4072
rect 90508 4060 90514 4072
rect 90729 4063 90787 4069
rect 90729 4060 90741 4063
rect 90508 4032 90741 4060
rect 90508 4020 90514 4032
rect 90729 4029 90741 4032
rect 90775 4029 90787 4063
rect 91554 4060 91560 4072
rect 91515 4032 91560 4060
rect 90729 4023 90787 4029
rect 91554 4020 91560 4032
rect 91612 4020 91618 4072
rect 91646 4020 91652 4072
rect 91704 4060 91710 4072
rect 92385 4063 92443 4069
rect 91704 4032 91876 4060
rect 91704 4020 91710 4032
rect 91848 3992 91876 4032
rect 92385 4029 92397 4063
rect 92431 4060 92443 4063
rect 92658 4060 92664 4072
rect 92431 4032 92664 4060
rect 92431 4029 92443 4032
rect 92385 4023 92443 4029
rect 92658 4020 92664 4032
rect 92716 4020 92722 4072
rect 93026 4060 93032 4072
rect 92987 4032 93032 4060
rect 93026 4020 93032 4032
rect 93084 4020 93090 4072
rect 94130 4060 94136 4072
rect 94091 4032 94136 4060
rect 94130 4020 94136 4032
rect 94188 4020 94194 4072
rect 94866 4060 94872 4072
rect 94827 4032 94872 4060
rect 94866 4020 94872 4032
rect 94924 4020 94930 4072
rect 95970 4060 95976 4072
rect 95931 4032 95976 4060
rect 95970 4020 95976 4032
rect 96028 4020 96034 4072
rect 96264 3992 96292 4100
rect 97994 4088 98000 4140
rect 98052 4128 98058 4140
rect 102870 4128 102876 4140
rect 98052 4100 102876 4128
rect 98052 4088 98058 4100
rect 102870 4088 102876 4100
rect 102928 4088 102934 4140
rect 104713 4131 104771 4137
rect 104713 4128 104725 4131
rect 103072 4100 104725 4128
rect 97074 4060 97080 4072
rect 97035 4032 97080 4060
rect 97074 4020 97080 4032
rect 97132 4020 97138 4072
rect 98178 4060 98184 4072
rect 98139 4032 98184 4060
rect 98178 4020 98184 4032
rect 98236 4020 98242 4072
rect 99282 4060 99288 4072
rect 99243 4032 99288 4060
rect 99282 4020 99288 4032
rect 99340 4020 99346 4072
rect 100386 4020 100392 4072
rect 100444 4060 100450 4072
rect 101217 4063 101275 4069
rect 101217 4060 101229 4063
rect 100444 4032 101229 4060
rect 100444 4020 100450 4032
rect 101217 4029 101229 4032
rect 101263 4029 101275 4063
rect 101217 4023 101275 4029
rect 101490 4020 101496 4072
rect 101548 4060 101554 4072
rect 101861 4063 101919 4069
rect 101861 4060 101873 4063
rect 101548 4032 101873 4060
rect 101548 4020 101554 4032
rect 101861 4029 101873 4032
rect 101907 4029 101919 4063
rect 102962 4060 102968 4072
rect 102923 4032 102968 4060
rect 101861 4023 101919 4029
rect 102962 4020 102968 4032
rect 103020 4020 103026 4072
rect 89180 3964 91784 3992
rect 91848 3964 96200 3992
rect 96264 3964 99374 3992
rect 91646 3924 91652 3936
rect 89088 3896 91652 3924
rect 87049 3887 87107 3893
rect 91646 3884 91652 3896
rect 91704 3884 91710 3936
rect 91756 3933 91784 3964
rect 91741 3927 91799 3933
rect 91741 3893 91753 3927
rect 91787 3893 91799 3927
rect 91741 3887 91799 3893
rect 91830 3884 91836 3936
rect 91888 3924 91894 3936
rect 92569 3927 92627 3933
rect 92569 3924 92581 3927
rect 91888 3896 92581 3924
rect 91888 3884 91894 3896
rect 92569 3893 92581 3896
rect 92615 3893 92627 3927
rect 93210 3924 93216 3936
rect 93171 3896 93216 3924
rect 92569 3887 92627 3893
rect 93210 3884 93216 3896
rect 93268 3884 93274 3936
rect 95050 3924 95056 3936
rect 95011 3896 95056 3924
rect 95050 3884 95056 3896
rect 95108 3884 95114 3936
rect 96172 3933 96200 3964
rect 96157 3927 96215 3933
rect 96157 3893 96169 3927
rect 96203 3893 96215 3927
rect 97258 3924 97264 3936
rect 97219 3896 97264 3924
rect 96157 3887 96215 3893
rect 97258 3884 97264 3896
rect 97316 3884 97322 3936
rect 98362 3924 98368 3936
rect 98323 3896 98368 3924
rect 98362 3884 98368 3896
rect 98420 3884 98426 3936
rect 99346 3924 99374 3964
rect 101030 3952 101036 4004
rect 101088 3992 101094 4004
rect 103072 3992 103100 4100
rect 104713 4097 104725 4100
rect 104759 4097 104771 4131
rect 104713 4091 104771 4097
rect 103701 4063 103759 4069
rect 103701 4029 103713 4063
rect 103747 4060 103759 4063
rect 103790 4060 103796 4072
rect 103747 4032 103796 4060
rect 103747 4029 103759 4032
rect 103701 4023 103759 4029
rect 103790 4020 103796 4032
rect 103848 4020 103854 4072
rect 104802 4060 104808 4072
rect 104763 4032 104808 4060
rect 104802 4020 104808 4032
rect 104860 4020 104866 4072
rect 105906 4020 105912 4072
rect 105964 4060 105970 4072
rect 106461 4063 106519 4069
rect 106461 4060 106473 4063
rect 105964 4032 106473 4060
rect 105964 4020 105970 4032
rect 106461 4029 106473 4032
rect 106507 4029 106519 4063
rect 106461 4023 106519 4029
rect 107010 4020 107016 4072
rect 107068 4060 107074 4072
rect 107105 4063 107163 4069
rect 107105 4060 107117 4063
rect 107068 4032 107117 4060
rect 107068 4020 107074 4032
rect 107105 4029 107117 4032
rect 107151 4029 107163 4063
rect 107105 4023 107163 4029
rect 111426 4020 111432 4072
rect 111484 4060 111490 4072
rect 111705 4063 111763 4069
rect 111705 4060 111717 4063
rect 111484 4032 111717 4060
rect 111484 4020 111490 4032
rect 111705 4029 111717 4032
rect 111751 4029 111763 4063
rect 112530 4060 112536 4072
rect 112491 4032 112536 4060
rect 111705 4023 111763 4029
rect 112530 4020 112536 4032
rect 112588 4020 112594 4072
rect 113634 4060 113640 4072
rect 113595 4032 113640 4060
rect 113634 4020 113640 4032
rect 113692 4020 113698 4072
rect 114738 4060 114744 4072
rect 114699 4032 114744 4060
rect 114738 4020 114744 4032
rect 114796 4020 114802 4072
rect 115842 4060 115848 4072
rect 115803 4032 115848 4060
rect 115842 4020 115848 4032
rect 115900 4020 115906 4072
rect 116946 4060 116952 4072
rect 116907 4032 116952 4060
rect 116946 4020 116952 4032
rect 117004 4020 117010 4072
rect 118050 4060 118056 4072
rect 118011 4032 118056 4060
rect 118050 4020 118056 4032
rect 118108 4020 118114 4072
rect 119154 4060 119160 4072
rect 119115 4032 119160 4060
rect 119154 4020 119160 4032
rect 119212 4020 119218 4072
rect 120166 4060 120172 4072
rect 120127 4032 120172 4060
rect 120166 4020 120172 4032
rect 120224 4020 120230 4072
rect 121089 4063 121147 4069
rect 121089 4029 121101 4063
rect 121135 4060 121147 4063
rect 121270 4060 121276 4072
rect 121135 4032 121276 4060
rect 121135 4029 121147 4032
rect 121089 4023 121147 4029
rect 121270 4020 121276 4032
rect 121328 4020 121334 4072
rect 122282 4020 122288 4072
rect 122340 4060 122346 4072
rect 122377 4063 122435 4069
rect 122377 4060 122389 4063
rect 122340 4032 122389 4060
rect 122340 4020 122346 4032
rect 122377 4029 122389 4032
rect 122423 4029 122435 4063
rect 123478 4060 123484 4072
rect 123439 4032 123484 4060
rect 122377 4023 122435 4029
rect 123478 4020 123484 4032
rect 123536 4020 123542 4072
rect 124582 4060 124588 4072
rect 124543 4032 124588 4060
rect 124582 4020 124588 4032
rect 124640 4020 124646 4072
rect 125686 4060 125692 4072
rect 125647 4032 125692 4060
rect 125686 4020 125692 4032
rect 125744 4020 125750 4072
rect 126790 4020 126796 4072
rect 126848 4060 126854 4072
rect 127437 4063 127495 4069
rect 127437 4060 127449 4063
rect 126848 4032 127449 4060
rect 126848 4020 126854 4032
rect 127437 4029 127449 4032
rect 127483 4029 127495 4063
rect 127437 4023 127495 4029
rect 127894 4020 127900 4072
rect 127952 4060 127958 4072
rect 128081 4063 128139 4069
rect 128081 4060 128093 4063
rect 127952 4032 128093 4060
rect 127952 4020 127958 4032
rect 128081 4029 128093 4032
rect 128127 4029 128139 4063
rect 131206 4060 131212 4072
rect 131167 4032 131212 4060
rect 128081 4023 128139 4029
rect 131206 4020 131212 4032
rect 131264 4020 131270 4072
rect 133414 4060 133420 4072
rect 133375 4032 133420 4060
rect 133414 4020 133420 4032
rect 133472 4020 133478 4072
rect 134518 4060 134524 4072
rect 134479 4032 134524 4060
rect 134518 4020 134524 4032
rect 134576 4020 134582 4072
rect 136726 4060 136732 4072
rect 136687 4032 136732 4060
rect 136726 4020 136732 4032
rect 136784 4020 136790 4072
rect 137830 4020 137836 4072
rect 137888 4060 137894 4072
rect 137925 4063 137983 4069
rect 137925 4060 137937 4063
rect 137888 4032 137937 4060
rect 137888 4020 137894 4032
rect 137925 4029 137937 4032
rect 137971 4029 137983 4063
rect 138934 4060 138940 4072
rect 138895 4032 138940 4060
rect 137925 4023 137983 4029
rect 138934 4020 138940 4032
rect 138992 4020 138998 4072
rect 140038 4060 140044 4072
rect 139999 4032 140044 4060
rect 140038 4020 140044 4032
rect 140096 4020 140102 4072
rect 141142 4060 141148 4072
rect 141103 4032 141148 4060
rect 141142 4020 141148 4032
rect 141200 4020 141206 4072
rect 142065 4063 142123 4069
rect 142065 4029 142077 4063
rect 142111 4060 142123 4063
rect 142246 4060 142252 4072
rect 142111 4032 142252 4060
rect 142111 4029 142123 4032
rect 142065 4023 142123 4029
rect 142246 4020 142252 4032
rect 142304 4020 142310 4072
rect 143353 4063 143411 4069
rect 143353 4029 143365 4063
rect 143399 4060 143411 4063
rect 143442 4060 143448 4072
rect 143399 4032 143448 4060
rect 143399 4029 143411 4032
rect 143353 4023 143411 4029
rect 143442 4020 143448 4032
rect 143500 4020 143506 4072
rect 144454 4060 144460 4072
rect 144415 4032 144460 4060
rect 144454 4020 144460 4032
rect 144512 4020 144518 4072
rect 145558 4060 145564 4072
rect 145519 4032 145564 4060
rect 145558 4020 145564 4032
rect 145616 4020 145622 4072
rect 146662 4060 146668 4072
rect 146623 4032 146668 4060
rect 146662 4020 146668 4032
rect 146720 4020 146726 4072
rect 147766 4020 147772 4072
rect 147824 4060 147830 4072
rect 148413 4063 148471 4069
rect 148413 4060 148425 4063
rect 147824 4032 148425 4060
rect 147824 4020 147830 4032
rect 148413 4029 148425 4032
rect 148459 4029 148471 4063
rect 148413 4023 148471 4029
rect 148870 4020 148876 4072
rect 148928 4060 148934 4072
rect 149057 4063 149115 4069
rect 149057 4060 149069 4063
rect 148928 4032 149069 4060
rect 148928 4020 148934 4032
rect 149057 4029 149069 4032
rect 149103 4029 149115 4063
rect 152182 4060 152188 4072
rect 152143 4032 152188 4060
rect 149057 4023 149115 4029
rect 152182 4020 152188 4032
rect 152240 4020 152246 4072
rect 153286 4020 153292 4072
rect 153344 4060 153350 4072
rect 153657 4063 153715 4069
rect 153657 4060 153669 4063
rect 153344 4032 153669 4060
rect 153344 4020 153350 4032
rect 153657 4029 153669 4032
rect 153703 4029 153715 4063
rect 154390 4060 154396 4072
rect 154351 4032 154396 4060
rect 153657 4023 153715 4029
rect 154390 4020 154396 4032
rect 154448 4020 154454 4072
rect 155494 4060 155500 4072
rect 155455 4032 155500 4060
rect 155494 4020 155500 4032
rect 155552 4020 155558 4072
rect 157702 4060 157708 4072
rect 157663 4032 157708 4060
rect 157702 4020 157708 4032
rect 157760 4020 157766 4072
rect 158806 4020 158812 4072
rect 158864 4060 158870 4072
rect 158901 4063 158959 4069
rect 158901 4060 158913 4063
rect 158864 4032 158913 4060
rect 158864 4020 158870 4032
rect 158901 4029 158913 4032
rect 158947 4029 158959 4063
rect 159910 4060 159916 4072
rect 159871 4032 159916 4060
rect 158901 4023 158959 4029
rect 159910 4020 159916 4032
rect 159968 4020 159974 4072
rect 161014 4060 161020 4072
rect 160975 4032 161020 4060
rect 161014 4020 161020 4032
rect 161072 4020 161078 4072
rect 162118 4060 162124 4072
rect 162079 4032 162124 4060
rect 162118 4020 162124 4032
rect 162176 4020 162182 4072
rect 165430 4060 165436 4072
rect 165391 4032 165436 4060
rect 165430 4020 165436 4032
rect 165488 4020 165494 4072
rect 166534 4060 166540 4072
rect 166495 4032 166540 4060
rect 166534 4020 166540 4032
rect 166592 4020 166598 4072
rect 167638 4060 167644 4072
rect 167599 4032 167644 4060
rect 167638 4020 167644 4032
rect 167696 4020 167702 4072
rect 168742 4020 168748 4072
rect 168800 4060 168806 4072
rect 169389 4063 169447 4069
rect 169389 4060 169401 4063
rect 168800 4032 169401 4060
rect 168800 4020 168806 4032
rect 169389 4029 169401 4032
rect 169435 4029 169447 4063
rect 169389 4023 169447 4029
rect 169846 4020 169852 4072
rect 169904 4060 169910 4072
rect 170033 4063 170091 4069
rect 170033 4060 170045 4063
rect 169904 4032 170045 4060
rect 169904 4020 169910 4032
rect 170033 4029 170045 4032
rect 170079 4029 170091 4063
rect 170033 4023 170091 4029
rect 173066 4020 173072 4072
rect 173124 4060 173130 4072
rect 173161 4063 173219 4069
rect 173161 4060 173173 4063
rect 173124 4032 173173 4060
rect 173124 4020 173130 4032
rect 173161 4029 173173 4032
rect 173207 4029 173219 4063
rect 173161 4023 173219 4029
rect 174262 4020 174268 4072
rect 174320 4060 174326 4072
rect 174633 4063 174691 4069
rect 174633 4060 174645 4063
rect 174320 4032 174645 4060
rect 174320 4020 174326 4032
rect 174633 4029 174645 4032
rect 174679 4029 174691 4063
rect 175734 4060 175740 4072
rect 175695 4032 175740 4060
rect 174633 4023 174691 4029
rect 175734 4020 175740 4032
rect 175792 4020 175798 4072
rect 176933 4063 176991 4069
rect 176933 4029 176945 4063
rect 176979 4060 176991 4063
rect 177298 4060 177304 4072
rect 176979 4032 177304 4060
rect 176979 4029 176991 4032
rect 176933 4023 176991 4029
rect 177298 4020 177304 4032
rect 177356 4020 177362 4072
rect 177393 4063 177451 4069
rect 177393 4029 177405 4063
rect 177439 4029 177451 4063
rect 177393 4023 177451 4029
rect 101088 3964 103100 3992
rect 101088 3952 101094 3964
rect 103514 3952 103520 4004
rect 103572 3992 103578 4004
rect 103572 3964 106688 3992
rect 103572 3952 103578 3964
rect 99469 3927 99527 3933
rect 99469 3924 99481 3927
rect 99346 3896 99481 3924
rect 99469 3893 99481 3896
rect 99515 3893 99527 3927
rect 101398 3924 101404 3936
rect 101359 3896 101404 3924
rect 99469 3887 99527 3893
rect 101398 3884 101404 3896
rect 101456 3884 101462 3936
rect 102042 3924 102048 3936
rect 102003 3896 102048 3924
rect 102042 3884 102048 3896
rect 102100 3884 102106 3936
rect 103054 3884 103060 3936
rect 103112 3924 103118 3936
rect 103149 3927 103207 3933
rect 103149 3924 103161 3927
rect 103112 3896 103161 3924
rect 103112 3884 103118 3896
rect 103149 3893 103161 3896
rect 103195 3893 103207 3927
rect 103882 3924 103888 3936
rect 103843 3896 103888 3924
rect 103149 3887 103207 3893
rect 103882 3884 103888 3896
rect 103940 3884 103946 3936
rect 106660 3933 106688 3964
rect 176838 3952 176844 4004
rect 176896 3992 176902 4004
rect 177408 3992 177436 4023
rect 176896 3964 177436 3992
rect 176896 3952 176902 3964
rect 104713 3927 104771 3933
rect 104713 3893 104725 3927
rect 104759 3924 104771 3927
rect 104989 3927 105047 3933
rect 104989 3924 105001 3927
rect 104759 3896 105001 3924
rect 104759 3893 104771 3896
rect 104713 3887 104771 3893
rect 104989 3893 105001 3896
rect 105035 3893 105047 3927
rect 104989 3887 105047 3893
rect 106645 3927 106703 3933
rect 106645 3893 106657 3927
rect 106691 3893 106703 3927
rect 107286 3924 107292 3936
rect 107247 3896 107292 3924
rect 106645 3887 106703 3893
rect 107286 3884 107292 3896
rect 107344 3884 107350 3936
rect 107470 3884 107476 3936
rect 107528 3924 107534 3936
rect 111889 3927 111947 3933
rect 111889 3924 111901 3927
rect 107528 3896 111901 3924
rect 107528 3884 107534 3896
rect 111889 3893 111901 3896
rect 111935 3893 111947 3927
rect 111889 3887 111947 3893
rect 1104 3834 178848 3856
rect 1104 3782 19606 3834
rect 19658 3782 19670 3834
rect 19722 3782 19734 3834
rect 19786 3782 19798 3834
rect 19850 3782 50326 3834
rect 50378 3782 50390 3834
rect 50442 3782 50454 3834
rect 50506 3782 50518 3834
rect 50570 3782 81046 3834
rect 81098 3782 81110 3834
rect 81162 3782 81174 3834
rect 81226 3782 81238 3834
rect 81290 3782 111766 3834
rect 111818 3782 111830 3834
rect 111882 3782 111894 3834
rect 111946 3782 111958 3834
rect 112010 3782 142486 3834
rect 142538 3782 142550 3834
rect 142602 3782 142614 3834
rect 142666 3782 142678 3834
rect 142730 3782 173206 3834
rect 173258 3782 173270 3834
rect 173322 3782 173334 3834
rect 173386 3782 173398 3834
rect 173450 3782 178848 3834
rect 1104 3760 178848 3782
rect 3142 3720 3148 3732
rect 3103 3692 3148 3720
rect 3142 3680 3148 3692
rect 3200 3680 3206 3732
rect 6273 3723 6331 3729
rect 6273 3689 6285 3723
rect 6319 3720 6331 3723
rect 10229 3723 10287 3729
rect 10229 3720 10241 3723
rect 6319 3692 10241 3720
rect 6319 3689 6331 3692
rect 6273 3683 6331 3689
rect 10229 3689 10241 3692
rect 10275 3689 10287 3723
rect 10229 3683 10287 3689
rect 11149 3723 11207 3729
rect 11149 3689 11161 3723
rect 11195 3720 11207 3723
rect 24673 3723 24731 3729
rect 24673 3720 24685 3723
rect 11195 3692 24685 3720
rect 11195 3689 11207 3692
rect 11149 3683 11207 3689
rect 24673 3689 24685 3692
rect 24719 3689 24731 3723
rect 33134 3720 33140 3732
rect 24673 3683 24731 3689
rect 27080 3692 33140 3720
rect 1673 3655 1731 3661
rect 1673 3621 1685 3655
rect 1719 3652 1731 3655
rect 1946 3652 1952 3664
rect 1719 3624 1952 3652
rect 1719 3621 1731 3624
rect 1673 3615 1731 3621
rect 1946 3612 1952 3624
rect 2004 3612 2010 3664
rect 9950 3612 9956 3664
rect 10008 3652 10014 3664
rect 12250 3652 12256 3664
rect 10008 3624 12112 3652
rect 12211 3624 12256 3652
rect 10008 3612 10014 3624
rect 2501 3587 2559 3593
rect 2501 3553 2513 3587
rect 2547 3553 2559 3587
rect 3326 3584 3332 3596
rect 3287 3556 3332 3584
rect 2501 3547 2559 3553
rect 1486 3476 1492 3528
rect 1544 3516 1550 3528
rect 2516 3516 2544 3547
rect 3326 3544 3332 3556
rect 3384 3544 3390 3596
rect 4798 3544 4804 3596
rect 4856 3584 4862 3596
rect 4985 3587 5043 3593
rect 4985 3584 4997 3587
rect 4856 3556 4997 3584
rect 4856 3544 4862 3556
rect 4985 3553 4997 3556
rect 5031 3553 5043 3587
rect 4985 3547 5043 3553
rect 6270 3544 6276 3596
rect 6328 3584 6334 3596
rect 6457 3587 6515 3593
rect 6457 3584 6469 3587
rect 6328 3556 6469 3584
rect 6328 3544 6334 3556
rect 6457 3553 6469 3556
rect 6503 3553 6515 3587
rect 9582 3584 9588 3596
rect 9543 3556 9588 3584
rect 6457 3547 6515 3553
rect 9582 3544 9588 3556
rect 9640 3544 9646 3596
rect 10318 3584 10324 3596
rect 10279 3556 10324 3584
rect 10318 3544 10324 3556
rect 10376 3544 10382 3596
rect 10686 3544 10692 3596
rect 10744 3584 10750 3596
rect 10965 3587 11023 3593
rect 10965 3584 10977 3587
rect 10744 3556 10977 3584
rect 10744 3544 10750 3556
rect 10965 3553 10977 3556
rect 11011 3553 11023 3587
rect 12084 3584 12112 3624
rect 12250 3612 12256 3624
rect 12308 3612 12314 3664
rect 12342 3612 12348 3664
rect 12400 3652 12406 3664
rect 13722 3652 13728 3664
rect 12400 3624 13584 3652
rect 13683 3624 13728 3652
rect 12400 3612 12406 3624
rect 13354 3584 13360 3596
rect 12084 3556 13360 3584
rect 10965 3547 11023 3553
rect 13354 3544 13360 3556
rect 13412 3544 13418 3596
rect 13556 3593 13584 3624
rect 13722 3612 13728 3624
rect 13780 3612 13786 3664
rect 14826 3652 14832 3664
rect 14787 3624 14832 3652
rect 14826 3612 14832 3624
rect 14884 3612 14890 3664
rect 15396 3624 15608 3652
rect 13541 3587 13599 3593
rect 13541 3553 13553 3587
rect 13587 3553 13599 3587
rect 13541 3547 13599 3553
rect 14185 3587 14243 3593
rect 14185 3553 14197 3587
rect 14231 3584 14243 3587
rect 15396 3584 15424 3624
rect 14231 3556 15424 3584
rect 15473 3587 15531 3593
rect 14231 3553 14243 3556
rect 14185 3547 14243 3553
rect 15473 3553 15485 3587
rect 15519 3553 15531 3587
rect 15580 3584 15608 3624
rect 15654 3612 15660 3664
rect 15712 3652 15718 3664
rect 18874 3652 18880 3664
rect 15712 3624 18736 3652
rect 18835 3624 18880 3652
rect 15712 3612 15718 3624
rect 16574 3584 16580 3596
rect 15580 3556 16580 3584
rect 15473 3547 15531 3553
rect 10134 3516 10140 3528
rect 1544 3488 2544 3516
rect 6886 3488 10140 3516
rect 1544 3476 1550 3488
rect 750 3408 756 3460
rect 808 3448 814 3460
rect 1765 3451 1823 3457
rect 1765 3448 1777 3451
rect 808 3420 1777 3448
rect 808 3408 814 3420
rect 1765 3417 1777 3420
rect 1811 3417 1823 3451
rect 1765 3411 1823 3417
rect 4801 3451 4859 3457
rect 4801 3417 4813 3451
rect 4847 3448 4859 3451
rect 6886 3448 6914 3488
rect 10134 3476 10140 3488
rect 10192 3476 10198 3528
rect 14734 3476 14740 3528
rect 14792 3516 14798 3528
rect 15488 3516 15516 3547
rect 16574 3544 16580 3556
rect 16632 3544 16638 3596
rect 16669 3587 16727 3593
rect 16669 3553 16681 3587
rect 16715 3553 16727 3587
rect 16669 3547 16727 3553
rect 14792 3488 15516 3516
rect 16684 3516 16712 3547
rect 16758 3544 16764 3596
rect 16816 3584 16822 3596
rect 16853 3587 16911 3593
rect 16853 3584 16865 3587
rect 16816 3556 16865 3584
rect 16816 3544 16822 3556
rect 16853 3553 16865 3556
rect 16899 3553 16911 3587
rect 16853 3547 16911 3553
rect 16942 3544 16948 3596
rect 17000 3584 17006 3596
rect 17313 3587 17371 3593
rect 17313 3584 17325 3587
rect 17000 3556 17325 3584
rect 17000 3544 17006 3556
rect 17313 3553 17325 3556
rect 17359 3553 17371 3587
rect 18046 3584 18052 3596
rect 18007 3556 18052 3584
rect 17313 3547 17371 3553
rect 18046 3544 18052 3556
rect 18104 3544 18110 3596
rect 18708 3584 18736 3624
rect 18874 3612 18880 3624
rect 18932 3612 18938 3664
rect 21085 3655 21143 3661
rect 19076 3624 21036 3652
rect 19076 3584 19104 3624
rect 18708 3556 19104 3584
rect 19150 3544 19156 3596
rect 19208 3584 19214 3596
rect 19981 3587 20039 3593
rect 19981 3584 19993 3587
rect 19208 3556 19993 3584
rect 19208 3544 19214 3556
rect 19981 3553 19993 3556
rect 20027 3553 20039 3587
rect 21008 3584 21036 3624
rect 21085 3621 21097 3655
rect 21131 3652 21143 3655
rect 27080 3652 27108 3692
rect 33134 3680 33140 3692
rect 33192 3680 33198 3732
rect 33226 3680 33232 3732
rect 33284 3720 33290 3732
rect 45462 3720 45468 3732
rect 33284 3692 45468 3720
rect 33284 3680 33290 3692
rect 45462 3680 45468 3692
rect 45520 3680 45526 3732
rect 70670 3720 70676 3732
rect 67192 3692 70676 3720
rect 21131 3624 24256 3652
rect 21131 3621 21143 3624
rect 21085 3615 21143 3621
rect 21266 3584 21272 3596
rect 21008 3556 21272 3584
rect 19981 3547 20039 3553
rect 21266 3544 21272 3556
rect 21324 3544 21330 3596
rect 21358 3544 21364 3596
rect 21416 3584 21422 3596
rect 21729 3587 21787 3593
rect 21729 3584 21741 3587
rect 21416 3556 21741 3584
rect 21416 3544 21422 3556
rect 21729 3553 21741 3556
rect 21775 3553 21787 3587
rect 22462 3584 22468 3596
rect 22423 3556 22468 3584
rect 21729 3547 21787 3553
rect 22462 3544 22468 3556
rect 22520 3544 22526 3596
rect 23566 3584 23572 3596
rect 23527 3556 23572 3584
rect 23566 3544 23572 3556
rect 23624 3544 23630 3596
rect 24228 3584 24256 3624
rect 24596 3624 27108 3652
rect 24596 3584 24624 3624
rect 28810 3612 28816 3664
rect 28868 3652 28874 3664
rect 40034 3652 40040 3664
rect 28868 3624 40040 3652
rect 28868 3612 28874 3624
rect 40034 3612 40040 3624
rect 40092 3612 40098 3664
rect 41414 3612 41420 3664
rect 41472 3652 41478 3664
rect 62206 3652 62212 3664
rect 41472 3624 62212 3652
rect 41472 3612 41478 3624
rect 62206 3612 62212 3624
rect 62264 3612 62270 3664
rect 67192 3661 67220 3692
rect 70670 3680 70676 3692
rect 70728 3680 70734 3732
rect 70762 3680 70768 3732
rect 70820 3720 70826 3732
rect 72694 3720 72700 3732
rect 70820 3692 72700 3720
rect 70820 3680 70826 3692
rect 72694 3680 72700 3692
rect 72752 3680 72758 3732
rect 72789 3723 72847 3729
rect 72789 3689 72801 3723
rect 72835 3720 72847 3723
rect 73246 3720 73252 3732
rect 72835 3692 73252 3720
rect 72835 3689 72847 3692
rect 72789 3683 72847 3689
rect 73246 3680 73252 3692
rect 73304 3680 73310 3732
rect 75181 3723 75239 3729
rect 75181 3689 75193 3723
rect 75227 3720 75239 3723
rect 75270 3720 75276 3732
rect 75227 3692 75276 3720
rect 75227 3689 75239 3692
rect 75181 3683 75239 3689
rect 75270 3680 75276 3692
rect 75328 3680 75334 3732
rect 75822 3680 75828 3732
rect 75880 3720 75886 3732
rect 79042 3720 79048 3732
rect 75880 3692 79048 3720
rect 75880 3680 75886 3692
rect 79042 3680 79048 3692
rect 79100 3680 79106 3732
rect 79410 3720 79416 3732
rect 79371 3692 79416 3720
rect 79410 3680 79416 3692
rect 79468 3680 79474 3732
rect 80054 3680 80060 3732
rect 80112 3720 80118 3732
rect 80112 3692 80560 3720
rect 80112 3680 80118 3692
rect 67177 3655 67235 3661
rect 67177 3621 67189 3655
rect 67223 3621 67235 3655
rect 67177 3615 67235 3621
rect 67591 3655 67649 3661
rect 67591 3621 67603 3655
rect 67637 3652 67649 3655
rect 68278 3652 68284 3664
rect 67637 3624 68140 3652
rect 68239 3624 68284 3652
rect 67637 3621 67649 3624
rect 67591 3615 67649 3621
rect 24228 3556 24624 3584
rect 24670 3544 24676 3596
rect 24728 3584 24734 3596
rect 25225 3587 25283 3593
rect 25225 3584 25237 3587
rect 24728 3556 25237 3584
rect 24728 3544 24734 3556
rect 25225 3553 25237 3556
rect 25271 3553 25283 3587
rect 25225 3547 25283 3553
rect 25774 3544 25780 3596
rect 25832 3584 25838 3596
rect 25869 3587 25927 3593
rect 25869 3584 25881 3587
rect 25832 3556 25881 3584
rect 25832 3544 25838 3556
rect 25869 3553 25881 3556
rect 25915 3553 25927 3587
rect 26878 3584 26884 3596
rect 26839 3556 26884 3584
rect 25869 3547 25927 3553
rect 26878 3544 26884 3556
rect 26936 3544 26942 3596
rect 27982 3584 27988 3596
rect 27943 3556 27988 3584
rect 27982 3544 27988 3556
rect 28040 3544 28046 3596
rect 28166 3544 28172 3596
rect 28224 3584 28230 3596
rect 30374 3584 30380 3596
rect 28224 3556 30380 3584
rect 28224 3544 28230 3556
rect 30374 3544 30380 3556
rect 30432 3544 30438 3596
rect 31294 3584 31300 3596
rect 31255 3556 31300 3584
rect 31294 3544 31300 3556
rect 31352 3544 31358 3596
rect 32398 3584 32404 3596
rect 32359 3556 32404 3584
rect 32398 3544 32404 3556
rect 32456 3544 32462 3596
rect 33502 3584 33508 3596
rect 33463 3556 33508 3584
rect 33502 3544 33508 3556
rect 33560 3544 33566 3596
rect 34606 3584 34612 3596
rect 34567 3556 34612 3584
rect 34606 3544 34612 3556
rect 34664 3544 34670 3596
rect 35710 3584 35716 3596
rect 35671 3556 35716 3584
rect 35710 3544 35716 3556
rect 35768 3544 35774 3596
rect 37458 3584 37464 3596
rect 36280 3556 37464 3584
rect 21542 3516 21548 3528
rect 16684 3488 21548 3516
rect 14792 3476 14798 3488
rect 21542 3476 21548 3488
rect 21600 3476 21606 3528
rect 22278 3476 22284 3528
rect 22336 3516 22342 3528
rect 24118 3516 24124 3528
rect 22336 3488 24124 3516
rect 22336 3476 22342 3488
rect 24118 3476 24124 3488
rect 24176 3476 24182 3528
rect 25314 3476 25320 3528
rect 25372 3516 25378 3528
rect 36280 3516 36308 3556
rect 37458 3544 37464 3556
rect 37516 3544 37522 3596
rect 37918 3584 37924 3596
rect 37879 3556 37924 3584
rect 37918 3544 37924 3556
rect 37976 3544 37982 3596
rect 38194 3544 38200 3596
rect 38252 3584 38258 3596
rect 39574 3584 39580 3596
rect 38252 3556 39580 3584
rect 38252 3544 38258 3556
rect 39574 3544 39580 3556
rect 39632 3544 39638 3596
rect 39758 3584 39764 3596
rect 39719 3556 39764 3584
rect 39758 3544 39764 3556
rect 39816 3544 39822 3596
rect 40862 3544 40868 3596
rect 40920 3584 40926 3596
rect 40957 3587 41015 3593
rect 40957 3584 40969 3587
rect 40920 3556 40969 3584
rect 40920 3544 40926 3556
rect 40957 3553 40969 3556
rect 41003 3553 41015 3587
rect 41966 3584 41972 3596
rect 41927 3556 41972 3584
rect 40957 3547 41015 3553
rect 41966 3544 41972 3556
rect 42024 3544 42030 3596
rect 43070 3584 43076 3596
rect 43031 3556 43076 3584
rect 43070 3544 43076 3556
rect 43128 3544 43134 3596
rect 44174 3584 44180 3596
rect 44135 3556 44180 3584
rect 44174 3544 44180 3556
rect 44232 3544 44238 3596
rect 45097 3587 45155 3593
rect 45097 3553 45109 3587
rect 45143 3584 45155 3587
rect 45278 3584 45284 3596
rect 45143 3556 45284 3584
rect 45143 3553 45155 3556
rect 45097 3547 45155 3553
rect 45278 3544 45284 3556
rect 45336 3544 45342 3596
rect 46382 3584 46388 3596
rect 46343 3556 46388 3584
rect 46382 3544 46388 3556
rect 46440 3544 46446 3596
rect 47486 3584 47492 3596
rect 47447 3556 47492 3584
rect 47486 3544 47492 3556
rect 47544 3544 47550 3596
rect 48590 3584 48596 3596
rect 48551 3556 48596 3584
rect 48590 3544 48596 3556
rect 48648 3544 48654 3596
rect 49694 3584 49700 3596
rect 49655 3556 49700 3584
rect 49694 3544 49700 3556
rect 49752 3544 49758 3596
rect 54110 3584 54116 3596
rect 54071 3556 54116 3584
rect 54110 3544 54116 3556
rect 54168 3544 54174 3596
rect 55214 3584 55220 3596
rect 55175 3556 55220 3584
rect 55214 3544 55220 3556
rect 55272 3544 55278 3596
rect 56318 3544 56324 3596
rect 56376 3584 56382 3596
rect 56689 3587 56747 3593
rect 56689 3584 56701 3587
rect 56376 3556 56701 3584
rect 56376 3544 56382 3556
rect 56689 3553 56701 3556
rect 56735 3553 56747 3587
rect 57422 3584 57428 3596
rect 57383 3556 57428 3584
rect 56689 3547 56747 3553
rect 57422 3544 57428 3556
rect 57480 3544 57486 3596
rect 58526 3584 58532 3596
rect 58487 3556 58532 3584
rect 58526 3544 58532 3556
rect 58584 3544 58590 3596
rect 59630 3584 59636 3596
rect 59591 3556 59636 3584
rect 59630 3544 59636 3556
rect 59688 3544 59694 3596
rect 60642 3584 60648 3596
rect 60603 3556 60648 3584
rect 60642 3544 60648 3556
rect 60700 3544 60706 3596
rect 61746 3544 61752 3596
rect 61804 3584 61810 3596
rect 61933 3587 61991 3593
rect 61933 3584 61945 3587
rect 61804 3556 61945 3584
rect 61804 3544 61810 3556
rect 61933 3553 61945 3556
rect 61979 3553 61991 3587
rect 62850 3584 62856 3596
rect 62811 3556 62856 3584
rect 61933 3547 61991 3553
rect 62850 3544 62856 3556
rect 62908 3544 62914 3596
rect 63954 3584 63960 3596
rect 63915 3556 63960 3584
rect 63954 3544 63960 3556
rect 64012 3544 64018 3596
rect 65058 3584 65064 3596
rect 65019 3556 65064 3584
rect 65058 3544 65064 3556
rect 65116 3544 65122 3596
rect 66073 3587 66131 3593
rect 66073 3553 66085 3587
rect 66119 3584 66131 3587
rect 66530 3584 66536 3596
rect 66119 3556 66536 3584
rect 66119 3553 66131 3556
rect 66073 3547 66131 3553
rect 66530 3544 66536 3556
rect 66588 3544 66594 3596
rect 67726 3544 67732 3596
rect 67784 3584 67790 3596
rect 67821 3587 67879 3593
rect 67821 3584 67833 3587
rect 67784 3556 67833 3584
rect 67784 3544 67790 3556
rect 67821 3553 67833 3556
rect 67867 3553 67879 3587
rect 68112 3584 68140 3624
rect 68278 3612 68284 3624
rect 68336 3612 68342 3664
rect 68695 3655 68753 3661
rect 68695 3621 68707 3655
rect 68741 3652 68753 3655
rect 69658 3652 69664 3664
rect 68741 3624 69664 3652
rect 68741 3621 68753 3624
rect 68695 3615 68753 3621
rect 69658 3612 69664 3624
rect 69716 3612 69722 3664
rect 69842 3661 69848 3664
rect 69799 3655 69848 3661
rect 69799 3621 69811 3655
rect 69845 3621 69848 3655
rect 69799 3615 69848 3621
rect 69842 3612 69848 3615
rect 69900 3612 69906 3664
rect 69934 3612 69940 3664
rect 69992 3652 69998 3664
rect 72418 3652 72424 3664
rect 69992 3624 72424 3652
rect 69992 3612 69998 3624
rect 72418 3612 72424 3624
rect 72476 3612 72482 3664
rect 76282 3612 76288 3664
rect 76340 3652 76346 3664
rect 76340 3624 76385 3652
rect 76340 3612 76346 3624
rect 76742 3612 76748 3664
rect 76800 3652 76806 3664
rect 80422 3652 80428 3664
rect 76800 3624 80284 3652
rect 80383 3624 80428 3652
rect 76800 3612 76806 3624
rect 69106 3584 69112 3596
rect 68112 3556 69112 3584
rect 67821 3547 67879 3553
rect 69106 3544 69112 3556
rect 69164 3544 69170 3596
rect 69382 3544 69388 3596
rect 69440 3593 69446 3596
rect 69440 3584 69452 3593
rect 69440 3556 69485 3584
rect 69440 3547 69452 3556
rect 69440 3544 69446 3547
rect 69566 3544 69572 3596
rect 69624 3584 69630 3596
rect 70489 3587 70547 3593
rect 70489 3584 70501 3587
rect 69624 3556 70501 3584
rect 69624 3544 69630 3556
rect 70489 3553 70501 3556
rect 70535 3553 70547 3587
rect 70489 3547 70547 3553
rect 70854 3544 70860 3596
rect 70912 3584 70918 3596
rect 71133 3587 71191 3593
rect 71133 3584 71145 3587
rect 70912 3556 71145 3584
rect 70912 3544 70918 3556
rect 71133 3553 71145 3556
rect 71179 3584 71191 3587
rect 71222 3584 71228 3596
rect 71179 3556 71228 3584
rect 71179 3553 71191 3556
rect 71133 3547 71191 3553
rect 71222 3544 71228 3556
rect 71280 3544 71286 3596
rect 73430 3584 73436 3596
rect 73391 3556 73436 3584
rect 73430 3544 73436 3556
rect 73488 3544 73494 3596
rect 74353 3587 74411 3593
rect 74353 3553 74365 3587
rect 74399 3584 74411 3587
rect 75730 3584 75736 3596
rect 74399 3556 75736 3584
rect 74399 3553 74411 3556
rect 74353 3547 74411 3553
rect 75730 3544 75736 3556
rect 75788 3544 75794 3596
rect 76006 3544 76012 3596
rect 76064 3584 76070 3596
rect 78214 3584 78220 3596
rect 76064 3556 78220 3584
rect 76064 3544 76070 3556
rect 78214 3544 78220 3556
rect 78272 3584 78278 3596
rect 78309 3587 78367 3593
rect 78309 3584 78321 3587
rect 78272 3556 78321 3584
rect 78272 3544 78278 3556
rect 78309 3553 78321 3556
rect 78355 3553 78367 3587
rect 80054 3584 80060 3596
rect 78309 3547 78367 3553
rect 78416 3556 80060 3584
rect 25372 3488 36308 3516
rect 25372 3476 25378 3488
rect 36446 3476 36452 3528
rect 36504 3516 36510 3528
rect 45002 3516 45008 3528
rect 36504 3488 45008 3516
rect 36504 3476 36510 3488
rect 45002 3476 45008 3488
rect 45060 3476 45066 3528
rect 72421 3519 72479 3525
rect 72421 3485 72433 3519
rect 72467 3516 72479 3519
rect 75822 3516 75828 3528
rect 72467 3488 75828 3516
rect 72467 3485 72479 3488
rect 72421 3479 72479 3485
rect 75822 3476 75828 3488
rect 75880 3476 75886 3528
rect 75917 3519 75975 3525
rect 75917 3485 75929 3519
rect 75963 3516 75975 3519
rect 78416 3516 78444 3556
rect 80054 3544 80060 3556
rect 80112 3544 80118 3596
rect 80256 3584 80284 3624
rect 80422 3612 80428 3624
rect 80480 3612 80486 3664
rect 80532 3652 80560 3692
rect 80606 3680 80612 3732
rect 80664 3720 80670 3732
rect 81069 3723 81127 3729
rect 80664 3692 80709 3720
rect 80664 3680 80670 3692
rect 81069 3689 81081 3723
rect 81115 3720 81127 3723
rect 81434 3720 81440 3732
rect 81115 3692 81440 3720
rect 81115 3689 81127 3692
rect 81069 3683 81127 3689
rect 81434 3680 81440 3692
rect 81492 3680 81498 3732
rect 81802 3720 81808 3732
rect 81636 3692 81808 3720
rect 81636 3652 81664 3692
rect 81802 3680 81808 3692
rect 81860 3680 81866 3732
rect 81897 3723 81955 3729
rect 81897 3689 81909 3723
rect 81943 3720 81955 3723
rect 83458 3720 83464 3732
rect 81943 3692 83464 3720
rect 81943 3689 81955 3692
rect 81897 3683 81955 3689
rect 83458 3680 83464 3692
rect 83516 3680 83522 3732
rect 85022 3720 85028 3732
rect 84028 3692 84884 3720
rect 84983 3692 85028 3720
rect 82170 3652 82176 3664
rect 80532 3624 81664 3652
rect 81728 3624 82176 3652
rect 80974 3584 80980 3596
rect 80256 3556 80980 3584
rect 80974 3544 80980 3556
rect 81032 3544 81038 3596
rect 81069 3587 81127 3593
rect 81069 3553 81081 3587
rect 81115 3584 81127 3587
rect 81165 3587 81223 3593
rect 81165 3584 81177 3587
rect 81115 3556 81177 3584
rect 81115 3553 81127 3556
rect 81069 3547 81127 3553
rect 81165 3553 81177 3556
rect 81211 3553 81223 3587
rect 81165 3547 81223 3553
rect 81345 3587 81403 3593
rect 81345 3553 81357 3587
rect 81391 3553 81403 3587
rect 81345 3547 81403 3553
rect 81437 3587 81495 3593
rect 81437 3553 81449 3587
rect 81483 3584 81495 3587
rect 81526 3584 81532 3596
rect 81483 3556 81532 3584
rect 81483 3553 81495 3556
rect 81437 3547 81495 3553
rect 75963 3488 78444 3516
rect 78493 3519 78551 3525
rect 75963 3485 75975 3488
rect 75917 3479 75975 3485
rect 78493 3485 78505 3519
rect 78539 3516 78551 3519
rect 80882 3516 80888 3528
rect 78539 3488 80888 3516
rect 78539 3485 78551 3488
rect 78493 3479 78551 3485
rect 80882 3476 80888 3488
rect 80940 3476 80946 3528
rect 4847 3420 6914 3448
rect 9769 3451 9827 3457
rect 4847 3417 4859 3420
rect 4801 3411 4859 3417
rect 9769 3417 9781 3451
rect 9815 3448 9827 3451
rect 22002 3448 22008 3460
rect 9815 3420 22008 3448
rect 9815 3417 9827 3420
rect 9769 3411 9827 3417
rect 22002 3408 22008 3420
rect 22060 3408 22066 3460
rect 24673 3451 24731 3457
rect 24673 3417 24685 3451
rect 24719 3448 24731 3451
rect 35342 3448 35348 3460
rect 24719 3420 35348 3448
rect 24719 3417 24731 3420
rect 24673 3411 24731 3417
rect 35342 3408 35348 3420
rect 35400 3408 35406 3460
rect 35434 3408 35440 3460
rect 35492 3448 35498 3460
rect 46198 3448 46204 3460
rect 35492 3420 46204 3448
rect 35492 3408 35498 3420
rect 46198 3408 46204 3420
rect 46256 3408 46262 3460
rect 61562 3408 61568 3460
rect 61620 3448 61626 3460
rect 68833 3451 68891 3457
rect 68833 3448 68845 3451
rect 61620 3420 68845 3448
rect 61620 3408 61626 3420
rect 68833 3417 68845 3420
rect 68879 3417 68891 3451
rect 68833 3411 68891 3417
rect 72694 3408 72700 3460
rect 72752 3448 72758 3460
rect 74718 3448 74724 3460
rect 72752 3420 74724 3448
rect 72752 3408 72758 3420
rect 74718 3408 74724 3420
rect 74776 3408 74782 3460
rect 74813 3451 74871 3457
rect 74813 3417 74825 3451
rect 74859 3448 74871 3451
rect 78858 3448 78864 3460
rect 74859 3420 78864 3448
rect 74859 3417 74871 3420
rect 74813 3411 74871 3417
rect 78858 3408 78864 3420
rect 78916 3408 78922 3460
rect 79042 3448 79048 3460
rect 79003 3420 79048 3448
rect 79042 3408 79048 3420
rect 79100 3408 79106 3460
rect 79226 3408 79232 3460
rect 79284 3448 79290 3460
rect 79597 3451 79655 3457
rect 79597 3448 79609 3451
rect 79284 3420 79609 3448
rect 79284 3408 79290 3420
rect 79597 3417 79609 3420
rect 79643 3417 79655 3451
rect 79597 3411 79655 3417
rect 80057 3451 80115 3457
rect 80057 3417 80069 3451
rect 80103 3448 80115 3451
rect 80103 3420 80560 3448
rect 80103 3417 80115 3420
rect 80057 3411 80115 3417
rect 2682 3380 2688 3392
rect 2643 3352 2688 3380
rect 2682 3340 2688 3352
rect 2740 3340 2746 3392
rect 10229 3383 10287 3389
rect 10229 3349 10241 3383
rect 10275 3380 10287 3383
rect 11974 3380 11980 3392
rect 10275 3352 11980 3380
rect 10275 3349 10287 3352
rect 10229 3343 10287 3349
rect 11974 3340 11980 3352
rect 12032 3340 12038 3392
rect 12158 3340 12164 3392
rect 12216 3380 12222 3392
rect 12345 3383 12403 3389
rect 12345 3380 12357 3383
rect 12216 3352 12357 3380
rect 12216 3340 12222 3352
rect 12345 3349 12357 3352
rect 12391 3349 12403 3383
rect 12345 3343 12403 3349
rect 13078 3340 13084 3392
rect 13136 3380 13142 3392
rect 14185 3383 14243 3389
rect 14185 3380 14197 3383
rect 13136 3352 14197 3380
rect 13136 3340 13142 3352
rect 14185 3349 14197 3352
rect 14231 3349 14243 3383
rect 14185 3343 14243 3349
rect 14366 3340 14372 3392
rect 14424 3380 14430 3392
rect 14921 3383 14979 3389
rect 14921 3380 14933 3383
rect 14424 3352 14933 3380
rect 14424 3340 14430 3352
rect 14921 3349 14933 3352
rect 14967 3349 14979 3383
rect 14921 3343 14979 3349
rect 15378 3340 15384 3392
rect 15436 3380 15442 3392
rect 18690 3380 18696 3392
rect 15436 3352 18696 3380
rect 15436 3340 15442 3352
rect 18690 3340 18696 3352
rect 18748 3340 18754 3392
rect 18782 3340 18788 3392
rect 18840 3380 18846 3392
rect 18969 3383 19027 3389
rect 18969 3380 18981 3383
rect 18840 3352 18981 3380
rect 18840 3340 18846 3352
rect 18969 3349 18981 3352
rect 19015 3349 19027 3383
rect 18969 3343 19027 3349
rect 19058 3340 19064 3392
rect 19116 3380 19122 3392
rect 20898 3380 20904 3392
rect 19116 3352 20904 3380
rect 19116 3340 19122 3352
rect 20898 3340 20904 3352
rect 20956 3340 20962 3392
rect 20990 3340 20996 3392
rect 21048 3380 21054 3392
rect 21177 3383 21235 3389
rect 21177 3380 21189 3383
rect 21048 3352 21189 3380
rect 21048 3340 21054 3352
rect 21177 3349 21189 3352
rect 21223 3349 21235 3383
rect 21177 3343 21235 3349
rect 22646 3340 22652 3392
rect 22704 3380 22710 3392
rect 34238 3380 34244 3392
rect 22704 3352 34244 3380
rect 22704 3340 22710 3352
rect 34238 3340 34244 3352
rect 34296 3340 34302 3392
rect 34330 3340 34336 3392
rect 34388 3380 34394 3392
rect 45370 3380 45376 3392
rect 34388 3352 45376 3380
rect 34388 3340 34394 3352
rect 45370 3340 45376 3352
rect 45428 3340 45434 3392
rect 67542 3380 67548 3392
rect 67455 3352 67548 3380
rect 67542 3340 67548 3352
rect 67600 3380 67606 3392
rect 68649 3383 68707 3389
rect 68649 3380 68661 3383
rect 67600 3352 68661 3380
rect 67600 3340 67606 3352
rect 68649 3349 68661 3352
rect 68695 3380 68707 3383
rect 69750 3380 69756 3392
rect 68695 3352 69756 3380
rect 68695 3349 68707 3352
rect 68649 3343 68707 3349
rect 69750 3340 69756 3352
rect 69808 3340 69814 3392
rect 69937 3383 69995 3389
rect 69937 3349 69949 3383
rect 69983 3380 69995 3383
rect 70026 3380 70032 3392
rect 69983 3352 70032 3380
rect 69983 3349 69995 3352
rect 69937 3343 69995 3349
rect 70026 3340 70032 3352
rect 70084 3340 70090 3392
rect 70486 3340 70492 3392
rect 70544 3380 70550 3392
rect 71222 3380 71228 3392
rect 70544 3352 71228 3380
rect 70544 3340 70550 3352
rect 71222 3340 71228 3352
rect 71280 3340 71286 3392
rect 71317 3383 71375 3389
rect 71317 3349 71329 3383
rect 71363 3380 71375 3383
rect 72326 3380 72332 3392
rect 71363 3352 72332 3380
rect 71363 3349 71375 3352
rect 71317 3343 71375 3349
rect 72326 3340 72332 3352
rect 72384 3380 72390 3392
rect 72789 3383 72847 3389
rect 72789 3380 72801 3383
rect 72384 3352 72801 3380
rect 72384 3340 72390 3352
rect 72789 3349 72801 3352
rect 72835 3349 72847 3383
rect 72970 3380 72976 3392
rect 72931 3352 72976 3380
rect 72789 3343 72847 3349
rect 72970 3340 72976 3352
rect 73028 3340 73034 3392
rect 73617 3383 73675 3389
rect 73617 3349 73629 3383
rect 73663 3380 73675 3383
rect 75086 3380 75092 3392
rect 73663 3352 75092 3380
rect 73663 3349 73675 3352
rect 73617 3343 73675 3349
rect 75086 3340 75092 3352
rect 75144 3380 75150 3392
rect 75181 3383 75239 3389
rect 75181 3380 75193 3383
rect 75144 3352 75193 3380
rect 75144 3340 75150 3352
rect 75181 3349 75193 3352
rect 75227 3349 75239 3383
rect 75181 3343 75239 3349
rect 75270 3340 75276 3392
rect 75328 3380 75334 3392
rect 75365 3383 75423 3389
rect 75365 3380 75377 3383
rect 75328 3352 75377 3380
rect 75328 3340 75334 3352
rect 75365 3349 75377 3352
rect 75411 3349 75423 3383
rect 76282 3380 76288 3392
rect 76243 3352 76288 3380
rect 75365 3343 75423 3349
rect 76282 3340 76288 3352
rect 76340 3340 76346 3392
rect 76469 3383 76527 3389
rect 76469 3349 76481 3383
rect 76515 3380 76527 3383
rect 76650 3380 76656 3392
rect 76515 3352 76656 3380
rect 76515 3349 76527 3352
rect 76469 3343 76527 3349
rect 76650 3340 76656 3352
rect 76708 3340 76714 3392
rect 77846 3340 77852 3392
rect 77904 3380 77910 3392
rect 79318 3380 79324 3392
rect 77904 3352 79324 3380
rect 77904 3340 77910 3352
rect 79318 3340 79324 3352
rect 79376 3380 79382 3392
rect 79413 3383 79471 3389
rect 79413 3380 79425 3383
rect 79376 3352 79425 3380
rect 79376 3340 79382 3352
rect 79413 3349 79425 3352
rect 79459 3380 79471 3383
rect 80425 3383 80483 3389
rect 80425 3380 80437 3383
rect 79459 3352 80437 3380
rect 79459 3349 79471 3352
rect 79413 3343 79471 3349
rect 80425 3349 80437 3352
rect 80471 3349 80483 3383
rect 80532 3380 80560 3420
rect 80606 3408 80612 3460
rect 80664 3448 80670 3460
rect 81360 3448 81388 3547
rect 81526 3544 81532 3556
rect 81584 3544 81590 3596
rect 81728 3593 81756 3624
rect 82170 3612 82176 3624
rect 82228 3612 82234 3664
rect 82354 3612 82360 3664
rect 82412 3652 82418 3664
rect 84028 3652 84056 3692
rect 82412 3624 84056 3652
rect 82412 3612 82418 3624
rect 81713 3587 81771 3593
rect 81713 3553 81725 3587
rect 81759 3553 81771 3587
rect 81713 3547 81771 3553
rect 81728 3516 81756 3547
rect 81802 3544 81808 3596
rect 81860 3584 81866 3596
rect 82909 3587 82967 3593
rect 82909 3584 82921 3587
rect 81860 3556 82921 3584
rect 81860 3544 81866 3556
rect 82909 3553 82921 3556
rect 82955 3553 82967 3587
rect 82909 3547 82967 3553
rect 83093 3587 83151 3593
rect 83093 3553 83105 3587
rect 83139 3553 83151 3587
rect 83093 3547 83151 3553
rect 83461 3587 83519 3593
rect 83461 3553 83473 3587
rect 83507 3584 83519 3587
rect 84102 3584 84108 3596
rect 83507 3556 84108 3584
rect 83507 3553 83519 3556
rect 83461 3547 83519 3553
rect 81452 3488 81756 3516
rect 81452 3460 81480 3488
rect 81894 3476 81900 3528
rect 81952 3516 81958 3528
rect 83108 3516 83136 3547
rect 84102 3544 84108 3556
rect 84160 3544 84166 3596
rect 84289 3587 84347 3593
rect 84289 3553 84301 3587
rect 84335 3584 84347 3587
rect 84378 3584 84384 3596
rect 84335 3556 84384 3584
rect 84335 3553 84347 3556
rect 84289 3547 84347 3553
rect 84378 3544 84384 3556
rect 84436 3544 84442 3596
rect 84856 3593 84884 3692
rect 85022 3680 85028 3692
rect 85080 3680 85086 3732
rect 85758 3680 85764 3732
rect 85816 3720 85822 3732
rect 86221 3723 86279 3729
rect 86221 3720 86233 3723
rect 85816 3692 86233 3720
rect 85816 3680 85822 3692
rect 86221 3689 86233 3692
rect 86267 3689 86279 3723
rect 86221 3683 86279 3689
rect 87233 3723 87291 3729
rect 87233 3689 87245 3723
rect 87279 3720 87291 3723
rect 87322 3720 87328 3732
rect 87279 3692 87328 3720
rect 87279 3689 87291 3692
rect 87233 3683 87291 3689
rect 87322 3680 87328 3692
rect 87380 3680 87386 3732
rect 88521 3723 88579 3729
rect 88521 3689 88533 3723
rect 88567 3720 88579 3723
rect 88702 3720 88708 3732
rect 88567 3692 88708 3720
rect 88567 3689 88579 3692
rect 88521 3683 88579 3689
rect 88702 3680 88708 3692
rect 88760 3680 88766 3732
rect 88886 3680 88892 3732
rect 88944 3720 88950 3732
rect 91005 3723 91063 3729
rect 91005 3720 91017 3723
rect 88944 3692 91017 3720
rect 88944 3680 88950 3692
rect 91005 3689 91017 3692
rect 91051 3689 91063 3723
rect 91646 3720 91652 3732
rect 91607 3692 91652 3720
rect 91005 3683 91063 3689
rect 91646 3680 91652 3692
rect 91704 3680 91710 3732
rect 94961 3723 95019 3729
rect 94961 3689 94973 3723
rect 95007 3720 95019 3723
rect 101674 3720 101680 3732
rect 95007 3692 101680 3720
rect 95007 3689 95019 3692
rect 94961 3683 95019 3689
rect 101674 3680 101680 3692
rect 101732 3680 101738 3732
rect 101766 3680 101772 3732
rect 101824 3720 101830 3732
rect 104253 3723 104311 3729
rect 104253 3720 104265 3723
rect 101824 3692 104265 3720
rect 101824 3680 101830 3692
rect 104253 3689 104265 3692
rect 104299 3689 104311 3723
rect 104253 3683 104311 3689
rect 105357 3723 105415 3729
rect 105357 3689 105369 3723
rect 105403 3689 105415 3723
rect 105357 3683 105415 3689
rect 107565 3723 107623 3729
rect 107565 3689 107577 3723
rect 107611 3689 107623 3723
rect 109310 3720 109316 3732
rect 109271 3692 109316 3720
rect 107565 3683 107623 3689
rect 85206 3612 85212 3664
rect 85264 3652 85270 3664
rect 86862 3652 86868 3664
rect 85264 3624 86868 3652
rect 85264 3612 85270 3624
rect 86862 3612 86868 3624
rect 86920 3612 86926 3664
rect 87049 3655 87107 3661
rect 87049 3652 87061 3655
rect 86972 3624 87061 3652
rect 84473 3587 84531 3593
rect 84473 3553 84485 3587
rect 84519 3584 84531 3587
rect 84841 3587 84899 3593
rect 84519 3556 84792 3584
rect 84519 3553 84531 3556
rect 84473 3547 84531 3553
rect 81952 3488 83136 3516
rect 83185 3519 83243 3525
rect 81952 3476 81958 3488
rect 83185 3485 83197 3519
rect 83231 3516 83243 3519
rect 83277 3519 83335 3525
rect 83277 3516 83289 3519
rect 83231 3488 83289 3516
rect 83231 3485 83243 3488
rect 83185 3479 83243 3485
rect 83277 3485 83289 3488
rect 83323 3516 83335 3519
rect 83550 3516 83556 3528
rect 83323 3488 83556 3516
rect 83323 3485 83335 3488
rect 83277 3479 83335 3485
rect 83550 3476 83556 3488
rect 83608 3516 83614 3528
rect 84565 3519 84623 3525
rect 84565 3516 84577 3519
rect 83608 3488 84577 3516
rect 83608 3476 83614 3488
rect 84565 3485 84577 3488
rect 84611 3516 84623 3519
rect 84654 3516 84660 3528
rect 84611 3488 84660 3516
rect 84611 3485 84623 3488
rect 84565 3479 84623 3485
rect 84654 3476 84660 3488
rect 84712 3476 84718 3528
rect 84764 3516 84792 3556
rect 84841 3553 84853 3587
rect 84887 3553 84899 3587
rect 85482 3584 85488 3596
rect 85443 3556 85488 3584
rect 84841 3547 84899 3553
rect 85482 3544 85488 3556
rect 85540 3544 85546 3596
rect 85666 3584 85672 3596
rect 85627 3556 85672 3584
rect 85666 3544 85672 3556
rect 85724 3544 85730 3596
rect 86037 3587 86095 3593
rect 86037 3553 86049 3587
rect 86083 3584 86095 3587
rect 86494 3584 86500 3596
rect 86083 3556 86500 3584
rect 86083 3553 86095 3556
rect 86037 3547 86095 3553
rect 86494 3544 86500 3556
rect 86552 3544 86558 3596
rect 85390 3516 85396 3528
rect 84764 3488 85396 3516
rect 85390 3476 85396 3488
rect 85448 3476 85454 3528
rect 85761 3519 85819 3525
rect 85761 3485 85773 3519
rect 85807 3516 85819 3519
rect 85853 3519 85911 3525
rect 85853 3516 85865 3519
rect 85807 3488 85865 3516
rect 85807 3485 85819 3488
rect 85761 3479 85819 3485
rect 85853 3485 85865 3488
rect 85899 3485 85911 3519
rect 86972 3516 87000 3624
rect 87049 3621 87061 3624
rect 87095 3621 87107 3655
rect 89530 3652 89536 3664
rect 89491 3624 89536 3652
rect 87049 3615 87107 3621
rect 89530 3612 89536 3624
rect 89588 3612 89594 3664
rect 89714 3612 89720 3664
rect 89772 3652 89778 3664
rect 93946 3652 93952 3664
rect 89772 3624 90864 3652
rect 93907 3624 93952 3652
rect 89772 3612 89778 3624
rect 87322 3544 87328 3596
rect 87380 3584 87386 3596
rect 89162 3584 89168 3596
rect 87380 3556 89168 3584
rect 87380 3544 87386 3556
rect 89162 3544 89168 3556
rect 89220 3544 89226 3596
rect 90174 3584 90180 3596
rect 90135 3556 90180 3584
rect 90174 3544 90180 3556
rect 90232 3544 90238 3596
rect 90836 3593 90864 3624
rect 93946 3612 93952 3624
rect 94004 3612 94010 3664
rect 95602 3612 95608 3664
rect 95660 3652 95666 3664
rect 101398 3652 101404 3664
rect 95660 3624 101404 3652
rect 95660 3612 95666 3624
rect 101398 3612 101404 3624
rect 101456 3612 101462 3664
rect 101858 3612 101864 3664
rect 101916 3652 101922 3664
rect 105372 3652 105400 3683
rect 101916 3624 105400 3652
rect 101916 3612 101922 3624
rect 90821 3587 90879 3593
rect 90821 3553 90833 3587
rect 90867 3553 90879 3587
rect 90821 3547 90879 3553
rect 90910 3544 90916 3596
rect 90968 3584 90974 3596
rect 91465 3587 91523 3593
rect 91465 3584 91477 3587
rect 90968 3556 91477 3584
rect 90968 3544 90974 3556
rect 91465 3553 91477 3556
rect 91511 3553 91523 3587
rect 91465 3547 91523 3553
rect 91922 3544 91928 3596
rect 91980 3584 91986 3596
rect 92109 3587 92167 3593
rect 92109 3584 92121 3587
rect 91980 3556 92121 3584
rect 91980 3544 91986 3556
rect 92109 3553 92121 3556
rect 92155 3553 92167 3587
rect 92109 3547 92167 3553
rect 94682 3544 94688 3596
rect 94740 3544 94746 3596
rect 95510 3544 95516 3596
rect 95568 3584 95574 3596
rect 96157 3587 96215 3593
rect 96157 3584 96169 3587
rect 95568 3556 96169 3584
rect 95568 3544 95574 3556
rect 96157 3553 96169 3556
rect 96203 3553 96215 3587
rect 96157 3547 96215 3553
rect 96246 3544 96252 3596
rect 96304 3584 96310 3596
rect 96801 3587 96859 3593
rect 96801 3584 96813 3587
rect 96304 3556 96813 3584
rect 96304 3544 96310 3556
rect 96801 3553 96813 3556
rect 96847 3553 96859 3587
rect 97442 3584 97448 3596
rect 97403 3556 97448 3584
rect 96801 3547 96859 3553
rect 97442 3544 97448 3556
rect 97500 3544 97506 3596
rect 98546 3544 98552 3596
rect 98604 3584 98610 3596
rect 98641 3587 98699 3593
rect 98641 3584 98653 3587
rect 98604 3556 98653 3584
rect 98604 3544 98610 3556
rect 98641 3553 98653 3556
rect 98687 3553 98699 3587
rect 99650 3584 99656 3596
rect 99611 3556 99656 3584
rect 98641 3547 98699 3553
rect 99650 3544 99656 3556
rect 99708 3544 99714 3596
rect 100297 3587 100355 3593
rect 100297 3553 100309 3587
rect 100343 3584 100355 3587
rect 100754 3584 100760 3596
rect 100343 3556 100760 3584
rect 100343 3553 100355 3556
rect 100297 3547 100355 3553
rect 100754 3544 100760 3556
rect 100812 3544 100818 3596
rect 101950 3544 101956 3596
rect 102008 3584 102014 3596
rect 102689 3587 102747 3593
rect 102689 3584 102701 3587
rect 102008 3556 102701 3584
rect 102008 3544 102014 3556
rect 102689 3553 102701 3556
rect 102735 3553 102747 3587
rect 104066 3584 104072 3596
rect 104027 3556 104072 3584
rect 102689 3547 102747 3553
rect 104066 3544 104072 3556
rect 104124 3544 104130 3596
rect 105170 3584 105176 3596
rect 105131 3556 105176 3584
rect 105170 3544 105176 3556
rect 105228 3544 105234 3596
rect 106274 3584 106280 3596
rect 106235 3556 106280 3584
rect 106274 3544 106280 3556
rect 106332 3544 106338 3596
rect 107378 3584 107384 3596
rect 107339 3556 107384 3584
rect 107378 3544 107384 3556
rect 107436 3544 107442 3596
rect 93302 3516 93308 3528
rect 86972 3488 93308 3516
rect 85853 3479 85911 3485
rect 80664 3420 81388 3448
rect 80664 3408 80670 3420
rect 81434 3408 81440 3460
rect 81492 3408 81498 3460
rect 81526 3408 81532 3460
rect 81584 3448 81590 3460
rect 82538 3448 82544 3460
rect 81584 3420 82544 3448
rect 81584 3408 81590 3420
rect 82538 3408 82544 3420
rect 82596 3408 82602 3460
rect 83645 3451 83703 3457
rect 83645 3417 83657 3451
rect 83691 3448 83703 3451
rect 83691 3420 84056 3448
rect 83691 3417 83703 3420
rect 83645 3411 83703 3417
rect 81066 3380 81072 3392
rect 80532 3352 81072 3380
rect 80425 3343 80483 3349
rect 81066 3340 81072 3352
rect 81124 3340 81130 3392
rect 81158 3340 81164 3392
rect 81216 3380 81222 3392
rect 83734 3380 83740 3392
rect 81216 3352 83740 3380
rect 81216 3340 81222 3352
rect 83734 3340 83740 3352
rect 83792 3340 83798 3392
rect 84028 3380 84056 3420
rect 84286 3408 84292 3460
rect 84344 3448 84350 3460
rect 85868 3448 85896 3479
rect 93302 3476 93308 3488
rect 93360 3476 93366 3528
rect 101398 3516 101404 3528
rect 95726 3488 101404 3516
rect 101398 3476 101404 3488
rect 101456 3476 101462 3528
rect 101582 3476 101588 3528
rect 101640 3516 101646 3528
rect 107580 3516 107608 3683
rect 109310 3680 109316 3692
rect 109368 3680 109374 3732
rect 109954 3720 109960 3732
rect 109915 3692 109960 3720
rect 109954 3680 109960 3692
rect 110012 3680 110018 3732
rect 108482 3544 108488 3596
rect 108540 3584 108546 3596
rect 109129 3587 109187 3593
rect 109129 3584 109141 3587
rect 108540 3556 109141 3584
rect 108540 3544 108546 3556
rect 109129 3553 109141 3556
rect 109175 3553 109187 3587
rect 109129 3547 109187 3553
rect 109218 3544 109224 3596
rect 109276 3584 109282 3596
rect 109773 3587 109831 3593
rect 109773 3584 109785 3587
rect 109276 3556 109785 3584
rect 109276 3544 109282 3556
rect 109773 3553 109785 3556
rect 109819 3553 109831 3587
rect 110690 3584 110696 3596
rect 110651 3556 110696 3584
rect 109773 3547 109831 3553
rect 110690 3544 110696 3556
rect 110748 3544 110754 3596
rect 111797 3587 111855 3593
rect 111797 3553 111809 3587
rect 111843 3584 111855 3587
rect 112070 3584 112076 3596
rect 111843 3556 112076 3584
rect 111843 3553 111855 3556
rect 111797 3547 111855 3553
rect 112070 3544 112076 3556
rect 112128 3544 112134 3596
rect 112898 3584 112904 3596
rect 112859 3556 112904 3584
rect 112898 3544 112904 3556
rect 112956 3544 112962 3596
rect 114002 3544 114008 3596
rect 114060 3584 114066 3596
rect 114373 3587 114431 3593
rect 114373 3584 114385 3587
rect 114060 3556 114385 3584
rect 114060 3544 114066 3556
rect 114373 3553 114385 3556
rect 114419 3553 114431 3587
rect 115106 3584 115112 3596
rect 115067 3556 115112 3584
rect 114373 3547 114431 3553
rect 115106 3544 115112 3556
rect 115164 3544 115170 3596
rect 116210 3584 116216 3596
rect 116171 3556 116216 3584
rect 116210 3544 116216 3556
rect 116268 3544 116274 3596
rect 117314 3584 117320 3596
rect 117275 3556 117320 3584
rect 117314 3544 117320 3556
rect 117372 3544 117378 3596
rect 118418 3584 118424 3596
rect 118379 3556 118424 3584
rect 118418 3544 118424 3556
rect 118476 3544 118482 3596
rect 119522 3544 119528 3596
rect 119580 3584 119586 3596
rect 119617 3587 119675 3593
rect 119617 3584 119629 3587
rect 119580 3556 119629 3584
rect 119580 3544 119586 3556
rect 119617 3553 119629 3556
rect 119663 3553 119675 3587
rect 120534 3584 120540 3596
rect 120495 3556 120540 3584
rect 119617 3547 119675 3553
rect 120534 3544 120540 3556
rect 120592 3544 120598 3596
rect 121638 3584 121644 3596
rect 121599 3556 121644 3584
rect 121638 3544 121644 3556
rect 121696 3544 121702 3596
rect 122742 3584 122748 3596
rect 122703 3556 122748 3584
rect 122742 3544 122748 3556
rect 122800 3544 122806 3596
rect 123757 3587 123815 3593
rect 123757 3553 123769 3587
rect 123803 3584 123815 3587
rect 123846 3584 123852 3596
rect 123803 3556 123852 3584
rect 123803 3553 123815 3556
rect 123757 3547 123815 3553
rect 123846 3544 123852 3556
rect 123904 3544 123910 3596
rect 124950 3584 124956 3596
rect 124911 3556 124956 3584
rect 124950 3544 124956 3556
rect 125008 3544 125014 3596
rect 126054 3584 126060 3596
rect 126015 3556 126060 3584
rect 126054 3544 126060 3556
rect 126112 3544 126118 3596
rect 126974 3544 126980 3596
rect 127032 3584 127038 3596
rect 127161 3587 127219 3593
rect 127161 3584 127173 3587
rect 127032 3556 127173 3584
rect 127032 3544 127038 3556
rect 127161 3553 127173 3556
rect 127207 3553 127219 3587
rect 128262 3584 128268 3596
rect 128223 3556 128268 3584
rect 127161 3547 127219 3553
rect 128262 3544 128268 3556
rect 128320 3544 128326 3596
rect 128998 3584 129004 3596
rect 128959 3556 129004 3584
rect 128998 3544 129004 3556
rect 129056 3544 129062 3596
rect 129366 3544 129372 3596
rect 129424 3584 129430 3596
rect 130105 3587 130163 3593
rect 130105 3584 130117 3587
rect 129424 3556 130117 3584
rect 129424 3544 129430 3556
rect 130105 3553 130117 3556
rect 130151 3553 130163 3587
rect 130105 3547 130163 3553
rect 130194 3544 130200 3596
rect 130252 3584 130258 3596
rect 130749 3587 130807 3593
rect 130749 3584 130761 3587
rect 130252 3556 130761 3584
rect 130252 3544 130258 3556
rect 130749 3553 130761 3556
rect 130795 3553 130807 3587
rect 130749 3547 130807 3553
rect 131574 3544 131580 3596
rect 131632 3584 131638 3596
rect 132405 3587 132463 3593
rect 132405 3584 132417 3587
rect 131632 3556 132417 3584
rect 131632 3544 131638 3556
rect 132405 3553 132417 3556
rect 132451 3553 132463 3587
rect 132405 3547 132463 3553
rect 133049 3587 133107 3593
rect 133049 3553 133061 3587
rect 133095 3553 133107 3587
rect 133782 3584 133788 3596
rect 133743 3556 133788 3584
rect 133049 3547 133107 3553
rect 101640 3488 107608 3516
rect 101640 3476 101646 3488
rect 132310 3476 132316 3528
rect 132368 3516 132374 3528
rect 133064 3516 133092 3547
rect 133782 3544 133788 3556
rect 133840 3544 133846 3596
rect 134886 3544 134892 3596
rect 134944 3584 134950 3596
rect 135349 3587 135407 3593
rect 135349 3584 135361 3587
rect 134944 3556 135361 3584
rect 134944 3544 134950 3556
rect 135349 3553 135361 3556
rect 135395 3553 135407 3587
rect 135349 3547 135407 3553
rect 135622 3544 135628 3596
rect 135680 3584 135686 3596
rect 135993 3587 136051 3593
rect 135993 3584 136005 3587
rect 135680 3556 136005 3584
rect 135680 3544 135686 3556
rect 135993 3553 136005 3556
rect 136039 3553 136051 3587
rect 137094 3584 137100 3596
rect 137055 3556 137100 3584
rect 135993 3547 136051 3553
rect 137094 3544 137100 3556
rect 137152 3544 137158 3596
rect 138198 3584 138204 3596
rect 138159 3556 138204 3584
rect 138198 3544 138204 3556
rect 138256 3544 138262 3596
rect 139302 3584 139308 3596
rect 139263 3556 139308 3584
rect 139302 3544 139308 3556
rect 139360 3544 139366 3596
rect 140406 3544 140412 3596
rect 140464 3584 140470 3596
rect 140593 3587 140651 3593
rect 140593 3584 140605 3587
rect 140464 3556 140605 3584
rect 140464 3544 140470 3556
rect 140593 3553 140605 3556
rect 140639 3553 140651 3587
rect 141510 3584 141516 3596
rect 141471 3556 141516 3584
rect 140593 3547 140651 3553
rect 141510 3544 141516 3556
rect 141568 3544 141574 3596
rect 142617 3587 142675 3593
rect 142617 3553 142629 3587
rect 142663 3584 142675 3587
rect 142798 3584 142804 3596
rect 142663 3556 142804 3584
rect 142663 3553 142675 3556
rect 142617 3547 142675 3553
rect 142798 3544 142804 3556
rect 142856 3544 142862 3596
rect 143718 3584 143724 3596
rect 143679 3556 143724 3584
rect 143718 3544 143724 3556
rect 143776 3544 143782 3596
rect 144733 3587 144791 3593
rect 144733 3553 144745 3587
rect 144779 3584 144791 3587
rect 144822 3584 144828 3596
rect 144779 3556 144828 3584
rect 144779 3553 144791 3556
rect 144733 3547 144791 3553
rect 144822 3544 144828 3556
rect 144880 3544 144886 3596
rect 145926 3584 145932 3596
rect 145887 3556 145932 3584
rect 145926 3544 145932 3556
rect 145984 3544 145990 3596
rect 147030 3584 147036 3596
rect 146991 3556 147036 3584
rect 147030 3544 147036 3556
rect 147088 3544 147094 3596
rect 148134 3584 148140 3596
rect 148095 3556 148140 3584
rect 148134 3544 148140 3556
rect 148192 3544 148198 3596
rect 149238 3584 149244 3596
rect 149199 3556 149244 3584
rect 149238 3544 149244 3556
rect 149296 3544 149302 3596
rect 149974 3584 149980 3596
rect 149935 3556 149980 3584
rect 149974 3544 149980 3556
rect 150032 3544 150038 3596
rect 150342 3544 150348 3596
rect 150400 3584 150406 3596
rect 151081 3587 151139 3593
rect 151081 3584 151093 3587
rect 150400 3556 151093 3584
rect 150400 3544 150406 3556
rect 151081 3553 151093 3556
rect 151127 3553 151139 3587
rect 151081 3547 151139 3553
rect 151170 3544 151176 3596
rect 151228 3584 151234 3596
rect 151725 3587 151783 3593
rect 151725 3584 151737 3587
rect 151228 3556 151737 3584
rect 151228 3544 151234 3556
rect 151725 3553 151737 3556
rect 151771 3553 151783 3587
rect 153654 3584 153660 3596
rect 153615 3556 153660 3584
rect 151725 3547 151783 3553
rect 153654 3544 153660 3556
rect 153712 3544 153718 3596
rect 154758 3584 154764 3596
rect 154719 3556 154764 3584
rect 154758 3544 154764 3556
rect 154816 3544 154822 3596
rect 155862 3544 155868 3596
rect 155920 3584 155926 3596
rect 156325 3587 156383 3593
rect 156325 3584 156337 3587
rect 155920 3556 156337 3584
rect 155920 3544 155926 3556
rect 156325 3553 156337 3556
rect 156371 3553 156383 3587
rect 156325 3547 156383 3553
rect 156598 3544 156604 3596
rect 156656 3584 156662 3596
rect 156969 3587 157027 3593
rect 156969 3584 156981 3587
rect 156656 3556 156981 3584
rect 156656 3544 156662 3556
rect 156969 3553 156981 3556
rect 157015 3553 157027 3587
rect 156969 3547 157027 3553
rect 158073 3587 158131 3593
rect 158073 3553 158085 3587
rect 158119 3584 158131 3587
rect 158162 3584 158168 3596
rect 158119 3556 158168 3584
rect 158119 3553 158131 3556
rect 158073 3547 158131 3553
rect 158162 3544 158168 3556
rect 158220 3544 158226 3596
rect 159174 3584 159180 3596
rect 159135 3556 159180 3584
rect 159174 3544 159180 3556
rect 159232 3544 159238 3596
rect 160278 3584 160284 3596
rect 160239 3556 160284 3584
rect 160278 3544 160284 3556
rect 160336 3544 160342 3596
rect 161382 3544 161388 3596
rect 161440 3584 161446 3596
rect 161569 3587 161627 3593
rect 161569 3584 161581 3587
rect 161440 3556 161581 3584
rect 161440 3544 161446 3556
rect 161569 3553 161581 3556
rect 161615 3553 161627 3587
rect 162486 3584 162492 3596
rect 162447 3556 162492 3584
rect 161569 3547 161627 3553
rect 162486 3544 162492 3556
rect 162544 3544 162550 3596
rect 163590 3584 163596 3596
rect 163551 3556 163596 3584
rect 163590 3544 163596 3556
rect 163648 3544 163654 3596
rect 164237 3587 164295 3593
rect 164237 3553 164249 3587
rect 164283 3553 164295 3587
rect 164237 3547 164295 3553
rect 132368 3488 133092 3516
rect 132368 3476 132374 3488
rect 163222 3476 163228 3528
rect 163280 3516 163286 3528
rect 164252 3516 164280 3547
rect 164418 3544 164424 3596
rect 164476 3584 164482 3596
rect 164881 3587 164939 3593
rect 164881 3584 164893 3587
rect 164476 3556 164893 3584
rect 164476 3544 164482 3556
rect 164881 3553 164893 3556
rect 164927 3553 164939 3587
rect 164881 3547 164939 3553
rect 165709 3587 165767 3593
rect 165709 3553 165721 3587
rect 165755 3584 165767 3587
rect 165798 3584 165804 3596
rect 165755 3556 165804 3584
rect 165755 3553 165767 3556
rect 165709 3547 165767 3553
rect 165798 3544 165804 3556
rect 165856 3544 165862 3596
rect 166902 3584 166908 3596
rect 166863 3556 166908 3584
rect 166902 3544 166908 3556
rect 166960 3544 166966 3596
rect 168006 3584 168012 3596
rect 167967 3556 168012 3584
rect 168006 3544 168012 3556
rect 168064 3544 168070 3596
rect 169110 3584 169116 3596
rect 169071 3556 169116 3584
rect 169110 3544 169116 3556
rect 169168 3544 169174 3596
rect 170214 3584 170220 3596
rect 170175 3556 170220 3584
rect 170214 3544 170220 3556
rect 170272 3544 170278 3596
rect 170950 3584 170956 3596
rect 170911 3556 170956 3584
rect 170950 3544 170956 3556
rect 171008 3544 171014 3596
rect 171318 3544 171324 3596
rect 171376 3584 171382 3596
rect 172057 3587 172115 3593
rect 172057 3584 172069 3587
rect 171376 3556 172069 3584
rect 171376 3544 171382 3556
rect 172057 3553 172069 3556
rect 172103 3553 172115 3587
rect 172057 3547 172115 3553
rect 172146 3544 172152 3596
rect 172204 3584 172210 3596
rect 172701 3587 172759 3593
rect 172701 3584 172713 3587
rect 172204 3556 172713 3584
rect 172204 3544 172210 3556
rect 172701 3553 172713 3556
rect 172747 3553 172759 3587
rect 172701 3547 172759 3553
rect 173526 3544 173532 3596
rect 173584 3584 173590 3596
rect 174357 3587 174415 3593
rect 174357 3584 174369 3587
rect 173584 3556 174369 3584
rect 173584 3544 173590 3556
rect 174357 3553 174369 3556
rect 174403 3553 174415 3587
rect 174357 3547 174415 3553
rect 174630 3544 174636 3596
rect 174688 3584 174694 3596
rect 175001 3587 175059 3593
rect 175001 3584 175013 3587
rect 174688 3556 175013 3584
rect 174688 3544 174694 3556
rect 175001 3553 175013 3556
rect 175047 3553 175059 3587
rect 175001 3547 175059 3553
rect 176381 3587 176439 3593
rect 176381 3553 176393 3587
rect 176427 3584 176439 3587
rect 177945 3587 178003 3593
rect 177945 3584 177957 3587
rect 176427 3556 177957 3584
rect 176427 3553 176439 3556
rect 176381 3547 176439 3553
rect 177945 3553 177957 3556
rect 177991 3553 178003 3587
rect 177945 3547 178003 3553
rect 163280 3488 164280 3516
rect 163280 3476 163286 3488
rect 84344 3420 85896 3448
rect 84344 3408 84350 3420
rect 84562 3380 84568 3392
rect 84028 3352 84568 3380
rect 84562 3340 84568 3352
rect 84620 3340 84626 3392
rect 85868 3380 85896 3420
rect 86681 3451 86739 3457
rect 86681 3417 86693 3451
rect 86727 3448 86739 3451
rect 86770 3448 86776 3460
rect 86727 3420 86776 3448
rect 86727 3417 86739 3420
rect 86681 3411 86739 3417
rect 86770 3408 86776 3420
rect 86828 3408 86834 3460
rect 88058 3408 88064 3460
rect 88116 3448 88122 3460
rect 88153 3451 88211 3457
rect 88153 3448 88165 3451
rect 88116 3420 88165 3448
rect 88116 3408 88122 3420
rect 88153 3417 88165 3420
rect 88199 3417 88211 3451
rect 90361 3451 90419 3457
rect 90361 3448 90373 3451
rect 88153 3411 88211 3417
rect 89364 3420 90373 3448
rect 86586 3380 86592 3392
rect 85868 3352 86592 3380
rect 86586 3340 86592 3352
rect 86644 3340 86650 3392
rect 87046 3380 87052 3392
rect 87007 3352 87052 3380
rect 87046 3340 87052 3352
rect 87104 3380 87110 3392
rect 88518 3380 88524 3392
rect 87104 3352 88524 3380
rect 87104 3340 87110 3352
rect 88518 3340 88524 3352
rect 88576 3340 88582 3392
rect 88705 3383 88763 3389
rect 88705 3349 88717 3383
rect 88751 3380 88763 3383
rect 89070 3380 89076 3392
rect 88751 3352 89076 3380
rect 88751 3349 88763 3352
rect 88705 3343 88763 3349
rect 89070 3340 89076 3352
rect 89128 3340 89134 3392
rect 89162 3340 89168 3392
rect 89220 3380 89226 3392
rect 89364 3380 89392 3420
rect 90361 3417 90373 3420
rect 90407 3417 90419 3451
rect 90361 3411 90419 3417
rect 90818 3408 90824 3460
rect 90876 3448 90882 3460
rect 92293 3451 92351 3457
rect 92293 3448 92305 3451
rect 90876 3420 92305 3448
rect 90876 3408 90882 3420
rect 92293 3417 92305 3420
rect 92339 3417 92351 3451
rect 92293 3411 92351 3417
rect 95142 3408 95148 3460
rect 95200 3448 95206 3460
rect 96985 3451 97043 3457
rect 96985 3448 96997 3451
rect 95200 3420 96997 3448
rect 95200 3408 95206 3420
rect 96985 3417 96997 3420
rect 97031 3417 97043 3451
rect 96985 3411 97043 3417
rect 98086 3408 98092 3460
rect 98144 3448 98150 3460
rect 99837 3451 99895 3457
rect 99837 3448 99849 3451
rect 98144 3420 99849 3448
rect 98144 3408 98150 3420
rect 99837 3417 99849 3420
rect 99883 3417 99895 3451
rect 102042 3448 102048 3460
rect 99837 3411 99895 3417
rect 100312 3420 102048 3448
rect 89220 3352 89392 3380
rect 89533 3383 89591 3389
rect 89220 3340 89226 3352
rect 89533 3349 89545 3383
rect 89579 3380 89591 3383
rect 89622 3380 89628 3392
rect 89579 3352 89628 3380
rect 89579 3349 89591 3352
rect 89533 3343 89591 3349
rect 89622 3340 89628 3352
rect 89680 3340 89686 3392
rect 89717 3383 89775 3389
rect 89717 3349 89729 3383
rect 89763 3380 89775 3383
rect 89806 3380 89812 3392
rect 89763 3352 89812 3380
rect 89763 3349 89775 3352
rect 89717 3343 89775 3349
rect 89806 3340 89812 3352
rect 89864 3340 89870 3392
rect 93486 3340 93492 3392
rect 93544 3380 93550 3392
rect 96341 3383 96399 3389
rect 96341 3380 96353 3383
rect 93544 3352 96353 3380
rect 93544 3340 93550 3352
rect 96341 3349 96353 3352
rect 96387 3349 96399 3383
rect 97626 3380 97632 3392
rect 97587 3352 97632 3380
rect 96341 3343 96399 3349
rect 97626 3340 97632 3352
rect 97684 3340 97690 3392
rect 98822 3380 98828 3392
rect 98783 3352 98828 3380
rect 98822 3340 98828 3352
rect 98880 3340 98886 3392
rect 98914 3340 98920 3392
rect 98972 3380 98978 3392
rect 100312 3380 100340 3420
rect 102042 3408 102048 3420
rect 102100 3408 102106 3460
rect 102318 3408 102324 3460
rect 102376 3448 102382 3460
rect 110877 3451 110935 3457
rect 110877 3448 110889 3451
rect 102376 3420 110889 3448
rect 102376 3408 102382 3420
rect 110877 3417 110889 3420
rect 110923 3417 110935 3451
rect 110877 3411 110935 3417
rect 178129 3451 178187 3457
rect 178129 3417 178141 3451
rect 178175 3448 178187 3451
rect 179414 3448 179420 3460
rect 178175 3420 179420 3448
rect 178175 3417 178187 3420
rect 178129 3411 178187 3417
rect 179414 3408 179420 3420
rect 179472 3408 179478 3460
rect 100478 3380 100484 3392
rect 98972 3352 100340 3380
rect 100439 3352 100484 3380
rect 98972 3340 98978 3352
rect 100478 3340 100484 3352
rect 100536 3340 100542 3392
rect 101125 3383 101183 3389
rect 101125 3349 101137 3383
rect 101171 3380 101183 3383
rect 101858 3380 101864 3392
rect 101171 3352 101864 3380
rect 101171 3349 101183 3352
rect 101125 3343 101183 3349
rect 101858 3340 101864 3352
rect 101916 3340 101922 3392
rect 102226 3380 102232 3392
rect 102187 3352 102232 3380
rect 102226 3340 102232 3352
rect 102284 3340 102290 3392
rect 102870 3380 102876 3392
rect 102831 3352 102876 3380
rect 102870 3340 102876 3352
rect 102928 3340 102934 3392
rect 106458 3380 106464 3392
rect 106419 3352 106464 3380
rect 106458 3340 106464 3352
rect 106516 3340 106522 3392
rect 131942 3380 131948 3392
rect 131903 3352 131948 3380
rect 131942 3340 131948 3352
rect 132000 3340 132006 3392
rect 152921 3383 152979 3389
rect 152921 3349 152933 3383
rect 152967 3380 152979 3383
rect 153746 3380 153752 3392
rect 152967 3352 153752 3380
rect 152967 3349 152979 3352
rect 152921 3343 152979 3349
rect 153746 3340 153752 3352
rect 153804 3340 153810 3392
rect 173894 3380 173900 3392
rect 173855 3352 173900 3380
rect 173894 3340 173900 3352
rect 173952 3340 173958 3392
rect 1104 3290 178848 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 34966 3290
rect 35018 3238 35030 3290
rect 35082 3238 35094 3290
rect 35146 3238 35158 3290
rect 35210 3238 65686 3290
rect 65738 3238 65750 3290
rect 65802 3238 65814 3290
rect 65866 3238 65878 3290
rect 65930 3238 96406 3290
rect 96458 3238 96470 3290
rect 96522 3238 96534 3290
rect 96586 3238 96598 3290
rect 96650 3238 127126 3290
rect 127178 3238 127190 3290
rect 127242 3238 127254 3290
rect 127306 3238 127318 3290
rect 127370 3238 157846 3290
rect 157898 3238 157910 3290
rect 157962 3238 157974 3290
rect 158026 3238 158038 3290
rect 158090 3238 178848 3290
rect 1104 3216 178848 3238
rect 2682 3136 2688 3188
rect 2740 3176 2746 3188
rect 2740 3148 12296 3176
rect 2740 3136 2746 3148
rect 9861 3111 9919 3117
rect 9861 3108 9873 3111
rect 3068 3080 9873 3108
rect 1670 3040 1676 3052
rect 1631 3012 1676 3040
rect 1670 3000 1676 3012
rect 1728 3000 1734 3052
rect 382 2932 388 2984
rect 440 2972 446 2984
rect 1397 2975 1455 2981
rect 1397 2972 1409 2975
rect 440 2944 1409 2972
rect 440 2932 446 2944
rect 1397 2941 1409 2944
rect 1443 2941 1455 2975
rect 1397 2935 1455 2941
rect 2222 2932 2228 2984
rect 2280 2972 2286 2984
rect 3068 2981 3096 3080
rect 9861 3077 9873 3080
rect 9907 3077 9919 3111
rect 9861 3071 9919 3077
rect 9950 3068 9956 3120
rect 10008 3108 10014 3120
rect 11882 3108 11888 3120
rect 10008 3080 11888 3108
rect 10008 3068 10014 3080
rect 11882 3068 11888 3080
rect 11940 3068 11946 3120
rect 4540 3012 11744 3040
rect 2317 2975 2375 2981
rect 2317 2972 2329 2975
rect 2280 2944 2329 2972
rect 2280 2932 2286 2944
rect 2317 2941 2329 2944
rect 2363 2941 2375 2975
rect 2317 2935 2375 2941
rect 3053 2975 3111 2981
rect 3053 2941 3065 2975
rect 3099 2941 3111 2975
rect 3694 2972 3700 2984
rect 3655 2944 3700 2972
rect 3053 2935 3111 2941
rect 3694 2932 3700 2944
rect 3752 2932 3758 2984
rect 4540 2981 4568 3012
rect 4525 2975 4583 2981
rect 4525 2941 4537 2975
rect 4571 2941 4583 2975
rect 5166 2972 5172 2984
rect 5127 2944 5172 2972
rect 4525 2935 4583 2941
rect 5166 2932 5172 2944
rect 5224 2932 5230 2984
rect 6638 2932 6644 2984
rect 6696 2972 6702 2984
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 6696 2944 6837 2972
rect 6696 2932 6702 2944
rect 6825 2941 6837 2944
rect 6871 2941 6883 2975
rect 6825 2935 6883 2941
rect 7742 2932 7748 2984
rect 7800 2972 7806 2984
rect 7929 2975 7987 2981
rect 7929 2972 7941 2975
rect 7800 2944 7941 2972
rect 7800 2932 7806 2944
rect 7929 2941 7941 2944
rect 7975 2941 7987 2975
rect 9214 2972 9220 2984
rect 9175 2944 9220 2972
rect 7929 2935 7987 2941
rect 9214 2932 9220 2944
rect 9272 2932 9278 2984
rect 9861 2975 9919 2981
rect 9861 2941 9873 2975
rect 9907 2972 9919 2975
rect 9907 2944 11192 2972
rect 9907 2941 9919 2944
rect 9861 2935 9919 2941
rect 10042 2904 10048 2916
rect 10003 2876 10048 2904
rect 10042 2864 10048 2876
rect 10100 2864 10106 2916
rect 10962 2904 10968 2916
rect 10923 2876 10968 2904
rect 10962 2864 10968 2876
rect 11020 2864 11026 2916
rect 2958 2796 2964 2848
rect 3016 2836 3022 2848
rect 3145 2839 3203 2845
rect 3145 2836 3157 2839
rect 3016 2808 3157 2836
rect 3016 2796 3022 2808
rect 3145 2805 3157 2808
rect 3191 2805 3203 2839
rect 4614 2836 4620 2848
rect 4575 2808 4620 2836
rect 3145 2799 3203 2805
rect 4614 2796 4620 2808
rect 4672 2796 4678 2848
rect 7745 2839 7803 2845
rect 7745 2805 7757 2839
rect 7791 2836 7803 2839
rect 9858 2836 9864 2848
rect 7791 2808 9864 2836
rect 7791 2805 7803 2808
rect 7745 2799 7803 2805
rect 9858 2796 9864 2808
rect 9916 2796 9922 2848
rect 9950 2796 9956 2848
rect 10008 2836 10014 2848
rect 10137 2839 10195 2845
rect 10137 2836 10149 2839
rect 10008 2808 10149 2836
rect 10008 2796 10014 2808
rect 10137 2805 10149 2808
rect 10183 2805 10195 2839
rect 11054 2836 11060 2848
rect 11015 2808 11060 2836
rect 10137 2799 10195 2805
rect 11054 2796 11060 2808
rect 11112 2796 11118 2848
rect 11164 2836 11192 2944
rect 11716 2904 11744 3012
rect 12066 2972 12072 2984
rect 12027 2944 12072 2972
rect 12066 2932 12072 2944
rect 12124 2932 12130 2984
rect 12268 2972 12296 3148
rect 13170 3136 13176 3188
rect 13228 3176 13234 3188
rect 15378 3176 15384 3188
rect 13228 3148 15384 3176
rect 13228 3136 13234 3148
rect 15378 3136 15384 3148
rect 15436 3136 15442 3188
rect 15470 3136 15476 3188
rect 15528 3176 15534 3188
rect 16301 3179 16359 3185
rect 16301 3176 16313 3179
rect 15528 3148 16313 3176
rect 15528 3136 15534 3148
rect 16301 3145 16313 3148
rect 16347 3145 16359 3179
rect 16301 3139 16359 3145
rect 16390 3136 16396 3188
rect 16448 3176 16454 3188
rect 16448 3148 21220 3176
rect 16448 3136 16454 3148
rect 12526 3068 12532 3120
rect 12584 3108 12590 3120
rect 17678 3108 17684 3120
rect 12584 3080 17356 3108
rect 17639 3080 17684 3108
rect 12584 3068 12590 3080
rect 12437 3043 12495 3049
rect 12437 3009 12449 3043
rect 12483 3040 12495 3043
rect 12483 3012 13308 3040
rect 12483 3009 12495 3012
rect 12437 3003 12495 3009
rect 12621 2975 12679 2981
rect 12621 2972 12633 2975
rect 12268 2944 12633 2972
rect 12621 2941 12633 2944
rect 12667 2941 12679 2975
rect 13280 2972 13308 3012
rect 13354 3000 13360 3052
rect 13412 3040 13418 3052
rect 15194 3040 15200 3052
rect 13412 3012 15200 3040
rect 13412 3000 13418 3012
rect 15194 3000 15200 3012
rect 15252 3040 15258 3052
rect 17328 3049 17356 3080
rect 17678 3068 17684 3080
rect 17736 3068 17742 3120
rect 21082 3108 21088 3120
rect 18800 3080 21088 3108
rect 15289 3043 15347 3049
rect 15289 3040 15301 3043
rect 15252 3012 15301 3040
rect 15252 3000 15258 3012
rect 15289 3009 15301 3012
rect 15335 3009 15347 3043
rect 15289 3003 15347 3009
rect 17313 3043 17371 3049
rect 17313 3009 17325 3043
rect 17359 3009 17371 3043
rect 18800 3040 18828 3080
rect 21082 3068 21088 3080
rect 21140 3068 21146 3120
rect 21192 3108 21220 3148
rect 21266 3136 21272 3188
rect 21324 3176 21330 3188
rect 24302 3176 24308 3188
rect 21324 3148 24308 3176
rect 21324 3136 21330 3148
rect 24302 3136 24308 3148
rect 24360 3136 24366 3188
rect 24486 3176 24492 3188
rect 24447 3148 24492 3176
rect 24486 3136 24492 3148
rect 24544 3136 24550 3188
rect 24578 3136 24584 3188
rect 24636 3176 24642 3188
rect 27249 3179 27307 3185
rect 24636 3148 25084 3176
rect 24636 3136 24642 3148
rect 22370 3108 22376 3120
rect 21192 3080 22376 3108
rect 22370 3068 22376 3080
rect 22428 3068 22434 3120
rect 25056 3108 25084 3148
rect 27249 3145 27261 3179
rect 27295 3176 27307 3179
rect 38654 3176 38660 3188
rect 27295 3148 38660 3176
rect 27295 3145 27307 3148
rect 27249 3139 27307 3145
rect 38654 3136 38660 3148
rect 38712 3136 38718 3188
rect 40954 3176 40960 3188
rect 39040 3148 40960 3176
rect 28074 3108 28080 3120
rect 25056 3080 28080 3108
rect 28074 3068 28080 3080
rect 28132 3068 28138 3120
rect 28166 3068 28172 3120
rect 28224 3108 28230 3120
rect 30650 3108 30656 3120
rect 28224 3080 30656 3108
rect 28224 3068 28230 3080
rect 30650 3068 30656 3080
rect 30708 3108 30714 3120
rect 31570 3108 31576 3120
rect 30708 3080 31576 3108
rect 30708 3068 30714 3080
rect 31570 3068 31576 3080
rect 31628 3068 31634 3120
rect 36446 3108 36452 3120
rect 31726 3080 36452 3108
rect 17313 3003 17371 3009
rect 18248 3012 18828 3040
rect 19245 3043 19303 3049
rect 13998 2972 14004 2984
rect 13280 2944 13860 2972
rect 13959 2944 14004 2972
rect 12621 2935 12679 2941
rect 13078 2904 13084 2916
rect 11716 2876 13084 2904
rect 13078 2864 13084 2876
rect 13136 2864 13142 2916
rect 13357 2907 13415 2913
rect 13357 2873 13369 2907
rect 13403 2904 13415 2907
rect 13832 2904 13860 2944
rect 13998 2932 14004 2944
rect 14056 2932 14062 2984
rect 14274 2972 14280 2984
rect 14235 2944 14280 2972
rect 14274 2932 14280 2944
rect 14332 2932 14338 2984
rect 15473 2975 15531 2981
rect 15473 2941 15485 2975
rect 15519 2972 15531 2975
rect 15654 2972 15660 2984
rect 15519 2944 15660 2972
rect 15519 2941 15531 2944
rect 15473 2935 15531 2941
rect 15654 2932 15660 2944
rect 15712 2932 15718 2984
rect 16390 2972 16396 2984
rect 16040 2944 16396 2972
rect 16040 2904 16068 2944
rect 16390 2932 16396 2944
rect 16448 2932 16454 2984
rect 17494 2972 17500 2984
rect 17455 2944 17500 2972
rect 17494 2932 17500 2944
rect 17552 2972 17558 2984
rect 18248 2981 18276 3012
rect 19245 3009 19257 3043
rect 19291 3040 19303 3043
rect 25406 3040 25412 3052
rect 19291 3012 25412 3040
rect 19291 3009 19303 3012
rect 19245 3003 19303 3009
rect 25406 3000 25412 3012
rect 25464 3000 25470 3052
rect 18233 2975 18291 2981
rect 17552 2944 18184 2972
rect 17552 2932 17558 2944
rect 16206 2904 16212 2916
rect 13403 2876 13768 2904
rect 13832 2876 16068 2904
rect 16167 2876 16212 2904
rect 13403 2873 13415 2876
rect 13357 2867 13415 2873
rect 13170 2836 13176 2848
rect 11164 2808 13176 2836
rect 13170 2796 13176 2808
rect 13228 2796 13234 2848
rect 13262 2796 13268 2848
rect 13320 2836 13326 2848
rect 13449 2839 13507 2845
rect 13449 2836 13461 2839
rect 13320 2808 13461 2836
rect 13320 2796 13326 2808
rect 13449 2805 13461 2808
rect 13495 2805 13507 2839
rect 13740 2836 13768 2876
rect 16206 2864 16212 2876
rect 16264 2864 16270 2916
rect 18156 2904 18184 2944
rect 18233 2941 18245 2975
rect 18279 2941 18291 2975
rect 18877 2975 18935 2981
rect 18877 2972 18889 2975
rect 18233 2935 18291 2941
rect 18340 2944 18889 2972
rect 18340 2904 18368 2944
rect 18877 2941 18889 2944
rect 18923 2941 18935 2975
rect 18877 2935 18935 2941
rect 19061 2975 19119 2981
rect 19061 2941 19073 2975
rect 19107 2941 19119 2975
rect 19061 2935 19119 2941
rect 17696 2876 18000 2904
rect 18156 2876 18368 2904
rect 18417 2907 18475 2913
rect 15562 2836 15568 2848
rect 13740 2808 15568 2836
rect 13449 2799 13507 2805
rect 15562 2796 15568 2808
rect 15620 2796 15626 2848
rect 15657 2839 15715 2845
rect 15657 2805 15669 2839
rect 15703 2836 15715 2839
rect 17696 2836 17724 2876
rect 15703 2808 17724 2836
rect 17972 2836 18000 2876
rect 18417 2873 18429 2907
rect 18463 2904 18475 2907
rect 18506 2904 18512 2916
rect 18463 2876 18512 2904
rect 18463 2873 18475 2876
rect 18417 2867 18475 2873
rect 18506 2864 18512 2876
rect 18564 2864 18570 2916
rect 18966 2864 18972 2916
rect 19024 2904 19030 2916
rect 19076 2904 19104 2935
rect 19886 2932 19892 2984
rect 19944 2972 19950 2984
rect 20165 2975 20223 2981
rect 20165 2972 20177 2975
rect 19944 2944 20177 2972
rect 19944 2932 19950 2944
rect 20165 2941 20177 2944
rect 20211 2941 20223 2975
rect 20622 2972 20628 2984
rect 20583 2944 20628 2972
rect 20165 2935 20223 2941
rect 20622 2932 20628 2944
rect 20680 2932 20686 2984
rect 20898 2972 20904 2984
rect 20859 2944 20904 2972
rect 20898 2932 20904 2944
rect 20956 2932 20962 2984
rect 22646 2972 22652 2984
rect 22607 2944 22652 2972
rect 22646 2932 22652 2944
rect 22704 2932 22710 2984
rect 23385 2975 23443 2981
rect 23385 2941 23397 2975
rect 23431 2972 23443 2975
rect 24302 2972 24308 2984
rect 23431 2944 24308 2972
rect 23431 2941 23443 2944
rect 23385 2935 23443 2941
rect 24302 2932 24308 2944
rect 24360 2932 24366 2984
rect 24397 2975 24455 2981
rect 24397 2941 24409 2975
rect 24443 2972 24455 2975
rect 24443 2944 24532 2972
rect 24443 2941 24455 2944
rect 24397 2935 24455 2941
rect 19024 2876 19104 2904
rect 19981 2907 20039 2913
rect 19024 2864 19030 2876
rect 19981 2873 19993 2907
rect 20027 2904 20039 2907
rect 22002 2904 22008 2916
rect 20027 2876 22008 2904
rect 20027 2873 20039 2876
rect 19981 2867 20039 2873
rect 22002 2864 22008 2876
rect 22060 2864 22066 2916
rect 24504 2904 24532 2944
rect 24578 2932 24584 2984
rect 24636 2972 24642 2984
rect 24636 2944 28948 2972
rect 24636 2932 24642 2944
rect 25314 2904 25320 2916
rect 24504 2876 25320 2904
rect 25314 2864 25320 2876
rect 25372 2864 25378 2916
rect 25498 2904 25504 2916
rect 25459 2876 25504 2904
rect 25498 2864 25504 2876
rect 25556 2864 25562 2916
rect 26605 2907 26663 2913
rect 26605 2873 26617 2907
rect 26651 2904 26663 2907
rect 27249 2907 27307 2913
rect 27249 2904 27261 2907
rect 26651 2876 27261 2904
rect 26651 2873 26663 2876
rect 26605 2867 26663 2873
rect 27249 2873 27261 2876
rect 27295 2873 27307 2907
rect 27890 2904 27896 2916
rect 27851 2876 27896 2904
rect 27249 2867 27307 2873
rect 27890 2864 27896 2876
rect 27948 2864 27954 2916
rect 28810 2904 28816 2916
rect 28771 2876 28816 2904
rect 28810 2864 28816 2876
rect 28868 2864 28874 2916
rect 28920 2904 28948 2944
rect 29086 2932 29092 2984
rect 29144 2972 29150 2984
rect 29457 2975 29515 2981
rect 29457 2972 29469 2975
rect 29144 2944 29469 2972
rect 29144 2932 29150 2944
rect 29457 2941 29469 2944
rect 29503 2941 29515 2975
rect 30190 2972 30196 2984
rect 30151 2944 30196 2972
rect 29457 2935 29515 2941
rect 30190 2932 30196 2944
rect 30248 2932 30254 2984
rect 31021 2975 31079 2981
rect 31021 2941 31033 2975
rect 31067 2972 31079 2975
rect 31726 2972 31754 3080
rect 36446 3068 36452 3080
rect 36504 3068 36510 3120
rect 39040 3108 39068 3148
rect 40954 3136 40960 3148
rect 41012 3136 41018 3188
rect 41046 3136 41052 3188
rect 41104 3176 41110 3188
rect 45094 3176 45100 3188
rect 41104 3148 45100 3176
rect 41104 3136 41110 3148
rect 45094 3136 45100 3148
rect 45152 3136 45158 3188
rect 66441 3179 66499 3185
rect 66441 3145 66453 3179
rect 66487 3176 66499 3179
rect 67542 3176 67548 3188
rect 66487 3148 67548 3176
rect 66487 3145 66499 3148
rect 66441 3139 66499 3145
rect 67542 3136 67548 3148
rect 67600 3136 67606 3188
rect 67634 3136 67640 3188
rect 67692 3176 67698 3188
rect 67729 3179 67787 3185
rect 67729 3176 67741 3179
rect 67692 3148 67741 3176
rect 67692 3136 67698 3148
rect 67729 3145 67741 3148
rect 67775 3145 67787 3179
rect 68554 3176 68560 3188
rect 67729 3139 67787 3145
rect 68112 3148 68560 3176
rect 38626 3080 39068 3108
rect 38626 3040 38654 3080
rect 39114 3068 39120 3120
rect 39172 3108 39178 3120
rect 48038 3108 48044 3120
rect 39172 3080 48044 3108
rect 39172 3068 39178 3080
rect 48038 3068 48044 3080
rect 48096 3068 48102 3120
rect 31956 3012 38654 3040
rect 31956 2981 31984 3012
rect 39022 3000 39028 3052
rect 39080 3040 39086 3052
rect 39080 3012 39804 3040
rect 39080 3000 39086 3012
rect 31067 2944 31754 2972
rect 31941 2975 31999 2981
rect 31067 2941 31079 2944
rect 31021 2935 31079 2941
rect 31941 2941 31953 2975
rect 31987 2941 31999 2975
rect 33226 2972 33232 2984
rect 33187 2944 33232 2972
rect 31941 2935 31999 2941
rect 33226 2932 33232 2944
rect 33284 2932 33290 2984
rect 34330 2972 34336 2984
rect 34291 2944 34336 2972
rect 34330 2932 34336 2944
rect 34388 2932 34394 2984
rect 35434 2972 35440 2984
rect 35395 2944 35440 2972
rect 35434 2932 35440 2944
rect 35492 2932 35498 2984
rect 36814 2932 36820 2984
rect 36872 2972 36878 2984
rect 39776 2981 39804 3012
rect 44266 3000 44272 3052
rect 44324 3040 44330 3052
rect 61562 3040 61568 3052
rect 44324 3012 61568 3040
rect 44324 3000 44330 3012
rect 61562 3000 61568 3012
rect 61620 3000 61626 3052
rect 68002 3040 68008 3052
rect 67100 3012 68008 3040
rect 37185 2975 37243 2981
rect 37185 2972 37197 2975
rect 36872 2944 37197 2972
rect 36872 2932 36878 2944
rect 37185 2941 37197 2944
rect 37231 2941 37243 2975
rect 39761 2975 39819 2981
rect 37185 2935 37243 2941
rect 38304 2944 39252 2972
rect 36262 2904 36268 2916
rect 28920 2876 36268 2904
rect 36262 2864 36268 2876
rect 36320 2864 36326 2916
rect 36541 2907 36599 2913
rect 36541 2873 36553 2907
rect 36587 2904 36599 2907
rect 38304 2904 38332 2944
rect 36587 2876 38332 2904
rect 36587 2873 36599 2876
rect 36541 2867 36599 2873
rect 38378 2864 38384 2916
rect 38436 2904 38442 2916
rect 39114 2904 39120 2916
rect 38436 2876 38481 2904
rect 39075 2876 39120 2904
rect 38436 2864 38442 2876
rect 39114 2864 39120 2876
rect 39172 2864 39178 2916
rect 39224 2904 39252 2944
rect 39761 2941 39773 2975
rect 39807 2941 39819 2975
rect 39761 2935 39819 2941
rect 40126 2932 40132 2984
rect 40184 2972 40190 2984
rect 40405 2975 40463 2981
rect 40405 2972 40417 2975
rect 40184 2944 40417 2972
rect 40184 2932 40190 2944
rect 40405 2941 40417 2944
rect 40451 2941 40463 2975
rect 41230 2972 41236 2984
rect 41191 2944 41236 2972
rect 40405 2935 40463 2941
rect 41230 2932 41236 2944
rect 41288 2932 41294 2984
rect 42334 2972 42340 2984
rect 42295 2944 42340 2972
rect 42334 2932 42340 2944
rect 42392 2932 42398 2984
rect 43438 2932 43444 2984
rect 43496 2972 43502 2984
rect 43533 2975 43591 2981
rect 43533 2972 43545 2975
rect 43496 2944 43545 2972
rect 43496 2932 43502 2944
rect 43533 2941 43545 2944
rect 43579 2941 43591 2975
rect 44542 2972 44548 2984
rect 44503 2944 44548 2972
rect 43533 2935 43591 2941
rect 44542 2932 44548 2944
rect 44600 2932 44606 2984
rect 45646 2972 45652 2984
rect 45607 2944 45652 2972
rect 45646 2932 45652 2944
rect 45704 2932 45710 2984
rect 46750 2972 46756 2984
rect 46711 2944 46756 2972
rect 46750 2932 46756 2944
rect 46808 2932 46814 2984
rect 47673 2975 47731 2981
rect 47673 2941 47685 2975
rect 47719 2972 47731 2975
rect 47854 2972 47860 2984
rect 47719 2944 47860 2972
rect 47719 2941 47731 2944
rect 47673 2935 47731 2941
rect 47854 2932 47860 2944
rect 47912 2932 47918 2984
rect 48958 2972 48964 2984
rect 48919 2944 48964 2972
rect 48958 2932 48964 2944
rect 49016 2932 49022 2984
rect 50062 2972 50068 2984
rect 50023 2944 50068 2972
rect 50062 2932 50068 2944
rect 50120 2932 50126 2984
rect 50798 2972 50804 2984
rect 50759 2944 50804 2972
rect 50798 2932 50804 2944
rect 50856 2932 50862 2984
rect 51629 2975 51687 2981
rect 51629 2941 51641 2975
rect 51675 2972 51687 2975
rect 51902 2972 51908 2984
rect 51675 2944 51908 2972
rect 51675 2941 51687 2944
rect 51629 2935 51687 2941
rect 51902 2932 51908 2944
rect 51960 2932 51966 2984
rect 52270 2972 52276 2984
rect 52231 2944 52276 2972
rect 52270 2932 52276 2944
rect 52328 2932 52334 2984
rect 52917 2975 52975 2981
rect 52917 2941 52929 2975
rect 52963 2972 52975 2975
rect 53006 2972 53012 2984
rect 52963 2944 53012 2972
rect 52963 2941 52975 2944
rect 52917 2935 52975 2941
rect 53006 2932 53012 2944
rect 53064 2932 53070 2984
rect 53374 2932 53380 2984
rect 53432 2972 53438 2984
rect 54021 2975 54079 2981
rect 54021 2972 54033 2975
rect 53432 2944 54033 2972
rect 53432 2932 53438 2944
rect 54021 2941 54033 2944
rect 54067 2941 54079 2975
rect 54021 2935 54079 2941
rect 54478 2932 54484 2984
rect 54536 2972 54542 2984
rect 54665 2975 54723 2981
rect 54665 2972 54677 2975
rect 54536 2944 54677 2972
rect 54536 2932 54542 2944
rect 54665 2941 54677 2944
rect 54711 2941 54723 2975
rect 55582 2972 55588 2984
rect 55543 2944 55588 2972
rect 54665 2935 54723 2941
rect 55582 2932 55588 2944
rect 55640 2932 55646 2984
rect 56686 2972 56692 2984
rect 56647 2944 56692 2972
rect 56686 2932 56692 2944
rect 56744 2932 56750 2984
rect 57790 2972 57796 2984
rect 57751 2944 57796 2972
rect 57790 2932 57796 2944
rect 57848 2932 57854 2984
rect 58894 2932 58900 2984
rect 58952 2972 58958 2984
rect 59265 2975 59323 2981
rect 59265 2972 59277 2975
rect 58952 2944 59277 2972
rect 58952 2932 58958 2944
rect 59265 2941 59277 2944
rect 59311 2941 59323 2975
rect 59998 2972 60004 2984
rect 59959 2944 60004 2972
rect 59265 2935 59323 2941
rect 59998 2932 60004 2944
rect 60056 2932 60062 2984
rect 61010 2972 61016 2984
rect 60971 2944 61016 2972
rect 61010 2932 61016 2944
rect 61068 2932 61074 2984
rect 62114 2972 62120 2984
rect 62075 2944 62120 2972
rect 62114 2932 62120 2944
rect 62172 2932 62178 2984
rect 63218 2972 63224 2984
rect 63179 2944 63224 2972
rect 63218 2932 63224 2944
rect 63276 2932 63282 2984
rect 64322 2932 64328 2984
rect 64380 2972 64386 2984
rect 64509 2975 64567 2981
rect 64509 2972 64521 2975
rect 64380 2944 64521 2972
rect 64380 2932 64386 2944
rect 64509 2941 64521 2944
rect 64555 2941 64567 2975
rect 65426 2972 65432 2984
rect 65387 2944 65432 2972
rect 64509 2935 64567 2941
rect 65426 2932 65432 2944
rect 65484 2932 65490 2984
rect 66622 2932 66628 2984
rect 66680 2972 66686 2984
rect 66717 2975 66775 2981
rect 66717 2972 66729 2975
rect 66680 2944 66729 2972
rect 66680 2932 66686 2944
rect 66717 2941 66729 2944
rect 66763 2941 66775 2975
rect 66717 2935 66775 2941
rect 48314 2904 48320 2916
rect 39224 2876 48320 2904
rect 48314 2864 48320 2876
rect 48372 2864 48378 2916
rect 66073 2907 66131 2913
rect 66073 2873 66085 2907
rect 66119 2873 66131 2907
rect 66073 2867 66131 2873
rect 66487 2907 66545 2913
rect 66487 2873 66499 2907
rect 66533 2904 66545 2907
rect 67100 2904 67128 3012
rect 68002 3000 68008 3012
rect 68060 3000 68066 3052
rect 67177 2975 67235 2981
rect 67177 2941 67189 2975
rect 67223 2972 67235 2975
rect 68112 2972 68140 3148
rect 68554 3136 68560 3148
rect 68612 3136 68618 3188
rect 68649 3179 68707 3185
rect 68649 3145 68661 3179
rect 68695 3176 68707 3179
rect 69934 3176 69940 3188
rect 68695 3148 69940 3176
rect 68695 3145 68707 3148
rect 68649 3139 68707 3145
rect 69934 3136 69940 3148
rect 69992 3136 69998 3188
rect 70121 3179 70179 3185
rect 70121 3145 70133 3179
rect 70167 3176 70179 3179
rect 71225 3179 71283 3185
rect 71225 3176 71237 3179
rect 70167 3148 71237 3176
rect 70167 3145 70179 3148
rect 70121 3139 70179 3145
rect 71225 3145 71237 3148
rect 71271 3176 71283 3179
rect 71866 3176 71872 3188
rect 71271 3148 71872 3176
rect 71271 3145 71283 3148
rect 71225 3139 71283 3145
rect 71866 3136 71872 3148
rect 71924 3176 71930 3188
rect 72326 3176 72332 3188
rect 71924 3148 72332 3176
rect 71924 3136 71930 3148
rect 72326 3136 72332 3148
rect 72384 3136 72390 3188
rect 72510 3176 72516 3188
rect 72471 3148 72516 3176
rect 72510 3136 72516 3148
rect 72568 3136 72574 3188
rect 72602 3136 72608 3188
rect 72660 3176 72666 3188
rect 74534 3176 74540 3188
rect 72660 3148 74540 3176
rect 72660 3136 72666 3148
rect 74534 3136 74540 3148
rect 74592 3136 74598 3188
rect 75086 3136 75092 3188
rect 75144 3176 75150 3188
rect 75365 3179 75423 3185
rect 75365 3176 75377 3179
rect 75144 3148 75377 3176
rect 75144 3136 75150 3148
rect 75365 3145 75377 3148
rect 75411 3176 75423 3179
rect 76282 3176 76288 3188
rect 75411 3148 76288 3176
rect 75411 3145 75423 3148
rect 75365 3139 75423 3145
rect 76282 3136 76288 3148
rect 76340 3176 76346 3188
rect 76377 3179 76435 3185
rect 76377 3176 76389 3179
rect 76340 3148 76389 3176
rect 76340 3136 76346 3148
rect 76377 3145 76389 3148
rect 76423 3145 76435 3179
rect 76558 3176 76564 3188
rect 76519 3148 76564 3176
rect 76377 3139 76435 3145
rect 76558 3136 76564 3148
rect 76616 3136 76622 3188
rect 77846 3136 77852 3188
rect 77904 3176 77910 3188
rect 78033 3179 78091 3185
rect 78033 3176 78045 3179
rect 77904 3148 78045 3176
rect 77904 3136 77910 3148
rect 78033 3145 78045 3148
rect 78079 3145 78091 3179
rect 78033 3139 78091 3145
rect 78122 3136 78128 3188
rect 78180 3176 78186 3188
rect 78217 3179 78275 3185
rect 78217 3176 78229 3179
rect 78180 3148 78229 3176
rect 78180 3136 78186 3148
rect 78217 3145 78229 3148
rect 78263 3145 78275 3179
rect 78217 3139 78275 3145
rect 79045 3179 79103 3185
rect 79045 3145 79057 3179
rect 79091 3176 79103 3179
rect 79318 3176 79324 3188
rect 79091 3148 79324 3176
rect 79091 3145 79103 3148
rect 79045 3139 79103 3145
rect 79318 3136 79324 3148
rect 79376 3136 79382 3188
rect 81158 3176 81164 3188
rect 80532 3148 81164 3176
rect 70026 3108 70032 3120
rect 67223 2944 68140 2972
rect 68204 3080 70032 3108
rect 67223 2941 67235 2944
rect 67177 2935 67235 2941
rect 66533 2876 67128 2904
rect 67591 2907 67649 2913
rect 66533 2873 66545 2876
rect 66487 2867 66545 2873
rect 67591 2873 67603 2907
rect 67637 2904 67649 2907
rect 68204 2904 68232 3080
rect 70026 3068 70032 3080
rect 70084 3068 70090 3120
rect 70302 3108 70308 3120
rect 70263 3080 70308 3108
rect 70302 3068 70308 3080
rect 70360 3068 70366 3120
rect 70394 3068 70400 3120
rect 70452 3108 70458 3120
rect 75914 3108 75920 3120
rect 70452 3080 75920 3108
rect 70452 3068 70458 3080
rect 75914 3068 75920 3080
rect 75972 3068 75978 3120
rect 76009 3111 76067 3117
rect 76009 3077 76021 3111
rect 76055 3108 76067 3111
rect 76742 3108 76748 3120
rect 76055 3080 76748 3108
rect 76055 3077 76067 3080
rect 76009 3071 76067 3077
rect 76742 3068 76748 3080
rect 76800 3068 76806 3120
rect 78677 3111 78735 3117
rect 78677 3077 78689 3111
rect 78723 3108 78735 3111
rect 80532 3108 80560 3148
rect 81158 3136 81164 3148
rect 81216 3136 81222 3188
rect 81253 3179 81311 3185
rect 81253 3145 81265 3179
rect 81299 3176 81311 3179
rect 81802 3176 81808 3188
rect 81299 3148 81808 3176
rect 81299 3145 81311 3148
rect 81253 3139 81311 3145
rect 81802 3136 81808 3148
rect 81860 3136 81866 3188
rect 83001 3179 83059 3185
rect 83001 3145 83013 3179
rect 83047 3176 83059 3179
rect 83274 3176 83280 3188
rect 83047 3148 83280 3176
rect 83047 3145 83059 3148
rect 83001 3139 83059 3145
rect 83274 3136 83280 3148
rect 83332 3136 83338 3188
rect 83918 3136 83924 3188
rect 83976 3176 83982 3188
rect 84289 3179 84347 3185
rect 84289 3176 84301 3179
rect 83976 3148 84301 3176
rect 83976 3136 83982 3148
rect 84289 3145 84301 3148
rect 84335 3145 84347 3179
rect 85758 3176 85764 3188
rect 84289 3139 84347 3145
rect 84764 3148 85764 3176
rect 80698 3108 80704 3120
rect 78723 3080 80560 3108
rect 80659 3080 80704 3108
rect 78723 3077 78735 3080
rect 78677 3071 78735 3077
rect 80698 3068 80704 3080
rect 80756 3068 80762 3120
rect 80882 3068 80888 3120
rect 80940 3108 80946 3120
rect 81526 3108 81532 3120
rect 80940 3080 81532 3108
rect 80940 3068 80946 3080
rect 81526 3068 81532 3080
rect 81584 3108 81590 3120
rect 81713 3111 81771 3117
rect 81713 3108 81725 3111
rect 81584 3080 81725 3108
rect 81584 3068 81590 3080
rect 81713 3077 81725 3080
rect 81759 3108 81771 3111
rect 82722 3108 82728 3120
rect 81759 3080 82728 3108
rect 81759 3077 81771 3080
rect 81713 3071 81771 3077
rect 82722 3068 82728 3080
rect 82780 3068 82786 3120
rect 83734 3068 83740 3120
rect 83792 3108 83798 3120
rect 84764 3108 84792 3148
rect 85758 3136 85764 3148
rect 85816 3136 85822 3188
rect 86328 3148 86549 3176
rect 83792 3080 84792 3108
rect 83792 3068 83798 3080
rect 84838 3068 84844 3120
rect 84896 3108 84902 3120
rect 86328 3108 86356 3148
rect 84896 3080 86356 3108
rect 86521 3108 86549 3148
rect 87690 3136 87696 3188
rect 87748 3176 87754 3188
rect 87877 3179 87935 3185
rect 87877 3176 87889 3179
rect 87748 3148 87889 3176
rect 87748 3136 87754 3148
rect 87877 3145 87889 3148
rect 87923 3145 87935 3179
rect 87877 3139 87935 3145
rect 88518 3136 88524 3188
rect 88576 3176 88582 3188
rect 88797 3179 88855 3185
rect 88797 3176 88809 3179
rect 88576 3148 88809 3176
rect 88576 3136 88582 3148
rect 88797 3145 88809 3148
rect 88843 3145 88855 3179
rect 98914 3176 98920 3188
rect 88797 3139 88855 3145
rect 88904 3148 98920 3176
rect 86957 3111 87015 3117
rect 86957 3108 86969 3111
rect 86521 3080 86969 3108
rect 84896 3068 84902 3080
rect 86957 3077 86969 3080
rect 87003 3077 87015 3111
rect 86957 3071 87015 3077
rect 87230 3068 87236 3120
rect 87288 3108 87294 3120
rect 88904 3108 88932 3148
rect 98914 3136 98920 3148
rect 98972 3136 98978 3188
rect 100478 3176 100484 3188
rect 99024 3148 100484 3176
rect 87288 3080 88932 3108
rect 90913 3111 90971 3117
rect 87288 3068 87294 3080
rect 68281 3043 68339 3049
rect 68281 3009 68293 3043
rect 68327 3040 68339 3043
rect 70762 3040 70768 3052
rect 68327 3012 70768 3040
rect 68327 3009 68339 3012
rect 68281 3003 68339 3009
rect 70762 3000 70768 3012
rect 70820 3000 70826 3052
rect 74902 3040 74908 3052
rect 70872 3012 74908 3040
rect 70872 2981 70900 3012
rect 74902 3000 74908 3012
rect 74960 3000 74966 3052
rect 74997 3043 75055 3049
rect 74997 3009 75009 3043
rect 75043 3040 75055 3043
rect 78858 3040 78864 3052
rect 75043 3012 78864 3040
rect 75043 3009 75055 3012
rect 74997 3003 75055 3009
rect 78858 3000 78864 3012
rect 78916 3000 78922 3052
rect 82078 3040 82084 3052
rect 79152 3012 82084 3040
rect 69753 2975 69811 2981
rect 67637 2876 68232 2904
rect 68572 2944 68968 2972
rect 67637 2873 67649 2876
rect 67591 2867 67649 2873
rect 21266 2836 21272 2848
rect 17972 2808 21272 2836
rect 15703 2805 15715 2808
rect 15657 2799 15715 2805
rect 21266 2796 21272 2808
rect 21324 2796 21330 2848
rect 22094 2796 22100 2848
rect 22152 2836 22158 2848
rect 22741 2839 22799 2845
rect 22741 2836 22753 2839
rect 22152 2808 22753 2836
rect 22152 2796 22158 2808
rect 22741 2805 22753 2808
rect 22787 2805 22799 2839
rect 22741 2799 22799 2805
rect 23198 2796 23204 2848
rect 23256 2836 23262 2848
rect 23477 2839 23535 2845
rect 23477 2836 23489 2839
rect 23256 2808 23489 2836
rect 23256 2796 23262 2808
rect 23477 2805 23489 2808
rect 23523 2805 23535 2839
rect 23477 2799 23535 2805
rect 25406 2796 25412 2848
rect 25464 2836 25470 2848
rect 25593 2839 25651 2845
rect 25593 2836 25605 2839
rect 25464 2808 25605 2836
rect 25464 2796 25470 2808
rect 25593 2805 25605 2808
rect 25639 2805 25651 2839
rect 25593 2799 25651 2805
rect 26510 2796 26516 2848
rect 26568 2836 26574 2848
rect 26697 2839 26755 2845
rect 26697 2836 26709 2839
rect 26568 2808 26709 2836
rect 26568 2796 26574 2808
rect 26697 2805 26709 2808
rect 26743 2805 26755 2839
rect 26697 2799 26755 2805
rect 27614 2796 27620 2848
rect 27672 2836 27678 2848
rect 27985 2839 28043 2845
rect 27985 2836 27997 2839
rect 27672 2808 27997 2836
rect 27672 2796 27678 2808
rect 27985 2805 27997 2808
rect 28031 2805 28043 2839
rect 27985 2799 28043 2805
rect 28718 2796 28724 2848
rect 28776 2836 28782 2848
rect 28905 2839 28963 2845
rect 28905 2836 28917 2839
rect 28776 2808 28917 2836
rect 28776 2796 28782 2808
rect 28905 2805 28917 2808
rect 28951 2805 28963 2839
rect 28905 2799 28963 2805
rect 30926 2796 30932 2848
rect 30984 2836 30990 2848
rect 31113 2839 31171 2845
rect 31113 2836 31125 2839
rect 30984 2808 31125 2836
rect 30984 2796 30990 2808
rect 31113 2805 31125 2808
rect 31159 2805 31171 2839
rect 32030 2836 32036 2848
rect 31991 2808 32036 2836
rect 31113 2799 31171 2805
rect 32030 2796 32036 2808
rect 32088 2796 32094 2848
rect 33134 2796 33140 2848
rect 33192 2836 33198 2848
rect 33321 2839 33379 2845
rect 33321 2836 33333 2839
rect 33192 2808 33333 2836
rect 33192 2796 33198 2808
rect 33321 2805 33333 2808
rect 33367 2805 33379 2839
rect 33321 2799 33379 2805
rect 34238 2796 34244 2848
rect 34296 2836 34302 2848
rect 34425 2839 34483 2845
rect 34425 2836 34437 2839
rect 34296 2808 34437 2836
rect 34296 2796 34302 2808
rect 34425 2805 34437 2808
rect 34471 2805 34483 2839
rect 34425 2799 34483 2805
rect 35342 2796 35348 2848
rect 35400 2836 35406 2848
rect 35529 2839 35587 2845
rect 35529 2836 35541 2839
rect 35400 2808 35541 2836
rect 35400 2796 35406 2808
rect 35529 2805 35541 2808
rect 35575 2805 35587 2839
rect 35529 2799 35587 2805
rect 36446 2796 36452 2848
rect 36504 2836 36510 2848
rect 36633 2839 36691 2845
rect 36633 2836 36645 2839
rect 36504 2808 36645 2836
rect 36504 2796 36510 2808
rect 36633 2805 36645 2808
rect 36679 2805 36691 2839
rect 36633 2799 36691 2805
rect 37550 2796 37556 2848
rect 37608 2836 37614 2848
rect 38473 2839 38531 2845
rect 38473 2836 38485 2839
rect 37608 2808 38485 2836
rect 37608 2796 37614 2808
rect 38473 2805 38485 2808
rect 38519 2805 38531 2839
rect 38473 2799 38531 2805
rect 38654 2796 38660 2848
rect 38712 2836 38718 2848
rect 39209 2839 39267 2845
rect 39209 2836 39221 2839
rect 38712 2808 39221 2836
rect 38712 2796 38718 2808
rect 39209 2805 39221 2808
rect 39255 2805 39267 2839
rect 66088 2836 66116 2867
rect 68572 2836 68600 2944
rect 68646 2864 68652 2916
rect 68704 2904 68710 2916
rect 68704 2876 68749 2904
rect 68704 2864 68710 2876
rect 68830 2836 68836 2848
rect 66088 2808 68600 2836
rect 68791 2808 68836 2836
rect 39209 2799 39267 2805
rect 68830 2796 68836 2808
rect 68888 2796 68894 2848
rect 68940 2836 68968 2944
rect 69753 2941 69765 2975
rect 69799 2972 69811 2975
rect 70857 2975 70915 2981
rect 69799 2944 70394 2972
rect 69799 2941 69811 2944
rect 69753 2935 69811 2941
rect 70210 2913 70216 2916
rect 70167 2907 70216 2913
rect 70167 2873 70179 2907
rect 70213 2873 70216 2907
rect 70167 2867 70216 2873
rect 70210 2864 70216 2867
rect 70268 2864 70274 2916
rect 70366 2904 70394 2944
rect 70857 2941 70869 2975
rect 70903 2941 70915 2975
rect 71501 2975 71559 2981
rect 70857 2935 70915 2941
rect 70964 2944 71452 2972
rect 70964 2904 70992 2944
rect 71314 2913 71320 2916
rect 70366 2876 70992 2904
rect 71271 2907 71320 2913
rect 71271 2873 71283 2907
rect 71317 2873 71320 2907
rect 71271 2867 71320 2873
rect 71314 2864 71320 2867
rect 71372 2864 71378 2916
rect 71424 2904 71452 2944
rect 71501 2941 71513 2975
rect 71547 2972 71559 2975
rect 71590 2972 71596 2984
rect 71547 2944 71596 2972
rect 71547 2941 71559 2944
rect 71501 2935 71559 2941
rect 71590 2932 71596 2944
rect 71648 2932 71654 2984
rect 71961 2975 72019 2981
rect 71961 2941 71973 2975
rect 72007 2972 72019 2975
rect 72142 2972 72148 2984
rect 72007 2944 72148 2972
rect 72007 2941 72019 2944
rect 71961 2935 72019 2941
rect 72142 2932 72148 2944
rect 72200 2932 72206 2984
rect 73614 2932 73620 2984
rect 73672 2972 73678 2984
rect 77205 2975 77263 2981
rect 73672 2944 73717 2972
rect 74920 2944 76788 2972
rect 73672 2932 73678 2944
rect 74920 2904 74948 2944
rect 71424 2876 74948 2904
rect 75365 2907 75423 2913
rect 75365 2873 75377 2907
rect 75411 2904 75423 2907
rect 75454 2904 75460 2916
rect 75411 2876 75460 2904
rect 75411 2873 75423 2876
rect 75365 2867 75423 2873
rect 75454 2864 75460 2876
rect 75512 2864 75518 2916
rect 76377 2907 76435 2913
rect 76377 2873 76389 2907
rect 76423 2904 76435 2907
rect 76650 2904 76656 2916
rect 76423 2876 76656 2904
rect 76423 2873 76435 2876
rect 76377 2867 76435 2873
rect 76650 2864 76656 2876
rect 76708 2864 76714 2916
rect 71590 2836 71596 2848
rect 68940 2808 71596 2836
rect 71590 2796 71596 2808
rect 71648 2796 71654 2848
rect 72329 2839 72387 2845
rect 72329 2805 72341 2839
rect 72375 2836 72387 2839
rect 73430 2836 73436 2848
rect 72375 2808 73436 2836
rect 72375 2805 72387 2808
rect 72329 2799 72387 2805
rect 73430 2796 73436 2808
rect 73488 2796 73494 2848
rect 73522 2796 73528 2848
rect 73580 2836 73586 2848
rect 73709 2839 73767 2845
rect 73709 2836 73721 2839
rect 73580 2808 73721 2836
rect 73580 2796 73586 2808
rect 73709 2805 73721 2808
rect 73755 2805 73767 2839
rect 75546 2836 75552 2848
rect 75507 2808 75552 2836
rect 73709 2799 73767 2805
rect 75546 2796 75552 2808
rect 75604 2796 75610 2848
rect 76760 2836 76788 2944
rect 77205 2941 77217 2975
rect 77251 2972 77263 2975
rect 77570 2972 77576 2984
rect 77251 2944 77576 2972
rect 77251 2941 77263 2944
rect 77205 2935 77263 2941
rect 77570 2932 77576 2944
rect 77628 2932 77634 2984
rect 77665 2975 77723 2981
rect 77665 2941 77677 2975
rect 77711 2972 77723 2975
rect 78950 2972 78956 2984
rect 77711 2944 78956 2972
rect 77711 2941 77723 2944
rect 77665 2935 77723 2941
rect 78950 2932 78956 2944
rect 79008 2932 79014 2984
rect 78033 2907 78091 2913
rect 78033 2873 78045 2907
rect 78079 2904 78091 2907
rect 78766 2904 78772 2916
rect 78079 2876 78772 2904
rect 78079 2873 78091 2876
rect 78033 2867 78091 2873
rect 78766 2864 78772 2876
rect 78824 2864 78830 2916
rect 79042 2904 79048 2916
rect 79003 2876 79048 2904
rect 79042 2864 79048 2876
rect 79100 2864 79106 2916
rect 79152 2836 79180 3012
rect 80054 2932 80060 2984
rect 80112 2972 80118 2984
rect 80241 2975 80299 2981
rect 80241 2972 80253 2975
rect 80112 2944 80253 2972
rect 80112 2932 80118 2944
rect 80241 2941 80253 2944
rect 80287 2941 80299 2975
rect 80241 2935 80299 2941
rect 80330 2932 80336 2984
rect 80388 2972 80394 2984
rect 80425 2975 80483 2981
rect 80425 2972 80437 2975
rect 80388 2944 80437 2972
rect 80388 2932 80394 2944
rect 80425 2941 80437 2944
rect 80471 2941 80483 2975
rect 80425 2935 80483 2941
rect 80517 2975 80575 2981
rect 80517 2941 80529 2975
rect 80563 2972 80575 2975
rect 80698 2972 80704 2984
rect 80563 2944 80704 2972
rect 80563 2941 80575 2944
rect 80517 2935 80575 2941
rect 80698 2932 80704 2944
rect 80756 2932 80762 2984
rect 80793 2975 80851 2981
rect 80793 2941 80805 2975
rect 80839 2972 80851 2975
rect 80882 2972 80888 2984
rect 80839 2944 80888 2972
rect 80839 2941 80851 2944
rect 80793 2935 80851 2941
rect 80882 2932 80888 2944
rect 80940 2932 80946 2984
rect 81452 2981 81480 3012
rect 82078 3000 82084 3012
rect 82136 3000 82142 3052
rect 82354 3000 82360 3052
rect 82412 3040 82418 3052
rect 85761 3043 85819 3049
rect 85761 3040 85773 3043
rect 82412 3012 85773 3040
rect 82412 3000 82418 3012
rect 85761 3009 85773 3012
rect 85807 3009 85819 3043
rect 86506 3043 86564 3049
rect 86506 3040 86518 3043
rect 85761 3003 85819 3009
rect 86328 3012 86518 3040
rect 81437 2975 81495 2981
rect 81437 2941 81449 2975
rect 81483 2941 81495 2975
rect 81437 2935 81495 2941
rect 81526 2932 81532 2984
rect 81584 2972 81590 2984
rect 81805 2975 81863 2981
rect 81584 2944 81629 2972
rect 81584 2932 81590 2944
rect 81805 2941 81817 2975
rect 81851 2972 81863 2975
rect 82170 2972 82176 2984
rect 81851 2944 82176 2972
rect 81851 2941 81863 2944
rect 81805 2935 81863 2941
rect 82170 2932 82176 2944
rect 82228 2932 82234 2984
rect 82262 2932 82268 2984
rect 82320 2972 82326 2984
rect 82449 2975 82507 2981
rect 82320 2944 82365 2972
rect 82320 2932 82326 2944
rect 82449 2941 82461 2975
rect 82495 2941 82507 2975
rect 82449 2935 82507 2941
rect 82464 2904 82492 2935
rect 82538 2932 82544 2984
rect 82596 2972 82602 2984
rect 82633 2975 82691 2981
rect 82633 2972 82645 2975
rect 82596 2944 82645 2972
rect 82596 2932 82602 2944
rect 82633 2941 82645 2944
rect 82679 2941 82691 2975
rect 82814 2972 82820 2984
rect 82775 2944 82820 2972
rect 82633 2935 82691 2941
rect 82814 2932 82820 2944
rect 82872 2932 82878 2984
rect 83553 2975 83611 2981
rect 83553 2941 83565 2975
rect 83599 2941 83611 2975
rect 83734 2972 83740 2984
rect 83695 2944 83740 2972
rect 83553 2935 83611 2941
rect 80072 2876 82492 2904
rect 76760 2808 79180 2836
rect 79229 2839 79287 2845
rect 79229 2805 79241 2839
rect 79275 2836 79287 2839
rect 79318 2836 79324 2848
rect 79275 2808 79324 2836
rect 79275 2805 79287 2808
rect 79229 2799 79287 2805
rect 79318 2796 79324 2808
rect 79376 2796 79382 2848
rect 79686 2796 79692 2848
rect 79744 2836 79750 2848
rect 80072 2836 80100 2876
rect 82722 2864 82728 2916
rect 82780 2904 82786 2916
rect 82998 2904 83004 2916
rect 82780 2876 83004 2904
rect 82780 2864 82786 2876
rect 82998 2864 83004 2876
rect 83056 2864 83062 2916
rect 79744 2808 80100 2836
rect 79744 2796 79750 2808
rect 80422 2796 80428 2848
rect 80480 2836 80486 2848
rect 82078 2836 82084 2848
rect 80480 2808 82084 2836
rect 80480 2796 80486 2808
rect 82078 2796 82084 2808
rect 82136 2796 82142 2848
rect 82170 2796 82176 2848
rect 82228 2836 82234 2848
rect 82630 2836 82636 2848
rect 82228 2808 82636 2836
rect 82228 2796 82234 2808
rect 82630 2796 82636 2808
rect 82688 2796 82694 2848
rect 83568 2836 83596 2935
rect 83734 2932 83740 2944
rect 83792 2932 83798 2984
rect 83829 2975 83887 2981
rect 83829 2941 83841 2975
rect 83875 2972 83887 2975
rect 83921 2975 83979 2981
rect 83921 2972 83933 2975
rect 83875 2944 83933 2972
rect 83875 2941 83887 2944
rect 83829 2935 83887 2941
rect 83921 2941 83933 2944
rect 83967 2941 83979 2975
rect 83921 2935 83979 2941
rect 83936 2904 83964 2935
rect 84010 2932 84016 2984
rect 84068 2972 84074 2984
rect 84105 2975 84163 2981
rect 84105 2972 84117 2975
rect 84068 2944 84117 2972
rect 84068 2932 84074 2944
rect 84105 2941 84117 2944
rect 84151 2941 84163 2975
rect 84105 2935 84163 2941
rect 84286 2932 84292 2984
rect 84344 2932 84350 2984
rect 84654 2932 84660 2984
rect 84712 2972 84718 2984
rect 84712 2944 85804 2972
rect 84712 2932 84718 2944
rect 84304 2904 84332 2932
rect 83936 2876 84332 2904
rect 85298 2864 85304 2916
rect 85356 2904 85362 2916
rect 85577 2907 85635 2913
rect 85577 2904 85589 2907
rect 85356 2876 85589 2904
rect 85356 2864 85362 2876
rect 85577 2873 85589 2876
rect 85623 2873 85635 2907
rect 85776 2904 85804 2944
rect 85850 2932 85856 2984
rect 85908 2972 85914 2984
rect 86221 2975 86279 2981
rect 86221 2972 86233 2975
rect 85908 2944 86233 2972
rect 85908 2932 85914 2944
rect 86221 2941 86233 2944
rect 86267 2941 86279 2975
rect 86221 2935 86279 2941
rect 86328 2904 86356 3012
rect 86506 3009 86518 3012
rect 86552 3009 86564 3043
rect 86506 3003 86564 3009
rect 86393 2975 86451 2981
rect 86393 2941 86405 2975
rect 86439 2941 86451 2975
rect 86586 2972 86592 2984
rect 86547 2944 86592 2972
rect 86393 2935 86451 2941
rect 85776 2876 86356 2904
rect 86420 2904 86448 2935
rect 86586 2932 86592 2944
rect 86644 2932 86650 2984
rect 86770 2972 86776 2984
rect 86731 2944 86776 2972
rect 86770 2932 86776 2944
rect 86828 2932 86834 2984
rect 87616 2981 87644 3080
rect 90913 3077 90925 3111
rect 90959 3108 90971 3111
rect 93118 3108 93124 3120
rect 90959 3080 93124 3108
rect 90959 3077 90971 3080
rect 90913 3071 90971 3077
rect 93118 3068 93124 3080
rect 93176 3068 93182 3120
rect 93302 3068 93308 3120
rect 93360 3108 93366 3120
rect 99024 3108 99052 3148
rect 100478 3136 100484 3148
rect 100536 3136 100542 3188
rect 101674 3136 101680 3188
rect 101732 3176 101738 3188
rect 110601 3179 110659 3185
rect 110601 3176 110613 3179
rect 101732 3148 110613 3176
rect 101732 3136 101738 3148
rect 110601 3145 110613 3148
rect 110647 3145 110659 3179
rect 110601 3139 110659 3145
rect 103882 3108 103888 3120
rect 93360 3080 99052 3108
rect 99346 3080 103888 3108
rect 93360 3068 93366 3080
rect 91557 3043 91615 3049
rect 91557 3009 91569 3043
rect 91603 3040 91615 3043
rect 93210 3040 93216 3052
rect 91603 3012 93216 3040
rect 91603 3009 91615 3012
rect 91557 3003 91615 3009
rect 93210 3000 93216 3012
rect 93268 3000 93274 3052
rect 93578 3000 93584 3052
rect 93636 3040 93642 3052
rect 96801 3043 96859 3049
rect 93636 3012 96752 3040
rect 93636 3000 93642 3012
rect 87601 2975 87659 2981
rect 87601 2941 87613 2975
rect 87647 2941 87659 2975
rect 87601 2935 87659 2941
rect 87690 2932 87696 2984
rect 87748 2972 87754 2984
rect 87966 2981 87972 2984
rect 87951 2975 87972 2981
rect 87748 2944 87793 2972
rect 87748 2932 87754 2944
rect 87951 2941 87963 2975
rect 87951 2935 87972 2941
rect 87966 2932 87972 2935
rect 88024 2932 88030 2984
rect 88150 2932 88156 2984
rect 88208 2972 88214 2984
rect 88334 2972 88340 2984
rect 88208 2944 88340 2972
rect 88208 2932 88214 2944
rect 88334 2932 88340 2944
rect 88392 2972 88398 2984
rect 88429 2975 88487 2981
rect 88429 2972 88441 2975
rect 88392 2944 88441 2972
rect 88392 2932 88398 2944
rect 88429 2941 88441 2944
rect 88475 2941 88487 2975
rect 88429 2935 88487 2941
rect 89438 2932 89444 2984
rect 89496 2972 89502 2984
rect 89533 2975 89591 2981
rect 89533 2972 89545 2975
rect 89496 2944 89545 2972
rect 89496 2932 89502 2944
rect 89533 2941 89545 2944
rect 89579 2941 89591 2975
rect 89533 2935 89591 2941
rect 92293 2975 92351 2981
rect 92293 2941 92305 2975
rect 92339 2972 92351 2975
rect 93302 2972 93308 2984
rect 92339 2944 93308 2972
rect 92339 2941 92351 2944
rect 92293 2935 92351 2941
rect 93302 2932 93308 2944
rect 93360 2932 93366 2984
rect 93397 2975 93455 2981
rect 93397 2941 93409 2975
rect 93443 2972 93455 2975
rect 94406 2972 94412 2984
rect 93443 2944 94412 2972
rect 93443 2941 93455 2944
rect 93397 2935 93455 2941
rect 94406 2932 94412 2944
rect 94464 2932 94470 2984
rect 94501 2975 94559 2981
rect 94501 2941 94513 2975
rect 94547 2972 94559 2975
rect 96062 2972 96068 2984
rect 94547 2944 96068 2972
rect 94547 2941 94559 2944
rect 94501 2935 94559 2941
rect 96062 2932 96068 2944
rect 96120 2932 96126 2984
rect 96157 2975 96215 2981
rect 96157 2941 96169 2975
rect 96203 2972 96215 2975
rect 96614 2972 96620 2984
rect 96203 2944 96620 2972
rect 96203 2941 96215 2944
rect 96157 2935 96215 2941
rect 96614 2932 96620 2944
rect 96672 2932 96678 2984
rect 96724 2972 96752 3012
rect 96801 3009 96813 3043
rect 96847 3040 96859 3043
rect 98454 3040 98460 3052
rect 96847 3012 98460 3040
rect 96847 3009 96859 3012
rect 96801 3003 96859 3009
rect 98454 3000 98460 3012
rect 98512 3000 98518 3052
rect 99346 3040 99374 3080
rect 103882 3068 103888 3080
rect 103940 3068 103946 3120
rect 101306 3040 101312 3052
rect 98840 3012 99374 3040
rect 101267 3012 101312 3040
rect 97813 2975 97871 2981
rect 96724 2944 97396 2972
rect 86494 2904 86500 2916
rect 86420 2876 86500 2904
rect 85577 2867 85635 2873
rect 86494 2864 86500 2876
rect 86552 2864 86558 2916
rect 86862 2864 86868 2916
rect 86920 2904 86926 2916
rect 87417 2907 87475 2913
rect 87417 2904 87429 2907
rect 86920 2876 87429 2904
rect 86920 2864 86926 2876
rect 87417 2873 87429 2876
rect 87463 2873 87475 2907
rect 87417 2867 87475 2873
rect 92198 2864 92204 2916
rect 92256 2904 92262 2916
rect 92256 2876 92704 2904
rect 92256 2864 92262 2876
rect 84286 2836 84292 2848
rect 83568 2808 84292 2836
rect 84286 2796 84292 2808
rect 84344 2796 84350 2848
rect 85482 2796 85488 2848
rect 85540 2836 85546 2848
rect 86586 2836 86592 2848
rect 85540 2808 86592 2836
rect 85540 2796 85546 2808
rect 86586 2796 86592 2808
rect 86644 2796 86650 2848
rect 86678 2796 86684 2848
rect 86736 2836 86742 2848
rect 87690 2836 87696 2848
rect 86736 2808 87696 2836
rect 86736 2796 86742 2808
rect 87690 2796 87696 2808
rect 87748 2796 87754 2848
rect 88426 2796 88432 2848
rect 88484 2836 88490 2848
rect 88797 2839 88855 2845
rect 88797 2836 88809 2839
rect 88484 2808 88809 2836
rect 88484 2796 88490 2808
rect 88797 2805 88809 2808
rect 88843 2805 88855 2839
rect 88797 2799 88855 2805
rect 88886 2796 88892 2848
rect 88944 2836 88950 2848
rect 88981 2839 89039 2845
rect 88981 2836 88993 2839
rect 88944 2808 88993 2836
rect 88944 2796 88950 2808
rect 88981 2805 88993 2808
rect 89027 2805 89039 2839
rect 88981 2799 89039 2805
rect 89162 2796 89168 2848
rect 89220 2836 89226 2848
rect 89625 2839 89683 2845
rect 89625 2836 89637 2839
rect 89220 2808 89637 2836
rect 89220 2796 89226 2808
rect 89625 2805 89637 2808
rect 89671 2805 89683 2839
rect 89625 2799 89683 2805
rect 90082 2796 90088 2848
rect 90140 2836 90146 2848
rect 92566 2836 92572 2848
rect 90140 2808 92572 2836
rect 90140 2796 90146 2808
rect 92566 2796 92572 2808
rect 92624 2796 92630 2848
rect 92676 2836 92704 2876
rect 92750 2864 92756 2916
rect 92808 2904 92814 2916
rect 97258 2904 97264 2916
rect 92808 2876 97264 2904
rect 92808 2864 92814 2876
rect 97258 2864 97264 2876
rect 97316 2864 97322 2916
rect 97368 2904 97396 2944
rect 97813 2941 97825 2975
rect 97859 2972 97871 2975
rect 98730 2972 98736 2984
rect 97859 2944 98736 2972
rect 97859 2941 97871 2944
rect 97813 2935 97871 2941
rect 98730 2932 98736 2944
rect 98788 2932 98794 2984
rect 98840 2904 98868 3012
rect 101306 3000 101312 3012
rect 101364 3000 101370 3052
rect 102134 3000 102140 3052
rect 102192 3000 102198 3052
rect 107470 3040 107476 3052
rect 103086 3012 107476 3040
rect 107470 3000 107476 3012
rect 107528 3000 107534 3052
rect 107749 3043 107807 3049
rect 107749 3009 107761 3043
rect 107795 3040 107807 3043
rect 109126 3040 109132 3052
rect 107795 3012 109132 3040
rect 107795 3009 107807 3012
rect 107749 3003 107807 3009
rect 109126 3000 109132 3012
rect 109184 3000 109190 3052
rect 109957 3043 110015 3049
rect 109957 3009 109969 3043
rect 110003 3040 110015 3043
rect 111610 3040 111616 3052
rect 110003 3012 111616 3040
rect 110003 3009 110015 3012
rect 109957 3003 110015 3009
rect 111610 3000 111616 3012
rect 111668 3000 111674 3052
rect 98917 2975 98975 2981
rect 98917 2941 98929 2975
rect 98963 2972 98975 2975
rect 99926 2972 99932 2984
rect 98963 2944 99932 2972
rect 98963 2941 98975 2944
rect 98917 2935 98975 2941
rect 99926 2932 99932 2944
rect 99984 2932 99990 2984
rect 100021 2975 100079 2981
rect 100021 2941 100033 2975
rect 100067 2972 100079 2975
rect 101122 2972 101128 2984
rect 100067 2944 101128 2972
rect 100067 2941 100079 2944
rect 100021 2935 100079 2941
rect 101122 2932 101128 2944
rect 101180 2932 101186 2984
rect 102152 2958 102180 3000
rect 103698 2972 103704 2984
rect 103659 2944 103704 2972
rect 103698 2932 103704 2944
rect 103756 2932 103762 2984
rect 104434 2972 104440 2984
rect 104395 2944 104440 2972
rect 104434 2932 104440 2944
rect 104492 2932 104498 2984
rect 105538 2972 105544 2984
rect 105499 2944 105544 2972
rect 105538 2932 105544 2944
rect 105596 2932 105602 2984
rect 106642 2972 106648 2984
rect 106603 2944 106648 2972
rect 106642 2932 106648 2944
rect 106700 2932 106706 2984
rect 108853 2975 108911 2981
rect 108853 2941 108865 2975
rect 108899 2972 108911 2975
rect 109862 2972 109868 2984
rect 108899 2944 109868 2972
rect 108899 2941 108911 2944
rect 108853 2935 108911 2941
rect 109862 2932 109868 2944
rect 109920 2932 109926 2984
rect 110417 2975 110475 2981
rect 110417 2941 110429 2975
rect 110463 2941 110475 2975
rect 110417 2935 110475 2941
rect 111889 2975 111947 2981
rect 111889 2941 111901 2975
rect 111935 2972 111947 2975
rect 112438 2972 112444 2984
rect 111935 2944 112444 2972
rect 111935 2941 111947 2944
rect 111889 2935 111947 2941
rect 97368 2876 98868 2904
rect 102870 2864 102876 2916
rect 102928 2904 102934 2916
rect 107194 2904 107200 2916
rect 102928 2876 107200 2904
rect 102928 2864 102934 2876
rect 107194 2864 107200 2876
rect 107252 2864 107258 2916
rect 109586 2864 109592 2916
rect 109644 2904 109650 2916
rect 110432 2904 110460 2935
rect 112438 2932 112444 2944
rect 112496 2932 112502 2984
rect 112533 2975 112591 2981
rect 112533 2941 112545 2975
rect 112579 2972 112591 2975
rect 113174 2972 113180 2984
rect 112579 2944 113180 2972
rect 112579 2941 112591 2944
rect 112533 2935 112591 2941
rect 113174 2932 113180 2944
rect 113232 2932 113238 2984
rect 113269 2975 113327 2981
rect 113269 2941 113281 2975
rect 113315 2972 113327 2975
rect 114278 2972 114284 2984
rect 113315 2944 114284 2972
rect 113315 2941 113327 2944
rect 113269 2935 113327 2941
rect 114278 2932 114284 2944
rect 114336 2932 114342 2984
rect 114373 2975 114431 2981
rect 114373 2941 114385 2975
rect 114419 2972 114431 2975
rect 115198 2972 115204 2984
rect 114419 2944 115204 2972
rect 114419 2941 114431 2944
rect 114373 2935 114431 2941
rect 115198 2932 115204 2944
rect 115256 2932 115262 2984
rect 115477 2975 115535 2981
rect 115477 2941 115489 2975
rect 115523 2972 115535 2975
rect 116394 2972 116400 2984
rect 115523 2944 116400 2972
rect 115523 2941 115535 2944
rect 115477 2935 115535 2941
rect 116394 2932 116400 2944
rect 116452 2932 116458 2984
rect 117130 2972 117136 2984
rect 117091 2944 117136 2972
rect 117130 2932 117136 2944
rect 117188 2932 117194 2984
rect 117774 2972 117780 2984
rect 117735 2944 117780 2972
rect 117774 2932 117780 2944
rect 117832 2932 117838 2984
rect 118786 2972 118792 2984
rect 118747 2944 118792 2972
rect 118786 2932 118792 2944
rect 118844 2932 118850 2984
rect 119890 2972 119896 2984
rect 119851 2944 119896 2972
rect 119890 2932 119896 2944
rect 119948 2932 119954 2984
rect 120905 2975 120963 2981
rect 120905 2941 120917 2975
rect 120951 2972 120963 2975
rect 121730 2972 121736 2984
rect 120951 2944 121736 2972
rect 120951 2941 120963 2944
rect 120905 2935 120963 2941
rect 121730 2932 121736 2944
rect 121788 2932 121794 2984
rect 122374 2972 122380 2984
rect 122335 2944 122380 2972
rect 122374 2932 122380 2944
rect 122432 2932 122438 2984
rect 123110 2972 123116 2984
rect 123071 2944 123116 2972
rect 123110 2932 123116 2944
rect 123168 2932 123174 2984
rect 124214 2972 124220 2984
rect 124175 2944 124220 2972
rect 124214 2932 124220 2944
rect 124272 2932 124278 2984
rect 125318 2972 125324 2984
rect 125279 2944 125324 2972
rect 125318 2932 125324 2944
rect 125376 2932 125382 2984
rect 126425 2975 126483 2981
rect 126425 2941 126437 2975
rect 126471 2972 126483 2975
rect 127066 2972 127072 2984
rect 126471 2944 127072 2972
rect 126471 2941 126483 2944
rect 126425 2935 126483 2941
rect 127066 2932 127072 2944
rect 127124 2932 127130 2984
rect 127618 2972 127624 2984
rect 127579 2944 127624 2972
rect 127618 2932 127624 2944
rect 127676 2932 127682 2984
rect 128630 2972 128636 2984
rect 128591 2944 128636 2972
rect 128630 2932 128636 2944
rect 128688 2932 128694 2984
rect 129734 2972 129740 2984
rect 129695 2944 129740 2972
rect 129734 2932 129740 2944
rect 129792 2932 129798 2984
rect 130838 2972 130844 2984
rect 130799 2944 130844 2972
rect 130838 2932 130844 2944
rect 130896 2932 130902 2984
rect 131301 2975 131359 2981
rect 131301 2941 131313 2975
rect 131347 2941 131359 2975
rect 133046 2972 133052 2984
rect 133007 2944 133052 2972
rect 131301 2935 131359 2941
rect 109644 2876 110460 2904
rect 109644 2864 109650 2876
rect 130470 2864 130476 2916
rect 130528 2904 130534 2916
rect 131316 2904 131344 2935
rect 133046 2932 133052 2944
rect 133104 2932 133110 2984
rect 134150 2972 134156 2984
rect 134111 2944 134156 2972
rect 134150 2932 134156 2944
rect 134208 2932 134214 2984
rect 135254 2972 135260 2984
rect 135215 2944 135260 2972
rect 135254 2932 135260 2944
rect 135312 2932 135318 2984
rect 136358 2972 136364 2984
rect 136319 2944 136364 2972
rect 136358 2932 136364 2944
rect 136416 2932 136422 2984
rect 136821 2975 136879 2981
rect 136821 2941 136833 2975
rect 136867 2941 136879 2975
rect 138106 2972 138112 2984
rect 138067 2944 138112 2972
rect 136821 2935 136879 2941
rect 130528 2876 131344 2904
rect 130528 2864 130534 2876
rect 135990 2864 135996 2916
rect 136048 2904 136054 2916
rect 136836 2904 136864 2935
rect 138106 2932 138112 2944
rect 138164 2932 138170 2984
rect 138750 2972 138756 2984
rect 138711 2944 138756 2972
rect 138750 2932 138756 2944
rect 138808 2932 138814 2984
rect 139670 2972 139676 2984
rect 139631 2944 139676 2972
rect 139670 2932 139676 2944
rect 139728 2932 139734 2984
rect 140774 2972 140780 2984
rect 140735 2944 140780 2972
rect 140774 2932 140780 2944
rect 140832 2932 140838 2984
rect 141878 2972 141884 2984
rect 141839 2944 141884 2972
rect 141878 2932 141884 2944
rect 141936 2932 141942 2984
rect 143350 2972 143356 2984
rect 143311 2944 143356 2972
rect 143350 2932 143356 2944
rect 143408 2932 143414 2984
rect 144086 2972 144092 2984
rect 144047 2944 144092 2972
rect 144086 2932 144092 2944
rect 144144 2932 144150 2984
rect 145190 2972 145196 2984
rect 145151 2944 145196 2972
rect 145190 2932 145196 2944
rect 145248 2932 145254 2984
rect 146294 2972 146300 2984
rect 146255 2944 146300 2972
rect 146294 2932 146300 2944
rect 146352 2932 146358 2984
rect 147398 2972 147404 2984
rect 147359 2944 147404 2972
rect 147398 2932 147404 2944
rect 147456 2932 147462 2984
rect 148594 2972 148600 2984
rect 148555 2944 148600 2972
rect 148594 2932 148600 2944
rect 148652 2932 148658 2984
rect 149606 2972 149612 2984
rect 149567 2944 149612 2972
rect 149606 2932 149612 2944
rect 149664 2932 149670 2984
rect 150710 2972 150716 2984
rect 150671 2944 150716 2972
rect 150710 2932 150716 2944
rect 150768 2932 150774 2984
rect 151814 2932 151820 2984
rect 151872 2972 151878 2984
rect 152550 2972 152556 2984
rect 151872 2944 151917 2972
rect 152511 2944 152556 2972
rect 151872 2932 151878 2944
rect 152550 2932 152556 2944
rect 152608 2932 152614 2984
rect 154022 2972 154028 2984
rect 153983 2944 154028 2972
rect 154022 2932 154028 2944
rect 154080 2932 154086 2984
rect 155126 2972 155132 2984
rect 155087 2944 155132 2972
rect 155126 2932 155132 2944
rect 155184 2932 155190 2984
rect 156230 2972 156236 2984
rect 156191 2944 156236 2972
rect 156230 2932 156236 2944
rect 156288 2932 156294 2984
rect 157334 2972 157340 2984
rect 157295 2944 157340 2972
rect 157334 2932 157340 2944
rect 157392 2932 157398 2984
rect 157797 2975 157855 2981
rect 157797 2941 157809 2975
rect 157843 2941 157855 2975
rect 159082 2972 159088 2984
rect 159043 2944 159088 2972
rect 157797 2935 157855 2941
rect 136048 2876 136864 2904
rect 136048 2864 136054 2876
rect 156966 2864 156972 2916
rect 157024 2904 157030 2916
rect 157812 2904 157840 2935
rect 159082 2932 159088 2944
rect 159140 2932 159146 2984
rect 159726 2972 159732 2984
rect 159687 2944 159732 2972
rect 159726 2932 159732 2944
rect 159784 2932 159790 2984
rect 160646 2972 160652 2984
rect 160607 2944 160652 2972
rect 160646 2932 160652 2944
rect 160704 2932 160710 2984
rect 161750 2972 161756 2984
rect 161711 2944 161756 2972
rect 161750 2932 161756 2944
rect 161808 2932 161814 2984
rect 162854 2972 162860 2984
rect 162815 2944 162860 2972
rect 162854 2932 162860 2944
rect 162912 2932 162918 2984
rect 164326 2972 164332 2984
rect 164287 2944 164332 2972
rect 164326 2932 164332 2944
rect 164384 2932 164390 2984
rect 165062 2972 165068 2984
rect 165023 2944 165068 2972
rect 165062 2932 165068 2944
rect 165120 2932 165126 2984
rect 166169 2975 166227 2981
rect 166169 2941 166181 2975
rect 166215 2972 166227 2975
rect 167086 2972 167092 2984
rect 166215 2944 167092 2972
rect 166215 2941 166227 2944
rect 166169 2935 166227 2941
rect 167086 2932 167092 2944
rect 167144 2932 167150 2984
rect 167270 2972 167276 2984
rect 167231 2944 167276 2972
rect 167270 2932 167276 2944
rect 167328 2932 167334 2984
rect 168374 2972 168380 2984
rect 168335 2944 168380 2972
rect 168374 2932 168380 2944
rect 168432 2932 168438 2984
rect 169573 2975 169631 2981
rect 169573 2941 169585 2975
rect 169619 2972 169631 2975
rect 169754 2972 169760 2984
rect 169619 2944 169760 2972
rect 169619 2941 169631 2944
rect 169573 2935 169631 2941
rect 169754 2932 169760 2944
rect 169812 2932 169818 2984
rect 170582 2972 170588 2984
rect 170543 2944 170588 2972
rect 170582 2932 170588 2944
rect 170640 2932 170646 2984
rect 171686 2972 171692 2984
rect 171647 2944 171692 2972
rect 171686 2932 171692 2944
rect 171744 2932 171750 2984
rect 172790 2972 172796 2984
rect 172751 2944 172796 2972
rect 172790 2932 172796 2944
rect 172848 2932 172854 2984
rect 173253 2975 173311 2981
rect 173253 2941 173265 2975
rect 173299 2941 173311 2975
rect 174998 2972 175004 2984
rect 174959 2944 175004 2972
rect 173253 2935 173311 2941
rect 157024 2876 157840 2904
rect 157024 2864 157030 2876
rect 172422 2864 172428 2916
rect 172480 2904 172486 2916
rect 173268 2904 173296 2935
rect 174998 2932 175004 2944
rect 175056 2932 175062 2984
rect 176102 2972 176108 2984
rect 176063 2944 176108 2972
rect 176102 2932 176108 2944
rect 176160 2932 176166 2984
rect 176930 2972 176936 2984
rect 176891 2944 176936 2972
rect 176930 2932 176936 2944
rect 176988 2932 176994 2984
rect 177298 2932 177304 2984
rect 177356 2972 177362 2984
rect 177945 2975 178003 2981
rect 177945 2972 177957 2975
rect 177356 2944 177957 2972
rect 177356 2932 177362 2944
rect 177945 2941 177957 2944
rect 177991 2941 178003 2975
rect 177945 2935 178003 2941
rect 172480 2876 173296 2904
rect 178129 2907 178187 2913
rect 172480 2864 172486 2876
rect 178129 2873 178141 2907
rect 178175 2904 178187 2907
rect 178310 2904 178316 2916
rect 178175 2876 178316 2904
rect 178175 2873 178187 2876
rect 178129 2867 178187 2873
rect 178310 2864 178316 2876
rect 178368 2864 178374 2916
rect 98822 2836 98828 2848
rect 92676 2808 98828 2836
rect 98822 2796 98828 2808
rect 98880 2796 98886 2848
rect 102318 2836 102324 2848
rect 102279 2808 102324 2836
rect 102318 2796 102324 2808
rect 102376 2796 102382 2848
rect 102502 2796 102508 2848
rect 102560 2836 102566 2848
rect 107286 2836 107292 2848
rect 102560 2808 107292 2836
rect 102560 2796 102566 2808
rect 107286 2796 107292 2808
rect 107344 2796 107350 2848
rect 1104 2746 178848 2768
rect 1104 2694 19606 2746
rect 19658 2694 19670 2746
rect 19722 2694 19734 2746
rect 19786 2694 19798 2746
rect 19850 2694 50326 2746
rect 50378 2694 50390 2746
rect 50442 2694 50454 2746
rect 50506 2694 50518 2746
rect 50570 2694 81046 2746
rect 81098 2694 81110 2746
rect 81162 2694 81174 2746
rect 81226 2694 81238 2746
rect 81290 2694 111766 2746
rect 111818 2694 111830 2746
rect 111882 2694 111894 2746
rect 111946 2694 111958 2746
rect 112010 2694 142486 2746
rect 142538 2694 142550 2746
rect 142602 2694 142614 2746
rect 142666 2694 142678 2746
rect 142730 2694 173206 2746
rect 173258 2694 173270 2746
rect 173322 2694 173334 2746
rect 173386 2694 173398 2746
rect 173450 2694 178848 2746
rect 1104 2672 178848 2694
rect 7374 2592 7380 2644
rect 7432 2632 7438 2644
rect 10505 2635 10563 2641
rect 10505 2632 10517 2635
rect 7432 2604 10517 2632
rect 7432 2592 7438 2604
rect 10505 2601 10517 2604
rect 10551 2601 10563 2635
rect 18598 2632 18604 2644
rect 10505 2595 10563 2601
rect 11164 2604 18604 2632
rect 5810 2564 5816 2576
rect 5771 2536 5816 2564
rect 5810 2524 5816 2536
rect 5868 2524 5874 2576
rect 11164 2573 11192 2604
rect 18598 2592 18604 2604
rect 18656 2592 18662 2644
rect 37274 2632 37280 2644
rect 31726 2604 37280 2632
rect 11149 2567 11207 2573
rect 11149 2533 11161 2567
rect 11195 2533 11207 2567
rect 31726 2564 31754 2604
rect 37274 2592 37280 2604
rect 37332 2592 37338 2644
rect 37369 2635 37427 2641
rect 37369 2601 37381 2635
rect 37415 2632 37427 2635
rect 65334 2632 65340 2644
rect 37415 2604 65340 2632
rect 37415 2601 37427 2604
rect 37369 2595 37427 2601
rect 65334 2592 65340 2604
rect 65392 2592 65398 2644
rect 71130 2632 71136 2644
rect 70366 2604 71136 2632
rect 11149 2527 11207 2533
rect 11348 2536 13124 2564
rect 106 2456 112 2508
rect 164 2496 170 2508
rect 1397 2499 1455 2505
rect 1397 2496 1409 2499
rect 164 2468 1409 2496
rect 164 2456 170 2468
rect 1397 2465 1409 2468
rect 1443 2465 1455 2499
rect 1670 2496 1676 2508
rect 1631 2468 1676 2496
rect 1397 2459 1455 2465
rect 1670 2456 1676 2468
rect 1728 2456 1734 2508
rect 2590 2456 2596 2508
rect 2648 2496 2654 2508
rect 2685 2499 2743 2505
rect 2685 2496 2697 2499
rect 2648 2468 2697 2496
rect 2648 2456 2654 2468
rect 2685 2465 2697 2468
rect 2731 2465 2743 2499
rect 2685 2459 2743 2465
rect 4062 2456 4068 2508
rect 4120 2496 4126 2508
rect 4341 2499 4399 2505
rect 4341 2496 4353 2499
rect 4120 2468 4353 2496
rect 4120 2456 4126 2468
rect 4341 2465 4353 2468
rect 4387 2465 4399 2499
rect 4341 2459 4399 2465
rect 5534 2456 5540 2508
rect 5592 2496 5598 2508
rect 5629 2499 5687 2505
rect 5629 2496 5641 2499
rect 5592 2468 5641 2496
rect 5592 2456 5598 2468
rect 5629 2465 5641 2468
rect 5675 2465 5687 2499
rect 5629 2459 5687 2465
rect 7006 2456 7012 2508
rect 7064 2496 7070 2508
rect 7101 2499 7159 2505
rect 7101 2496 7113 2499
rect 7064 2468 7113 2496
rect 7064 2456 7070 2468
rect 7101 2465 7113 2468
rect 7147 2465 7159 2499
rect 7101 2459 7159 2465
rect 7745 2499 7803 2505
rect 7745 2465 7757 2499
rect 7791 2496 7803 2499
rect 8110 2496 8116 2508
rect 7791 2468 8116 2496
rect 7791 2465 7803 2468
rect 7745 2459 7803 2465
rect 8110 2456 8116 2468
rect 8168 2456 8174 2508
rect 8478 2496 8484 2508
rect 8439 2468 8484 2496
rect 8478 2456 8484 2468
rect 8536 2456 8542 2508
rect 9674 2496 9680 2508
rect 9635 2468 9680 2496
rect 9674 2456 9680 2468
rect 9732 2456 9738 2508
rect 10413 2499 10471 2505
rect 10413 2465 10425 2499
rect 10459 2496 10471 2499
rect 11348 2496 11376 2536
rect 10459 2468 11376 2496
rect 10459 2465 10471 2468
rect 10413 2459 10471 2465
rect 11422 2456 11428 2508
rect 11480 2496 11486 2508
rect 12253 2499 12311 2505
rect 12253 2496 12265 2499
rect 11480 2468 12265 2496
rect 11480 2456 11486 2468
rect 12253 2465 12265 2468
rect 12299 2465 12311 2499
rect 12253 2459 12311 2465
rect 5902 2388 5908 2440
rect 5960 2428 5966 2440
rect 9861 2431 9919 2437
rect 9861 2428 9873 2431
rect 5960 2400 9873 2428
rect 5960 2388 5966 2400
rect 9861 2397 9873 2400
rect 9907 2397 9919 2431
rect 12894 2428 12900 2440
rect 12855 2400 12900 2428
rect 9861 2391 9919 2397
rect 12894 2388 12900 2400
rect 12952 2388 12958 2440
rect 13096 2428 13124 2536
rect 13188 2536 31754 2564
rect 31941 2567 31999 2573
rect 13188 2505 13216 2536
rect 31941 2533 31953 2567
rect 31987 2564 31999 2567
rect 32122 2564 32128 2576
rect 31987 2536 32128 2564
rect 31987 2533 31999 2536
rect 31941 2527 31999 2533
rect 32122 2524 32128 2536
rect 32180 2524 32186 2576
rect 36538 2524 36544 2576
rect 36596 2564 36602 2576
rect 39761 2567 39819 2573
rect 39761 2564 39773 2567
rect 36596 2536 39773 2564
rect 36596 2524 36602 2536
rect 39761 2533 39773 2536
rect 39807 2533 39819 2567
rect 40494 2564 40500 2576
rect 40455 2536 40500 2564
rect 39761 2527 39819 2533
rect 40494 2524 40500 2536
rect 40552 2524 40558 2576
rect 41138 2524 41144 2576
rect 41196 2564 41202 2576
rect 45094 2564 45100 2576
rect 41196 2536 42932 2564
rect 45055 2536 45100 2564
rect 41196 2524 41202 2536
rect 13173 2499 13231 2505
rect 13173 2465 13185 2499
rect 13219 2465 13231 2499
rect 13173 2459 13231 2465
rect 15102 2456 15108 2508
rect 15160 2496 15166 2508
rect 15197 2499 15255 2505
rect 15197 2496 15209 2499
rect 15160 2468 15209 2496
rect 15160 2456 15166 2468
rect 15197 2465 15209 2468
rect 15243 2465 15255 2499
rect 15197 2459 15255 2465
rect 16206 2456 16212 2508
rect 16264 2496 16270 2508
rect 16301 2499 16359 2505
rect 16301 2496 16313 2499
rect 16264 2468 16313 2496
rect 16264 2456 16270 2468
rect 16301 2465 16313 2468
rect 16347 2465 16359 2499
rect 16301 2459 16359 2465
rect 17310 2456 17316 2508
rect 17368 2496 17374 2508
rect 17681 2499 17739 2505
rect 17681 2496 17693 2499
rect 17368 2468 17693 2496
rect 17368 2456 17374 2468
rect 17681 2465 17693 2468
rect 17727 2465 17739 2499
rect 17681 2459 17739 2465
rect 18693 2499 18751 2505
rect 18693 2465 18705 2499
rect 18739 2496 18751 2499
rect 18739 2468 21680 2496
rect 18739 2465 18751 2468
rect 18693 2459 18751 2465
rect 17954 2428 17960 2440
rect 13096 2400 17960 2428
rect 17954 2388 17960 2400
rect 18012 2388 18018 2440
rect 18414 2428 18420 2440
rect 18375 2400 18420 2428
rect 18414 2388 18420 2400
rect 18472 2388 18478 2440
rect 19518 2388 19524 2440
rect 19576 2428 19582 2440
rect 20257 2431 20315 2437
rect 20257 2428 20269 2431
rect 19576 2400 20269 2428
rect 19576 2388 19582 2400
rect 20257 2397 20269 2400
rect 20303 2397 20315 2431
rect 20530 2428 20536 2440
rect 20491 2400 20536 2428
rect 20257 2391 20315 2397
rect 20530 2388 20536 2400
rect 20588 2388 20594 2440
rect 21652 2428 21680 2468
rect 21726 2456 21732 2508
rect 21784 2496 21790 2508
rect 21821 2499 21879 2505
rect 21821 2496 21833 2499
rect 21784 2468 21833 2496
rect 21784 2456 21790 2468
rect 21821 2465 21833 2468
rect 21867 2465 21879 2499
rect 21821 2459 21879 2465
rect 22830 2456 22836 2508
rect 22888 2496 22894 2508
rect 23017 2499 23075 2505
rect 23017 2496 23029 2499
rect 22888 2468 23029 2496
rect 22888 2456 22894 2468
rect 23017 2465 23029 2468
rect 23063 2465 23075 2499
rect 23017 2459 23075 2465
rect 23934 2456 23940 2508
rect 23992 2496 23998 2508
rect 24029 2499 24087 2505
rect 24029 2496 24041 2499
rect 23992 2468 24041 2496
rect 23992 2456 23998 2468
rect 24029 2465 24041 2468
rect 24075 2465 24087 2499
rect 24029 2459 24087 2465
rect 25038 2456 25044 2508
rect 25096 2496 25102 2508
rect 25685 2499 25743 2505
rect 25685 2496 25697 2499
rect 25096 2468 25697 2496
rect 25096 2456 25102 2468
rect 25685 2465 25697 2468
rect 25731 2465 25743 2499
rect 25685 2459 25743 2465
rect 26142 2456 26148 2508
rect 26200 2496 26206 2508
rect 26421 2499 26479 2505
rect 26421 2496 26433 2499
rect 26200 2468 26433 2496
rect 26200 2456 26206 2468
rect 26421 2465 26433 2468
rect 26467 2465 26479 2499
rect 26421 2459 26479 2465
rect 27157 2499 27215 2505
rect 27157 2465 27169 2499
rect 27203 2496 27215 2499
rect 27246 2496 27252 2508
rect 27203 2468 27252 2496
rect 27203 2465 27215 2468
rect 27157 2459 27215 2465
rect 27246 2456 27252 2468
rect 27304 2456 27310 2508
rect 28350 2456 28356 2508
rect 28408 2496 28414 2508
rect 28445 2499 28503 2505
rect 28445 2496 28457 2499
rect 28408 2468 28457 2496
rect 28408 2456 28414 2468
rect 28445 2465 28457 2468
rect 28491 2465 28503 2499
rect 28445 2459 28503 2465
rect 29454 2456 29460 2508
rect 29512 2496 29518 2508
rect 29549 2499 29607 2505
rect 29549 2496 29561 2499
rect 29512 2468 29561 2496
rect 29512 2456 29518 2468
rect 29549 2465 29561 2468
rect 29595 2465 29607 2499
rect 29549 2459 29607 2465
rect 30558 2456 30564 2508
rect 30616 2496 30622 2508
rect 31021 2499 31079 2505
rect 31021 2496 31033 2499
rect 30616 2468 31033 2496
rect 30616 2456 30622 2468
rect 31021 2465 31033 2468
rect 31067 2465 31079 2499
rect 31021 2459 31079 2465
rect 31662 2456 31668 2508
rect 31720 2496 31726 2508
rect 31757 2499 31815 2505
rect 31757 2496 31769 2499
rect 31720 2468 31769 2496
rect 31720 2456 31726 2468
rect 31757 2465 31769 2468
rect 31803 2465 31815 2499
rect 32490 2496 32496 2508
rect 32451 2468 32496 2496
rect 31757 2459 31815 2465
rect 32490 2456 32496 2468
rect 32548 2456 32554 2508
rect 32766 2456 32772 2508
rect 32824 2496 32830 2508
rect 33689 2499 33747 2505
rect 33689 2496 33701 2499
rect 32824 2468 33701 2496
rect 32824 2456 32830 2468
rect 33689 2465 33701 2468
rect 33735 2465 33747 2499
rect 33689 2459 33747 2465
rect 33870 2456 33876 2508
rect 33928 2496 33934 2508
rect 34425 2499 34483 2505
rect 34425 2496 34437 2499
rect 33928 2468 34437 2496
rect 33928 2456 33934 2468
rect 34425 2465 34437 2468
rect 34471 2465 34483 2499
rect 34425 2459 34483 2465
rect 35161 2499 35219 2505
rect 35161 2465 35173 2499
rect 35207 2496 35219 2499
rect 35250 2496 35256 2508
rect 35207 2468 35256 2496
rect 35207 2465 35219 2468
rect 35161 2459 35219 2465
rect 35250 2456 35256 2468
rect 35308 2456 35314 2508
rect 36078 2456 36084 2508
rect 36136 2496 36142 2508
rect 36357 2499 36415 2505
rect 36357 2496 36369 2499
rect 36136 2468 36369 2496
rect 36136 2456 36142 2468
rect 36357 2465 36369 2468
rect 36403 2465 36415 2499
rect 36357 2459 36415 2465
rect 37182 2456 37188 2508
rect 37240 2496 37246 2508
rect 37277 2499 37335 2505
rect 37277 2496 37289 2499
rect 37240 2468 37289 2496
rect 37240 2456 37246 2468
rect 37277 2465 37289 2468
rect 37323 2465 37335 2499
rect 37277 2459 37335 2465
rect 38286 2456 38292 2508
rect 38344 2496 38350 2508
rect 39025 2499 39083 2505
rect 39025 2496 39037 2499
rect 38344 2468 39037 2496
rect 38344 2456 38350 2468
rect 39025 2465 39037 2468
rect 39071 2465 39083 2499
rect 39025 2459 39083 2465
rect 39942 2456 39948 2508
rect 40000 2496 40006 2508
rect 41693 2499 41751 2505
rect 41693 2496 41705 2499
rect 40000 2468 41705 2496
rect 40000 2456 40006 2468
rect 41693 2465 41705 2468
rect 41739 2465 41751 2499
rect 41693 2459 41751 2465
rect 41782 2456 41788 2508
rect 41840 2496 41846 2508
rect 42797 2499 42855 2505
rect 42797 2496 42809 2499
rect 41840 2468 42809 2496
rect 41840 2456 41846 2468
rect 42797 2465 42809 2468
rect 42843 2465 42855 2499
rect 42904 2496 42932 2536
rect 45094 2524 45100 2536
rect 45152 2524 45158 2576
rect 45186 2524 45192 2576
rect 45244 2564 45250 2576
rect 45833 2567 45891 2573
rect 45833 2564 45845 2567
rect 45244 2536 45845 2564
rect 45244 2524 45250 2536
rect 45833 2533 45845 2536
rect 45879 2533 45891 2567
rect 47210 2564 47216 2576
rect 47171 2536 47216 2564
rect 45833 2527 45891 2533
rect 47210 2524 47216 2536
rect 47268 2524 47274 2576
rect 49786 2524 49792 2576
rect 49844 2564 49850 2576
rect 50525 2567 50583 2573
rect 50525 2564 50537 2567
rect 49844 2536 50537 2564
rect 49844 2524 49850 2536
rect 50525 2533 50537 2536
rect 50571 2533 50583 2567
rect 50525 2527 50583 2533
rect 50982 2524 50988 2576
rect 51040 2564 51046 2576
rect 52365 2567 52423 2573
rect 52365 2564 52377 2567
rect 51040 2536 52377 2564
rect 51040 2524 51046 2536
rect 52365 2533 52377 2536
rect 52411 2533 52423 2567
rect 52365 2527 52423 2533
rect 52822 2524 52828 2576
rect 52880 2564 52886 2576
rect 53837 2567 53895 2573
rect 53837 2564 53849 2567
rect 52880 2536 53849 2564
rect 52880 2524 52886 2536
rect 53837 2533 53849 2536
rect 53883 2533 53895 2567
rect 53837 2527 53895 2533
rect 54018 2524 54024 2576
rect 54076 2564 54082 2576
rect 55033 2567 55091 2573
rect 55033 2564 55045 2567
rect 54076 2536 55045 2564
rect 54076 2524 54082 2536
rect 55033 2533 55045 2536
rect 55079 2533 55091 2567
rect 61286 2564 61292 2576
rect 55033 2527 55091 2533
rect 55186 2536 61292 2564
rect 44361 2499 44419 2505
rect 44361 2496 44373 2499
rect 42904 2468 44373 2496
rect 42797 2459 42855 2465
rect 44361 2465 44373 2468
rect 44407 2465 44419 2499
rect 44361 2459 44419 2465
rect 44450 2456 44456 2508
rect 44508 2496 44514 2508
rect 48314 2496 48320 2508
rect 44508 2468 47164 2496
rect 48275 2468 48320 2496
rect 44508 2456 44514 2468
rect 33778 2428 33784 2440
rect 21652 2400 33784 2428
rect 33778 2388 33784 2400
rect 33836 2388 33842 2440
rect 47026 2428 47032 2440
rect 33888 2400 47032 2428
rect 4525 2363 4583 2369
rect 4525 2329 4537 2363
rect 4571 2360 4583 2363
rect 26602 2360 26608 2372
rect 4571 2332 26234 2360
rect 26563 2332 26608 2360
rect 4571 2329 4583 2332
rect 4525 2323 4583 2329
rect 2774 2292 2780 2304
rect 2735 2264 2780 2292
rect 2774 2252 2780 2264
rect 2832 2252 2838 2304
rect 7190 2292 7196 2304
rect 7151 2264 7196 2292
rect 7190 2252 7196 2264
rect 7248 2252 7254 2304
rect 8570 2292 8576 2304
rect 8531 2264 8576 2292
rect 8570 2252 8576 2264
rect 8628 2252 8634 2304
rect 8846 2252 8852 2304
rect 8904 2292 8910 2304
rect 11241 2295 11299 2301
rect 11241 2292 11253 2295
rect 8904 2264 11253 2292
rect 8904 2252 8910 2264
rect 11241 2261 11253 2264
rect 11287 2261 11299 2295
rect 15286 2292 15292 2304
rect 15247 2264 15292 2292
rect 11241 2255 11299 2261
rect 15286 2252 15292 2264
rect 15344 2252 15350 2304
rect 16390 2292 16396 2304
rect 16351 2264 16396 2292
rect 16390 2252 16396 2264
rect 16448 2252 16454 2304
rect 17770 2292 17776 2304
rect 17731 2264 17776 2292
rect 17770 2252 17776 2264
rect 17828 2252 17834 2304
rect 21910 2292 21916 2304
rect 21871 2264 21916 2292
rect 21910 2252 21916 2264
rect 21968 2252 21974 2304
rect 23106 2292 23112 2304
rect 23067 2264 23112 2292
rect 23106 2252 23112 2264
rect 23164 2252 23170 2304
rect 24118 2292 24124 2304
rect 24079 2264 24124 2292
rect 24118 2252 24124 2264
rect 24176 2252 24182 2304
rect 25777 2295 25835 2301
rect 25777 2261 25789 2295
rect 25823 2292 25835 2295
rect 25958 2292 25964 2304
rect 25823 2264 25964 2292
rect 25823 2261 25835 2264
rect 25777 2255 25835 2261
rect 25958 2252 25964 2264
rect 26016 2252 26022 2304
rect 26206 2292 26234 2332
rect 26602 2320 26608 2332
rect 26660 2320 26666 2372
rect 27338 2360 27344 2372
rect 27299 2332 27344 2360
rect 27338 2320 27344 2332
rect 27396 2320 27402 2372
rect 28626 2360 28632 2372
rect 28587 2332 28632 2360
rect 28626 2320 28632 2332
rect 28684 2320 28690 2372
rect 29730 2360 29736 2372
rect 29691 2332 29736 2360
rect 29730 2320 29736 2332
rect 29788 2320 29794 2372
rect 29822 2320 29828 2372
rect 29880 2360 29886 2372
rect 33888 2369 33916 2400
rect 47026 2388 47032 2400
rect 47084 2388 47090 2440
rect 47136 2428 47164 2468
rect 48314 2456 48320 2468
rect 48372 2456 48378 2508
rect 49697 2499 49755 2505
rect 49697 2465 49709 2499
rect 49743 2496 49755 2499
rect 49878 2496 49884 2508
rect 49743 2468 49884 2496
rect 49743 2465 49755 2468
rect 49697 2459 49755 2465
rect 49878 2456 49884 2468
rect 49936 2456 49942 2508
rect 51166 2496 51172 2508
rect 51127 2468 51172 2496
rect 51166 2456 51172 2468
rect 51224 2456 51230 2508
rect 53098 2496 53104 2508
rect 53059 2468 53104 2496
rect 53098 2456 53104 2468
rect 53156 2456 53162 2508
rect 55186 2496 55214 2536
rect 61286 2524 61292 2536
rect 61344 2524 61350 2576
rect 61473 2567 61531 2573
rect 61473 2533 61485 2567
rect 61519 2564 61531 2567
rect 62758 2564 62764 2576
rect 61519 2536 62764 2564
rect 61519 2533 61531 2536
rect 61473 2527 61531 2533
rect 62758 2524 62764 2536
rect 62816 2524 62822 2576
rect 63037 2567 63095 2573
rect 63037 2533 63049 2567
rect 63083 2564 63095 2567
rect 63494 2564 63500 2576
rect 63083 2536 63500 2564
rect 63083 2533 63095 2536
rect 63037 2527 63095 2533
rect 63494 2524 63500 2536
rect 63552 2524 63558 2576
rect 63773 2567 63831 2573
rect 63773 2533 63785 2567
rect 63819 2564 63831 2567
rect 65242 2564 65248 2576
rect 63819 2536 65248 2564
rect 63819 2533 63831 2536
rect 63773 2527 63831 2533
rect 65242 2524 65248 2536
rect 65300 2524 65306 2576
rect 66806 2564 66812 2576
rect 65720 2536 66812 2564
rect 56042 2496 56048 2508
rect 53208 2468 55214 2496
rect 56003 2468 56048 2496
rect 53208 2428 53236 2468
rect 56042 2456 56048 2468
rect 56100 2456 56106 2508
rect 57698 2496 57704 2508
rect 57659 2468 57704 2496
rect 57698 2456 57704 2468
rect 57756 2456 57762 2508
rect 58437 2499 58495 2505
rect 58437 2465 58449 2499
rect 58483 2496 58495 2499
rect 59078 2496 59084 2508
rect 58483 2468 59084 2496
rect 58483 2465 58495 2468
rect 58437 2459 58495 2465
rect 59078 2456 59084 2468
rect 59136 2456 59142 2508
rect 59173 2499 59231 2505
rect 59173 2465 59185 2499
rect 59219 2496 59231 2499
rect 59906 2496 59912 2508
rect 59219 2468 59912 2496
rect 59219 2465 59231 2468
rect 59173 2459 59231 2465
rect 59906 2456 59912 2468
rect 59964 2456 59970 2508
rect 60369 2499 60427 2505
rect 60369 2465 60381 2499
rect 60415 2496 60427 2499
rect 60918 2496 60924 2508
rect 60415 2468 60924 2496
rect 60415 2465 60427 2468
rect 60369 2459 60427 2465
rect 60918 2456 60924 2468
rect 60976 2456 60982 2508
rect 64509 2499 64567 2505
rect 64509 2465 64521 2499
rect 64555 2496 64567 2499
rect 65720 2496 65748 2536
rect 66806 2524 66812 2536
rect 66864 2524 66870 2576
rect 66993 2567 67051 2573
rect 66993 2533 67005 2567
rect 67039 2564 67051 2567
rect 67818 2564 67824 2576
rect 67039 2536 67824 2564
rect 67039 2533 67051 2536
rect 66993 2527 67051 2533
rect 67818 2524 67824 2536
rect 67876 2524 67882 2576
rect 68373 2567 68431 2573
rect 68373 2533 68385 2567
rect 68419 2564 68431 2567
rect 69014 2564 69020 2576
rect 68419 2536 69020 2564
rect 68419 2533 68431 2536
rect 68373 2527 68431 2533
rect 69014 2524 69020 2536
rect 69072 2524 69078 2576
rect 69201 2567 69259 2573
rect 69201 2533 69213 2567
rect 69247 2564 69259 2567
rect 70366 2564 70394 2604
rect 71130 2592 71136 2604
rect 71188 2592 71194 2644
rect 71314 2592 71320 2644
rect 71372 2632 71378 2644
rect 74537 2635 74595 2641
rect 74537 2632 74549 2635
rect 71372 2604 74549 2632
rect 71372 2592 71378 2604
rect 74537 2601 74549 2604
rect 74583 2601 74595 2635
rect 74537 2595 74595 2601
rect 77754 2592 77760 2644
rect 77812 2632 77818 2644
rect 81894 2632 81900 2644
rect 77812 2604 81900 2632
rect 77812 2592 77818 2604
rect 81894 2592 81900 2604
rect 81952 2592 81958 2644
rect 82909 2635 82967 2641
rect 82909 2601 82921 2635
rect 82955 2632 82967 2635
rect 83366 2632 83372 2644
rect 82955 2604 83372 2632
rect 82955 2601 82967 2604
rect 82909 2595 82967 2601
rect 83366 2592 83372 2604
rect 83424 2592 83430 2644
rect 84102 2632 84108 2644
rect 83568 2604 84108 2632
rect 69247 2536 70394 2564
rect 71869 2567 71927 2573
rect 69247 2533 69259 2536
rect 69201 2527 69259 2533
rect 71869 2533 71881 2567
rect 71915 2564 71927 2567
rect 73430 2564 73436 2576
rect 71915 2536 73436 2564
rect 71915 2533 71927 2536
rect 71869 2527 71927 2533
rect 73430 2524 73436 2536
rect 73488 2524 73494 2576
rect 73706 2564 73712 2576
rect 73667 2536 73712 2564
rect 73706 2524 73712 2536
rect 73764 2524 73770 2576
rect 73798 2524 73804 2576
rect 73856 2564 73862 2576
rect 74445 2567 74503 2573
rect 74445 2564 74457 2567
rect 73856 2536 74457 2564
rect 73856 2524 73862 2536
rect 74445 2533 74457 2536
rect 74491 2533 74503 2567
rect 75178 2564 75184 2576
rect 75139 2536 75184 2564
rect 74445 2527 74503 2533
rect 75178 2524 75184 2536
rect 75236 2524 75242 2576
rect 76561 2567 76619 2573
rect 76561 2533 76573 2567
rect 76607 2564 76619 2567
rect 76837 2567 76895 2573
rect 76837 2564 76849 2567
rect 76607 2536 76849 2564
rect 76607 2533 76619 2536
rect 76561 2527 76619 2533
rect 76837 2533 76849 2536
rect 76883 2564 76895 2567
rect 77110 2564 77116 2576
rect 76883 2536 77116 2564
rect 76883 2533 76895 2536
rect 76837 2527 76895 2533
rect 77110 2524 77116 2536
rect 77168 2524 77174 2576
rect 77570 2524 77576 2576
rect 77628 2564 77634 2576
rect 79045 2567 79103 2573
rect 79045 2564 79057 2567
rect 77628 2536 79057 2564
rect 77628 2524 77634 2536
rect 79045 2533 79057 2536
rect 79091 2533 79103 2567
rect 79045 2527 79103 2533
rect 80057 2567 80115 2573
rect 80057 2533 80069 2567
rect 80103 2564 80115 2567
rect 80333 2567 80391 2573
rect 80333 2564 80345 2567
rect 80103 2536 80345 2564
rect 80103 2533 80115 2536
rect 80057 2527 80115 2533
rect 80333 2533 80345 2536
rect 80379 2564 80391 2567
rect 80606 2564 80612 2576
rect 80379 2536 80612 2564
rect 80379 2533 80391 2536
rect 80333 2527 80391 2533
rect 80606 2524 80612 2536
rect 80664 2524 80670 2576
rect 81802 2524 81808 2576
rect 81860 2564 81866 2576
rect 83568 2564 83596 2604
rect 84102 2592 84108 2604
rect 84160 2592 84166 2644
rect 84286 2632 84292 2644
rect 84247 2604 84292 2632
rect 84286 2592 84292 2604
rect 84344 2592 84350 2644
rect 84378 2592 84384 2644
rect 84436 2632 84442 2644
rect 85301 2635 85359 2641
rect 85301 2632 85313 2635
rect 84436 2604 85313 2632
rect 84436 2592 84442 2604
rect 85301 2601 85313 2604
rect 85347 2601 85359 2635
rect 85301 2595 85359 2601
rect 85482 2592 85488 2644
rect 85540 2632 85546 2644
rect 85540 2604 86080 2632
rect 85540 2592 85546 2604
rect 81860 2536 83596 2564
rect 81860 2524 81866 2536
rect 83642 2524 83648 2576
rect 83700 2564 83706 2576
rect 83700 2536 85620 2564
rect 83700 2524 83706 2536
rect 64555 2468 65748 2496
rect 65889 2499 65947 2505
rect 64555 2465 64567 2468
rect 64509 2459 64567 2465
rect 65889 2465 65901 2499
rect 65935 2496 65947 2499
rect 67910 2496 67916 2508
rect 65935 2468 67916 2496
rect 65935 2465 65947 2468
rect 65889 2459 65947 2465
rect 67910 2456 67916 2468
rect 67968 2456 67974 2508
rect 68002 2456 68008 2508
rect 68060 2496 68066 2508
rect 69845 2499 69903 2505
rect 69845 2496 69857 2499
rect 68060 2468 69857 2496
rect 68060 2456 68066 2468
rect 69845 2465 69857 2468
rect 69891 2465 69903 2499
rect 69845 2459 69903 2465
rect 69934 2456 69940 2508
rect 69992 2496 69998 2508
rect 72513 2499 72571 2505
rect 72513 2496 72525 2499
rect 69992 2468 72525 2496
rect 69992 2456 69998 2468
rect 72513 2465 72525 2468
rect 72559 2465 72571 2499
rect 72513 2459 72571 2465
rect 75822 2456 75828 2508
rect 75880 2496 75886 2508
rect 77757 2499 77815 2505
rect 77757 2496 77769 2499
rect 75880 2468 77769 2496
rect 75880 2456 75886 2468
rect 77757 2465 77769 2468
rect 77803 2465 77815 2499
rect 77757 2459 77815 2465
rect 80238 2456 80244 2508
rect 80296 2496 80302 2508
rect 82170 2496 82176 2508
rect 80296 2468 82032 2496
rect 82131 2468 82176 2496
rect 80296 2456 80302 2468
rect 47136 2400 53236 2428
rect 53282 2388 53288 2440
rect 53340 2428 53346 2440
rect 77205 2431 77263 2437
rect 53340 2400 75500 2428
rect 53340 2388 53346 2400
rect 32677 2363 32735 2369
rect 32677 2360 32689 2363
rect 29880 2332 32689 2360
rect 29880 2320 29886 2332
rect 32677 2329 32689 2332
rect 32723 2329 32735 2363
rect 32677 2323 32735 2329
rect 33873 2363 33931 2369
rect 33873 2329 33885 2363
rect 33919 2329 33931 2363
rect 33873 2323 33931 2329
rect 35345 2363 35403 2369
rect 35345 2329 35357 2363
rect 35391 2360 35403 2363
rect 35391 2332 59216 2360
rect 35391 2329 35403 2332
rect 35345 2323 35403 2329
rect 30834 2292 30840 2304
rect 26206 2264 30840 2292
rect 30834 2252 30840 2264
rect 30892 2252 30898 2304
rect 31110 2292 31116 2304
rect 31071 2264 31116 2292
rect 31110 2252 31116 2264
rect 31168 2252 31174 2304
rect 34514 2292 34520 2304
rect 34475 2264 34520 2292
rect 34514 2252 34520 2264
rect 34572 2252 34578 2304
rect 36449 2295 36507 2301
rect 36449 2261 36461 2295
rect 36495 2292 36507 2295
rect 37274 2292 37280 2304
rect 36495 2264 37280 2292
rect 36495 2261 36507 2264
rect 36449 2255 36507 2261
rect 37274 2252 37280 2264
rect 37332 2252 37338 2304
rect 37366 2252 37372 2304
rect 37424 2292 37430 2304
rect 38838 2292 38844 2304
rect 37424 2264 38844 2292
rect 37424 2252 37430 2264
rect 38838 2252 38844 2264
rect 38896 2252 38902 2304
rect 39114 2292 39120 2304
rect 39075 2264 39120 2292
rect 39114 2252 39120 2264
rect 39172 2252 39178 2304
rect 39390 2252 39396 2304
rect 39448 2292 39454 2304
rect 39853 2295 39911 2301
rect 39853 2292 39865 2295
rect 39448 2264 39865 2292
rect 39448 2252 39454 2264
rect 39853 2261 39865 2264
rect 39899 2261 39911 2295
rect 39853 2255 39911 2261
rect 40494 2252 40500 2304
rect 40552 2292 40558 2304
rect 40589 2295 40647 2301
rect 40589 2292 40601 2295
rect 40552 2264 40601 2292
rect 40552 2252 40558 2264
rect 40589 2261 40601 2264
rect 40635 2261 40647 2295
rect 40589 2255 40647 2261
rect 41598 2252 41604 2304
rect 41656 2292 41662 2304
rect 41785 2295 41843 2301
rect 41785 2292 41797 2295
rect 41656 2264 41797 2292
rect 41656 2252 41662 2264
rect 41785 2261 41797 2264
rect 41831 2261 41843 2295
rect 41785 2255 41843 2261
rect 42702 2252 42708 2304
rect 42760 2292 42766 2304
rect 42889 2295 42947 2301
rect 42889 2292 42901 2295
rect 42760 2264 42901 2292
rect 42760 2252 42766 2264
rect 42889 2261 42901 2264
rect 42935 2261 42947 2295
rect 42889 2255 42947 2261
rect 43806 2252 43812 2304
rect 43864 2292 43870 2304
rect 44453 2295 44511 2301
rect 44453 2292 44465 2295
rect 43864 2264 44465 2292
rect 43864 2252 43870 2264
rect 44453 2261 44465 2264
rect 44499 2261 44511 2295
rect 44453 2255 44511 2261
rect 44910 2252 44916 2304
rect 44968 2292 44974 2304
rect 45189 2295 45247 2301
rect 45189 2292 45201 2295
rect 44968 2264 45201 2292
rect 44968 2252 44974 2264
rect 45189 2261 45201 2264
rect 45235 2261 45247 2295
rect 45189 2255 45247 2261
rect 45925 2295 45983 2301
rect 45925 2261 45937 2295
rect 45971 2292 45983 2295
rect 46014 2292 46020 2304
rect 45971 2264 46020 2292
rect 45971 2261 45983 2264
rect 45925 2255 45983 2261
rect 46014 2252 46020 2264
rect 46072 2252 46078 2304
rect 47118 2252 47124 2304
rect 47176 2292 47182 2304
rect 47305 2295 47363 2301
rect 47305 2292 47317 2295
rect 47176 2264 47317 2292
rect 47176 2252 47182 2264
rect 47305 2261 47317 2264
rect 47351 2261 47363 2295
rect 47305 2255 47363 2261
rect 48222 2252 48228 2304
rect 48280 2292 48286 2304
rect 48409 2295 48467 2301
rect 48409 2292 48421 2295
rect 48280 2264 48421 2292
rect 48280 2252 48286 2264
rect 48409 2261 48421 2264
rect 48455 2261 48467 2295
rect 48409 2255 48467 2261
rect 49326 2252 49332 2304
rect 49384 2292 49390 2304
rect 49789 2295 49847 2301
rect 49789 2292 49801 2295
rect 49384 2264 49801 2292
rect 49384 2252 49390 2264
rect 49789 2261 49801 2264
rect 49835 2261 49847 2295
rect 49789 2255 49847 2261
rect 50430 2252 50436 2304
rect 50488 2292 50494 2304
rect 50617 2295 50675 2301
rect 50617 2292 50629 2295
rect 50488 2264 50629 2292
rect 50488 2252 50494 2264
rect 50617 2261 50629 2264
rect 50663 2261 50675 2295
rect 50617 2255 50675 2261
rect 51534 2252 51540 2304
rect 51592 2292 51598 2304
rect 52457 2295 52515 2301
rect 52457 2292 52469 2295
rect 51592 2264 52469 2292
rect 51592 2252 51598 2264
rect 52457 2261 52469 2264
rect 52503 2261 52515 2295
rect 52457 2255 52515 2261
rect 52638 2252 52644 2304
rect 52696 2292 52702 2304
rect 53193 2295 53251 2301
rect 53193 2292 53205 2295
rect 52696 2264 53205 2292
rect 52696 2252 52702 2264
rect 53193 2261 53205 2264
rect 53239 2261 53251 2295
rect 53193 2255 53251 2261
rect 53742 2252 53748 2304
rect 53800 2292 53806 2304
rect 53929 2295 53987 2301
rect 53929 2292 53941 2295
rect 53800 2264 53941 2292
rect 53800 2252 53806 2264
rect 53929 2261 53941 2264
rect 53975 2261 53987 2295
rect 53929 2255 53987 2261
rect 54846 2252 54852 2304
rect 54904 2292 54910 2304
rect 55125 2295 55183 2301
rect 55125 2292 55137 2295
rect 54904 2264 55137 2292
rect 54904 2252 54910 2264
rect 55125 2261 55137 2264
rect 55171 2261 55183 2295
rect 55125 2255 55183 2261
rect 55950 2252 55956 2304
rect 56008 2292 56014 2304
rect 56137 2295 56195 2301
rect 56137 2292 56149 2295
rect 56008 2264 56149 2292
rect 56008 2252 56014 2264
rect 56137 2261 56149 2264
rect 56183 2261 56195 2295
rect 56137 2255 56195 2261
rect 57054 2252 57060 2304
rect 57112 2292 57118 2304
rect 57793 2295 57851 2301
rect 57793 2292 57805 2295
rect 57112 2264 57805 2292
rect 57112 2252 57118 2264
rect 57793 2261 57805 2264
rect 57839 2261 57851 2295
rect 57793 2255 57851 2261
rect 58158 2252 58164 2304
rect 58216 2292 58222 2304
rect 58529 2295 58587 2301
rect 58529 2292 58541 2295
rect 58216 2264 58541 2292
rect 58216 2252 58222 2264
rect 58529 2261 58541 2264
rect 58575 2261 58587 2295
rect 59188 2292 59216 2332
rect 59262 2320 59268 2372
rect 59320 2360 59326 2372
rect 59357 2363 59415 2369
rect 59357 2360 59369 2363
rect 59320 2332 59369 2360
rect 59320 2320 59326 2332
rect 59357 2329 59369 2332
rect 59403 2329 59415 2363
rect 64230 2360 64236 2372
rect 59357 2323 59415 2329
rect 59464 2332 64236 2360
rect 59464 2292 59492 2332
rect 64230 2320 64236 2332
rect 64288 2320 64294 2372
rect 64690 2360 64696 2372
rect 64651 2332 64696 2360
rect 64690 2320 64696 2332
rect 64748 2320 64754 2372
rect 71406 2320 71412 2372
rect 71464 2360 71470 2372
rect 71501 2363 71559 2369
rect 71501 2360 71513 2363
rect 71464 2332 71513 2360
rect 71464 2320 71470 2332
rect 71501 2329 71513 2332
rect 71547 2329 71559 2363
rect 73893 2363 73951 2369
rect 73893 2360 73905 2363
rect 71501 2323 71559 2329
rect 71700 2332 73905 2360
rect 59188 2264 59492 2292
rect 58529 2255 58587 2261
rect 60274 2252 60280 2304
rect 60332 2292 60338 2304
rect 60461 2295 60519 2301
rect 60461 2292 60473 2295
rect 60332 2264 60473 2292
rect 60332 2252 60338 2264
rect 60461 2261 60473 2264
rect 60507 2261 60519 2295
rect 60461 2255 60519 2261
rect 61378 2252 61384 2304
rect 61436 2292 61442 2304
rect 61565 2295 61623 2301
rect 61565 2292 61577 2295
rect 61436 2264 61577 2292
rect 61436 2252 61442 2264
rect 61565 2261 61577 2264
rect 61611 2261 61623 2295
rect 61565 2255 61623 2261
rect 62482 2252 62488 2304
rect 62540 2292 62546 2304
rect 63129 2295 63187 2301
rect 63129 2292 63141 2295
rect 62540 2264 63141 2292
rect 62540 2252 62546 2264
rect 63129 2261 63141 2264
rect 63175 2261 63187 2295
rect 63129 2255 63187 2261
rect 63586 2252 63592 2304
rect 63644 2292 63650 2304
rect 63865 2295 63923 2301
rect 63865 2292 63877 2295
rect 63644 2264 63877 2292
rect 63644 2252 63650 2264
rect 63865 2261 63877 2264
rect 63911 2261 63923 2295
rect 65978 2292 65984 2304
rect 65939 2264 65984 2292
rect 63865 2255 63923 2261
rect 65978 2252 65984 2264
rect 66036 2252 66042 2304
rect 66898 2252 66904 2304
rect 66956 2292 66962 2304
rect 67085 2295 67143 2301
rect 67085 2292 67097 2295
rect 66956 2264 67097 2292
rect 66956 2252 66962 2264
rect 67085 2261 67097 2264
rect 67131 2261 67143 2295
rect 67085 2255 67143 2261
rect 68002 2252 68008 2304
rect 68060 2292 68066 2304
rect 68465 2295 68523 2301
rect 68465 2292 68477 2295
rect 68060 2264 68477 2292
rect 68060 2252 68066 2264
rect 68465 2261 68477 2264
rect 68511 2261 68523 2295
rect 68465 2255 68523 2261
rect 69106 2252 69112 2304
rect 69164 2292 69170 2304
rect 69293 2295 69351 2301
rect 69293 2292 69305 2295
rect 69164 2264 69305 2292
rect 69164 2252 69170 2264
rect 69293 2261 69305 2264
rect 69339 2261 69351 2295
rect 69293 2255 69351 2261
rect 70210 2252 70216 2304
rect 70268 2292 70274 2304
rect 71700 2292 71728 2332
rect 73893 2329 73905 2332
rect 73939 2329 73951 2363
rect 75365 2363 75423 2369
rect 75365 2360 75377 2363
rect 73893 2323 73951 2329
rect 74000 2332 75377 2360
rect 71866 2292 71872 2304
rect 70268 2264 71728 2292
rect 71827 2264 71872 2292
rect 70268 2252 70274 2264
rect 71866 2252 71872 2264
rect 71924 2252 71930 2304
rect 71958 2252 71964 2304
rect 72016 2292 72022 2304
rect 72053 2295 72111 2301
rect 72053 2292 72065 2295
rect 72016 2264 72065 2292
rect 72016 2252 72022 2264
rect 72053 2261 72065 2264
rect 72099 2261 72111 2295
rect 72053 2255 72111 2261
rect 72418 2252 72424 2304
rect 72476 2292 72482 2304
rect 74000 2292 74028 2332
rect 75365 2329 75377 2332
rect 75411 2329 75423 2363
rect 75365 2323 75423 2329
rect 72476 2264 74028 2292
rect 75472 2292 75500 2400
rect 77205 2397 77217 2431
rect 77251 2428 77263 2431
rect 81802 2428 81808 2440
rect 77251 2400 81808 2428
rect 77251 2397 77263 2400
rect 77205 2391 77263 2397
rect 81802 2388 81808 2400
rect 81860 2388 81866 2440
rect 82004 2428 82032 2468
rect 82170 2456 82176 2468
rect 82228 2456 82234 2508
rect 82262 2456 82268 2508
rect 82320 2496 82326 2508
rect 82357 2499 82415 2505
rect 82357 2496 82369 2499
rect 82320 2468 82369 2496
rect 82320 2456 82326 2468
rect 82357 2465 82369 2468
rect 82403 2465 82415 2499
rect 82538 2496 82544 2508
rect 82499 2468 82544 2496
rect 82357 2459 82415 2465
rect 82538 2456 82544 2468
rect 82596 2456 82602 2508
rect 82725 2499 82783 2505
rect 82725 2465 82737 2499
rect 82771 2496 82783 2499
rect 82814 2496 82820 2508
rect 82771 2468 82820 2496
rect 82771 2465 82783 2468
rect 82725 2459 82783 2465
rect 82449 2431 82507 2437
rect 82449 2428 82461 2431
rect 82004 2400 82461 2428
rect 82449 2397 82461 2400
rect 82495 2428 82507 2431
rect 82630 2428 82636 2440
rect 82495 2400 82636 2428
rect 82495 2397 82507 2400
rect 82449 2391 82507 2397
rect 82630 2388 82636 2400
rect 82688 2388 82694 2440
rect 76282 2320 76288 2372
rect 76340 2360 76346 2372
rect 76340 2332 76880 2360
rect 76340 2320 76346 2332
rect 76852 2301 76880 2332
rect 77018 2320 77024 2372
rect 77076 2360 77082 2372
rect 79229 2363 79287 2369
rect 79229 2360 79241 2363
rect 77076 2332 79241 2360
rect 77076 2320 77082 2332
rect 79229 2329 79241 2332
rect 79275 2329 79287 2363
rect 79229 2323 79287 2329
rect 80701 2363 80759 2369
rect 80701 2329 80713 2363
rect 80747 2360 80759 2363
rect 82740 2360 82768 2459
rect 82814 2456 82820 2468
rect 82872 2456 82878 2508
rect 84473 2499 84531 2505
rect 84473 2465 84485 2499
rect 84519 2465 84531 2499
rect 84473 2459 84531 2465
rect 84488 2428 84516 2459
rect 84562 2456 84568 2508
rect 84620 2496 84626 2508
rect 84838 2496 84844 2508
rect 84620 2468 84665 2496
rect 84799 2468 84844 2496
rect 84620 2456 84626 2468
rect 84838 2456 84844 2468
rect 84896 2456 84902 2508
rect 85482 2496 85488 2508
rect 85443 2468 85488 2496
rect 85482 2456 85488 2468
rect 85540 2456 85546 2508
rect 85592 2505 85620 2536
rect 85577 2499 85635 2505
rect 85577 2465 85589 2499
rect 85623 2465 85635 2499
rect 85850 2496 85856 2508
rect 85811 2468 85856 2496
rect 85577 2459 85635 2465
rect 85850 2456 85856 2468
rect 85908 2456 85914 2508
rect 86052 2496 86080 2604
rect 86126 2592 86132 2644
rect 86184 2632 86190 2644
rect 89806 2632 89812 2644
rect 86184 2604 89714 2632
rect 89767 2604 89812 2632
rect 86184 2592 86190 2604
rect 86586 2524 86592 2576
rect 86644 2564 86650 2576
rect 86770 2564 86776 2576
rect 86644 2536 86776 2564
rect 86644 2524 86650 2536
rect 86770 2524 86776 2536
rect 86828 2524 86834 2576
rect 86865 2567 86923 2573
rect 86865 2533 86877 2567
rect 86911 2564 86923 2567
rect 87141 2567 87199 2573
rect 87141 2564 87153 2567
rect 86911 2536 87153 2564
rect 86911 2533 86923 2536
rect 86865 2527 86923 2533
rect 87141 2533 87153 2536
rect 87187 2564 87199 2567
rect 87322 2564 87328 2576
rect 87187 2536 87328 2564
rect 87187 2533 87199 2536
rect 87141 2527 87199 2533
rect 87322 2524 87328 2536
rect 87380 2524 87386 2576
rect 87877 2567 87935 2573
rect 87877 2533 87889 2567
rect 87923 2564 87935 2567
rect 88150 2564 88156 2576
rect 87923 2536 88156 2564
rect 87923 2533 87935 2536
rect 87877 2527 87935 2533
rect 88150 2524 88156 2536
rect 88208 2524 88214 2576
rect 89686 2564 89714 2604
rect 89806 2592 89812 2604
rect 89864 2592 89870 2644
rect 93394 2592 93400 2644
rect 93452 2632 93458 2644
rect 95881 2635 95939 2641
rect 95881 2632 95893 2635
rect 93452 2604 95893 2632
rect 93452 2592 93458 2604
rect 95881 2601 95893 2604
rect 95927 2601 95939 2635
rect 106458 2632 106464 2644
rect 95881 2595 95939 2601
rect 103486 2604 106464 2632
rect 90453 2567 90511 2573
rect 90453 2564 90465 2567
rect 88260 2536 89484 2564
rect 89686 2536 90465 2564
rect 87230 2496 87236 2508
rect 86052 2468 87236 2496
rect 87230 2456 87236 2468
rect 87288 2456 87294 2508
rect 87414 2456 87420 2508
rect 87472 2496 87478 2508
rect 88058 2496 88064 2508
rect 87472 2468 88064 2496
rect 87472 2456 87478 2468
rect 88058 2456 88064 2468
rect 88116 2456 88122 2508
rect 84488 2400 85620 2428
rect 80747 2332 82768 2360
rect 80747 2329 80759 2332
rect 80701 2323 80759 2329
rect 82998 2320 83004 2372
rect 83056 2360 83062 2372
rect 85592 2360 85620 2400
rect 86218 2388 86224 2440
rect 86276 2428 86282 2440
rect 87509 2431 87567 2437
rect 86276 2400 87460 2428
rect 86276 2388 86282 2400
rect 87432 2360 87460 2400
rect 87509 2397 87521 2431
rect 87555 2428 87567 2431
rect 87690 2428 87696 2440
rect 87555 2400 87696 2428
rect 87555 2397 87567 2400
rect 87509 2391 87567 2397
rect 87690 2388 87696 2400
rect 87748 2388 87754 2440
rect 87874 2388 87880 2440
rect 87932 2428 87938 2440
rect 88260 2428 88288 2536
rect 88518 2496 88524 2508
rect 88479 2468 88524 2496
rect 88518 2456 88524 2468
rect 88576 2496 88582 2508
rect 88576 2468 89208 2496
rect 88576 2456 88582 2468
rect 87932 2400 88288 2428
rect 87932 2388 87938 2400
rect 89180 2360 89208 2468
rect 89456 2428 89484 2536
rect 90453 2533 90465 2536
rect 90499 2533 90511 2567
rect 92382 2564 92388 2576
rect 92343 2536 92388 2564
rect 90453 2527 90511 2533
rect 92382 2524 92388 2536
rect 92440 2524 92446 2576
rect 93118 2564 93124 2576
rect 93079 2536 93124 2564
rect 93118 2524 93124 2536
rect 93176 2524 93182 2576
rect 93210 2524 93216 2576
rect 93268 2564 93274 2576
rect 93857 2567 93915 2573
rect 93857 2564 93869 2567
rect 93268 2536 93869 2564
rect 93268 2524 93274 2536
rect 93857 2533 93869 2536
rect 93903 2533 93915 2567
rect 93857 2527 93915 2533
rect 94406 2524 94412 2576
rect 94464 2564 94470 2576
rect 95789 2567 95847 2573
rect 95789 2564 95801 2567
rect 94464 2536 95801 2564
rect 94464 2524 94470 2536
rect 95789 2533 95801 2536
rect 95835 2533 95847 2567
rect 95789 2527 95847 2533
rect 96062 2524 96068 2576
rect 96120 2564 96126 2576
rect 96525 2567 96583 2573
rect 96525 2564 96537 2567
rect 96120 2536 96537 2564
rect 96120 2524 96126 2536
rect 96525 2533 96537 2536
rect 96571 2533 96583 2567
rect 96525 2527 96583 2533
rect 96614 2524 96620 2576
rect 96672 2564 96678 2576
rect 97721 2567 97779 2573
rect 97721 2564 97733 2567
rect 96672 2536 97733 2564
rect 96672 2524 96678 2536
rect 97721 2533 97733 2536
rect 97767 2533 97779 2567
rect 98454 2564 98460 2576
rect 98415 2536 98460 2564
rect 97721 2527 97779 2533
rect 98454 2524 98460 2536
rect 98512 2524 98518 2576
rect 98730 2524 98736 2576
rect 98788 2564 98794 2576
rect 99193 2567 99251 2573
rect 99193 2564 99205 2567
rect 98788 2536 99205 2564
rect 98788 2524 98794 2536
rect 99193 2533 99205 2536
rect 99239 2533 99251 2567
rect 99193 2527 99251 2533
rect 99926 2524 99932 2576
rect 99984 2564 99990 2576
rect 100389 2567 100447 2573
rect 100389 2564 100401 2567
rect 99984 2536 100401 2564
rect 99984 2524 99990 2536
rect 100389 2533 100401 2536
rect 100435 2533 100447 2567
rect 101122 2564 101128 2576
rect 101083 2536 101128 2564
rect 100389 2527 100447 2533
rect 101122 2524 101128 2536
rect 101180 2524 101186 2576
rect 101858 2564 101864 2576
rect 101819 2536 101864 2564
rect 101858 2524 101864 2536
rect 101916 2524 101922 2576
rect 102226 2524 102232 2576
rect 102284 2564 102290 2576
rect 103057 2567 103115 2573
rect 103057 2564 103069 2567
rect 102284 2536 103069 2564
rect 102284 2524 102290 2536
rect 103057 2533 103069 2536
rect 103103 2533 103115 2567
rect 103057 2527 103115 2533
rect 103146 2524 103152 2576
rect 103204 2564 103210 2576
rect 103486 2564 103514 2604
rect 106458 2592 106464 2604
rect 106516 2592 106522 2644
rect 107194 2592 107200 2644
rect 107252 2632 107258 2644
rect 111153 2635 111211 2641
rect 111153 2632 111165 2635
rect 107252 2604 111165 2632
rect 107252 2592 107258 2604
rect 111153 2601 111165 2604
rect 111199 2601 111211 2635
rect 111153 2595 111211 2601
rect 103204 2536 103514 2564
rect 103204 2524 103210 2536
rect 103698 2524 103704 2576
rect 103756 2564 103762 2576
rect 103793 2567 103851 2573
rect 103793 2564 103805 2567
rect 103756 2536 103805 2564
rect 103756 2524 103762 2536
rect 103793 2533 103805 2536
rect 103839 2533 103851 2567
rect 103793 2527 103851 2533
rect 104434 2524 104440 2576
rect 104492 2564 104498 2576
rect 104529 2567 104587 2573
rect 104529 2564 104541 2567
rect 104492 2536 104541 2564
rect 104492 2524 104498 2536
rect 104529 2533 104541 2536
rect 104575 2533 104587 2567
rect 104529 2527 104587 2533
rect 105538 2524 105544 2576
rect 105596 2564 105602 2576
rect 105725 2567 105783 2573
rect 105725 2564 105737 2567
rect 105596 2536 105737 2564
rect 105596 2524 105602 2536
rect 105725 2533 105737 2536
rect 105771 2533 105783 2567
rect 105725 2527 105783 2533
rect 106642 2524 106648 2576
rect 106700 2564 106706 2576
rect 106737 2567 106795 2573
rect 106737 2564 106749 2567
rect 106700 2536 106749 2564
rect 106700 2524 106706 2536
rect 106737 2533 106749 2536
rect 106783 2533 106795 2567
rect 109126 2564 109132 2576
rect 109087 2536 109132 2564
rect 106737 2527 106795 2533
rect 109126 2524 109132 2536
rect 109184 2524 109190 2576
rect 109862 2564 109868 2576
rect 109823 2536 109868 2564
rect 109862 2524 109868 2536
rect 109920 2524 109926 2576
rect 111610 2524 111616 2576
rect 111668 2564 111674 2576
rect 111797 2567 111855 2573
rect 111797 2564 111809 2567
rect 111668 2536 111809 2564
rect 111668 2524 111674 2536
rect 111797 2533 111809 2536
rect 111843 2533 111855 2567
rect 111797 2527 111855 2533
rect 112438 2524 112444 2576
rect 112496 2564 112502 2576
rect 112533 2567 112591 2573
rect 112533 2564 112545 2567
rect 112496 2536 112545 2564
rect 112496 2524 112502 2536
rect 112533 2533 112545 2536
rect 112579 2533 112591 2567
rect 112533 2527 112591 2533
rect 113174 2524 113180 2576
rect 113232 2564 113238 2576
rect 113729 2567 113787 2573
rect 113729 2564 113741 2567
rect 113232 2536 113741 2564
rect 113232 2524 113238 2536
rect 113729 2533 113741 2536
rect 113775 2533 113787 2567
rect 113729 2527 113787 2533
rect 114278 2524 114284 2576
rect 114336 2564 114342 2576
rect 114465 2567 114523 2573
rect 114465 2564 114477 2567
rect 114336 2536 114477 2564
rect 114336 2524 114342 2536
rect 114465 2533 114477 2536
rect 114511 2533 114523 2567
rect 115198 2564 115204 2576
rect 115159 2536 115204 2564
rect 114465 2527 114523 2533
rect 115198 2524 115204 2536
rect 115256 2524 115262 2576
rect 116394 2564 116400 2576
rect 116355 2536 116400 2564
rect 116394 2524 116400 2536
rect 116452 2524 116458 2576
rect 117130 2564 117136 2576
rect 117091 2536 117136 2564
rect 117130 2524 117136 2536
rect 117188 2524 117194 2576
rect 117774 2524 117780 2576
rect 117832 2564 117838 2576
rect 117869 2567 117927 2573
rect 117869 2564 117881 2567
rect 117832 2536 117881 2564
rect 117832 2524 117838 2536
rect 117869 2533 117881 2536
rect 117915 2533 117927 2567
rect 117869 2527 117927 2533
rect 118786 2524 118792 2576
rect 118844 2564 118850 2576
rect 119065 2567 119123 2573
rect 119065 2564 119077 2567
rect 118844 2536 119077 2564
rect 118844 2524 118850 2536
rect 119065 2533 119077 2536
rect 119111 2533 119123 2567
rect 119065 2527 119123 2533
rect 119890 2524 119896 2576
rect 119948 2564 119954 2576
rect 119985 2567 120043 2573
rect 119985 2564 119997 2567
rect 119948 2536 119997 2564
rect 119948 2524 119954 2536
rect 119985 2533 119997 2536
rect 120031 2533 120043 2567
rect 121730 2564 121736 2576
rect 121691 2536 121736 2564
rect 119985 2527 120043 2533
rect 121730 2524 121736 2536
rect 121788 2524 121794 2576
rect 122374 2524 122380 2576
rect 122432 2564 122438 2576
rect 122469 2567 122527 2573
rect 122469 2564 122481 2567
rect 122432 2536 122481 2564
rect 122432 2524 122438 2536
rect 122469 2533 122481 2536
rect 122515 2533 122527 2567
rect 122469 2527 122527 2533
rect 123110 2524 123116 2576
rect 123168 2564 123174 2576
rect 123205 2567 123263 2573
rect 123205 2564 123217 2567
rect 123168 2536 123217 2564
rect 123168 2524 123174 2536
rect 123205 2533 123217 2536
rect 123251 2533 123263 2567
rect 123205 2527 123263 2533
rect 124214 2524 124220 2576
rect 124272 2564 124278 2576
rect 124401 2567 124459 2573
rect 124401 2564 124413 2567
rect 124272 2536 124413 2564
rect 124272 2524 124278 2536
rect 124401 2533 124413 2536
rect 124447 2533 124459 2567
rect 124401 2527 124459 2533
rect 125318 2524 125324 2576
rect 125376 2564 125382 2576
rect 125413 2567 125471 2573
rect 125413 2564 125425 2567
rect 125376 2536 125425 2564
rect 125376 2524 125382 2536
rect 125413 2533 125425 2536
rect 125459 2533 125471 2567
rect 127066 2564 127072 2576
rect 127027 2536 127072 2564
rect 125413 2527 125471 2533
rect 127066 2524 127072 2536
rect 127124 2524 127130 2576
rect 127618 2524 127624 2576
rect 127676 2564 127682 2576
rect 127805 2567 127863 2573
rect 127805 2564 127817 2567
rect 127676 2536 127817 2564
rect 127676 2524 127682 2536
rect 127805 2533 127817 2536
rect 127851 2533 127863 2567
rect 127805 2527 127863 2533
rect 128541 2567 128599 2573
rect 128541 2533 128553 2567
rect 128587 2564 128599 2567
rect 128630 2564 128636 2576
rect 128587 2536 128636 2564
rect 128587 2533 128599 2536
rect 128541 2527 128599 2533
rect 128630 2524 128636 2536
rect 128688 2524 128694 2576
rect 129734 2524 129740 2576
rect 129792 2564 129798 2576
rect 129829 2567 129887 2573
rect 129829 2564 129841 2567
rect 129792 2536 129841 2564
rect 129792 2524 129798 2536
rect 129829 2533 129841 2536
rect 129875 2533 129887 2567
rect 129829 2527 129887 2533
rect 130838 2524 130844 2576
rect 130896 2564 130902 2576
rect 130933 2567 130991 2573
rect 130933 2564 130945 2567
rect 130896 2536 130945 2564
rect 130896 2524 130902 2536
rect 130933 2533 130945 2536
rect 130979 2533 130991 2567
rect 130933 2527 130991 2533
rect 131942 2524 131948 2576
rect 132000 2564 132006 2576
rect 132405 2567 132463 2573
rect 132405 2564 132417 2567
rect 132000 2536 132417 2564
rect 132000 2524 132006 2536
rect 132405 2533 132417 2536
rect 132451 2533 132463 2567
rect 132405 2527 132463 2533
rect 133046 2524 133052 2576
rect 133104 2564 133110 2576
rect 133141 2567 133199 2573
rect 133141 2564 133153 2567
rect 133104 2536 133153 2564
rect 133104 2524 133110 2536
rect 133141 2533 133153 2536
rect 133187 2533 133199 2567
rect 133141 2527 133199 2533
rect 134150 2524 134156 2576
rect 134208 2564 134214 2576
rect 135073 2567 135131 2573
rect 135073 2564 135085 2567
rect 134208 2536 135085 2564
rect 134208 2524 134214 2536
rect 135073 2533 135085 2536
rect 135119 2533 135131 2567
rect 135073 2527 135131 2533
rect 135254 2524 135260 2576
rect 135312 2564 135318 2576
rect 135809 2567 135867 2573
rect 135809 2564 135821 2567
rect 135312 2536 135821 2564
rect 135312 2524 135318 2536
rect 135809 2533 135821 2536
rect 135855 2533 135867 2567
rect 135809 2527 135867 2533
rect 136358 2524 136364 2576
rect 136416 2564 136422 2576
rect 136545 2567 136603 2573
rect 136545 2564 136557 2567
rect 136416 2536 136557 2564
rect 136416 2524 136422 2536
rect 136545 2533 136557 2536
rect 136591 2533 136603 2567
rect 136545 2527 136603 2533
rect 137741 2567 137799 2573
rect 137741 2533 137753 2567
rect 137787 2564 137799 2567
rect 138106 2564 138112 2576
rect 137787 2536 138112 2564
rect 137787 2533 137799 2536
rect 137741 2527 137799 2533
rect 138106 2524 138112 2536
rect 138164 2524 138170 2576
rect 138661 2567 138719 2573
rect 138661 2533 138673 2567
rect 138707 2564 138719 2567
rect 138750 2564 138756 2576
rect 138707 2536 138756 2564
rect 138707 2533 138719 2536
rect 138661 2527 138719 2533
rect 138750 2524 138756 2536
rect 138808 2524 138814 2576
rect 139670 2524 139676 2576
rect 139728 2564 139734 2576
rect 140409 2567 140467 2573
rect 140409 2564 140421 2567
rect 139728 2536 140421 2564
rect 139728 2524 139734 2536
rect 140409 2533 140421 2536
rect 140455 2533 140467 2567
rect 140409 2527 140467 2533
rect 140774 2524 140780 2576
rect 140832 2564 140838 2576
rect 141145 2567 141203 2573
rect 141145 2564 141157 2567
rect 140832 2536 141157 2564
rect 140832 2524 140838 2536
rect 141145 2533 141157 2536
rect 141191 2533 141203 2567
rect 141878 2564 141884 2576
rect 141839 2536 141884 2564
rect 141145 2527 141203 2533
rect 141878 2524 141884 2536
rect 141936 2524 141942 2576
rect 143077 2567 143135 2573
rect 143077 2533 143089 2567
rect 143123 2564 143135 2567
rect 143350 2564 143356 2576
rect 143123 2536 143356 2564
rect 143123 2533 143135 2536
rect 143077 2527 143135 2533
rect 143350 2524 143356 2536
rect 143408 2524 143414 2576
rect 144086 2524 144092 2576
rect 144144 2564 144150 2576
rect 144181 2567 144239 2573
rect 144181 2564 144193 2567
rect 144144 2536 144193 2564
rect 144144 2524 144150 2536
rect 144181 2533 144193 2536
rect 144227 2533 144239 2567
rect 144181 2527 144239 2533
rect 145190 2524 145196 2576
rect 145248 2564 145254 2576
rect 145745 2567 145803 2573
rect 145745 2564 145757 2567
rect 145248 2536 145757 2564
rect 145248 2524 145254 2536
rect 145745 2533 145757 2536
rect 145791 2533 145803 2567
rect 145745 2527 145803 2533
rect 146294 2524 146300 2576
rect 146352 2564 146358 2576
rect 146481 2567 146539 2573
rect 146481 2564 146493 2567
rect 146352 2536 146493 2564
rect 146352 2524 146358 2536
rect 146481 2533 146493 2536
rect 146527 2533 146539 2567
rect 146481 2527 146539 2533
rect 147217 2567 147275 2573
rect 147217 2533 147229 2567
rect 147263 2564 147275 2567
rect 147398 2564 147404 2576
rect 147263 2536 147404 2564
rect 147263 2533 147275 2536
rect 147217 2527 147275 2533
rect 147398 2524 147404 2536
rect 147456 2524 147462 2576
rect 148594 2564 148600 2576
rect 148555 2536 148600 2564
rect 148594 2524 148600 2536
rect 148652 2524 148658 2576
rect 149606 2524 149612 2576
rect 149664 2564 149670 2576
rect 149701 2567 149759 2573
rect 149701 2564 149713 2567
rect 149664 2536 149713 2564
rect 149664 2524 149670 2536
rect 149701 2533 149713 2536
rect 149747 2533 149759 2567
rect 149701 2527 149759 2533
rect 150710 2524 150716 2576
rect 150768 2564 150774 2576
rect 151081 2567 151139 2573
rect 151081 2564 151093 2567
rect 150768 2536 151093 2564
rect 150768 2524 150774 2536
rect 151081 2533 151093 2536
rect 151127 2533 151139 2567
rect 151081 2527 151139 2533
rect 151814 2524 151820 2576
rect 151872 2564 151878 2576
rect 151909 2567 151967 2573
rect 151909 2564 151921 2567
rect 151872 2536 151921 2564
rect 151872 2524 151878 2536
rect 151909 2533 151921 2536
rect 151955 2533 151967 2567
rect 153746 2564 153752 2576
rect 153707 2536 153752 2564
rect 151909 2527 151967 2533
rect 153746 2524 153752 2536
rect 153804 2524 153810 2576
rect 154022 2524 154028 2576
rect 154080 2564 154086 2576
rect 154485 2567 154543 2573
rect 154485 2564 154497 2567
rect 154080 2536 154497 2564
rect 154080 2524 154086 2536
rect 154485 2533 154497 2536
rect 154531 2533 154543 2567
rect 154485 2527 154543 2533
rect 155126 2524 155132 2576
rect 155184 2564 155190 2576
rect 155221 2567 155279 2573
rect 155221 2564 155233 2567
rect 155184 2536 155233 2564
rect 155184 2524 155190 2536
rect 155221 2533 155233 2536
rect 155267 2533 155279 2567
rect 155221 2527 155279 2533
rect 156230 2524 156236 2576
rect 156288 2564 156294 2576
rect 156417 2567 156475 2573
rect 156417 2564 156429 2567
rect 156288 2536 156429 2564
rect 156288 2524 156294 2536
rect 156417 2533 156429 2536
rect 156463 2533 156475 2567
rect 156417 2527 156475 2533
rect 157334 2524 157340 2576
rect 157392 2564 157398 2576
rect 157429 2567 157487 2573
rect 157429 2564 157441 2567
rect 157392 2536 157441 2564
rect 157392 2524 157398 2536
rect 157429 2533 157441 2536
rect 157475 2533 157487 2567
rect 159082 2564 159088 2576
rect 159043 2536 159088 2564
rect 157429 2527 157487 2533
rect 159082 2524 159088 2536
rect 159140 2524 159146 2576
rect 159726 2524 159732 2576
rect 159784 2564 159790 2576
rect 159821 2567 159879 2573
rect 159821 2564 159833 2567
rect 159784 2536 159833 2564
rect 159784 2524 159790 2536
rect 159821 2533 159833 2536
rect 159867 2533 159879 2567
rect 159821 2527 159879 2533
rect 160557 2567 160615 2573
rect 160557 2533 160569 2567
rect 160603 2564 160615 2567
rect 160646 2564 160652 2576
rect 160603 2536 160652 2564
rect 160603 2533 160615 2536
rect 160557 2527 160615 2533
rect 160646 2524 160652 2536
rect 160704 2524 160710 2576
rect 161750 2524 161756 2576
rect 161808 2564 161814 2576
rect 161845 2567 161903 2573
rect 161845 2564 161857 2567
rect 161808 2536 161857 2564
rect 161808 2524 161814 2536
rect 161845 2533 161857 2536
rect 161891 2533 161903 2567
rect 161845 2527 161903 2533
rect 162854 2524 162860 2576
rect 162912 2564 162918 2576
rect 162949 2567 163007 2573
rect 162949 2564 162961 2567
rect 162912 2536 162961 2564
rect 162912 2524 162918 2536
rect 162949 2533 162961 2536
rect 162995 2533 163007 2567
rect 162949 2527 163007 2533
rect 164326 2524 164332 2576
rect 164384 2564 164390 2576
rect 164421 2567 164479 2573
rect 164421 2564 164433 2567
rect 164384 2536 164433 2564
rect 164384 2524 164390 2536
rect 164421 2533 164433 2536
rect 164467 2533 164479 2567
rect 164421 2527 164479 2533
rect 165062 2524 165068 2576
rect 165120 2564 165126 2576
rect 165157 2567 165215 2573
rect 165157 2564 165169 2567
rect 165120 2536 165169 2564
rect 165120 2524 165126 2536
rect 165157 2533 165169 2536
rect 165203 2533 165215 2567
rect 167086 2564 167092 2576
rect 167047 2536 167092 2564
rect 165157 2527 165215 2533
rect 167086 2524 167092 2536
rect 167144 2524 167150 2576
rect 167270 2524 167276 2576
rect 167328 2564 167334 2576
rect 167825 2567 167883 2573
rect 167825 2564 167837 2567
rect 167328 2536 167837 2564
rect 167328 2524 167334 2536
rect 167825 2533 167837 2536
rect 167871 2533 167883 2567
rect 167825 2527 167883 2533
rect 168374 2524 168380 2576
rect 168432 2564 168438 2576
rect 168561 2567 168619 2573
rect 168561 2564 168573 2567
rect 168432 2536 168573 2564
rect 168432 2524 168438 2536
rect 168561 2533 168573 2536
rect 168607 2533 168619 2567
rect 169754 2564 169760 2576
rect 169715 2536 169760 2564
rect 168561 2527 168619 2533
rect 169754 2524 169760 2536
rect 169812 2524 169818 2576
rect 170582 2524 170588 2576
rect 170640 2564 170646 2576
rect 170677 2567 170735 2573
rect 170677 2564 170689 2567
rect 170640 2536 170689 2564
rect 170640 2524 170646 2536
rect 170677 2533 170689 2536
rect 170723 2533 170735 2567
rect 170677 2527 170735 2533
rect 171686 2524 171692 2576
rect 171744 2564 171750 2576
rect 172425 2567 172483 2573
rect 172425 2564 172437 2567
rect 171744 2536 172437 2564
rect 171744 2524 171750 2536
rect 172425 2533 172437 2536
rect 172471 2533 172483 2567
rect 172425 2527 172483 2533
rect 172790 2524 172796 2576
rect 172848 2564 172854 2576
rect 173161 2567 173219 2573
rect 173161 2564 173173 2567
rect 172848 2536 173173 2564
rect 172848 2524 172854 2536
rect 173161 2533 173173 2536
rect 173207 2533 173219 2567
rect 173894 2564 173900 2576
rect 173855 2536 173900 2564
rect 173161 2527 173219 2533
rect 173894 2524 173900 2536
rect 173952 2524 173958 2576
rect 174998 2524 175004 2576
rect 175056 2564 175062 2576
rect 175093 2567 175151 2573
rect 175093 2564 175105 2567
rect 175056 2536 175105 2564
rect 175056 2524 175062 2536
rect 175093 2533 175105 2536
rect 175139 2533 175151 2567
rect 175093 2527 175151 2533
rect 176102 2524 176108 2576
rect 176160 2564 176166 2576
rect 176197 2567 176255 2573
rect 176197 2564 176209 2567
rect 176160 2536 176209 2564
rect 176160 2524 176166 2536
rect 176197 2533 176209 2536
rect 176243 2533 176255 2567
rect 176197 2527 176255 2533
rect 176930 2524 176936 2576
rect 176988 2564 176994 2576
rect 177761 2567 177819 2573
rect 177761 2564 177773 2567
rect 176988 2536 177773 2564
rect 176988 2524 176994 2536
rect 177761 2533 177773 2536
rect 177807 2533 177819 2567
rect 177761 2527 177819 2533
rect 89717 2499 89775 2505
rect 89717 2465 89729 2499
rect 89763 2496 89775 2499
rect 89990 2496 89996 2508
rect 89763 2468 89996 2496
rect 89763 2465 89775 2468
rect 89717 2459 89775 2465
rect 89990 2456 89996 2468
rect 90048 2456 90054 2508
rect 90266 2456 90272 2508
rect 90324 2496 90330 2508
rect 91189 2499 91247 2505
rect 91189 2496 91201 2499
rect 90324 2468 91201 2496
rect 90324 2456 90330 2468
rect 91189 2465 91201 2468
rect 91235 2465 91247 2499
rect 91189 2459 91247 2465
rect 92290 2456 92296 2508
rect 92348 2496 92354 2508
rect 92348 2468 92796 2496
rect 92348 2456 92354 2468
rect 92569 2431 92627 2437
rect 92569 2428 92581 2431
rect 89456 2400 92581 2428
rect 92569 2397 92581 2400
rect 92615 2397 92627 2431
rect 92768 2428 92796 2468
rect 93302 2456 93308 2508
rect 93360 2496 93366 2508
rect 95053 2499 95111 2505
rect 95053 2496 95065 2499
rect 93360 2468 95065 2496
rect 93360 2456 93366 2468
rect 95053 2465 95065 2468
rect 95099 2465 95111 2499
rect 95053 2459 95111 2465
rect 95142 2456 95148 2508
rect 95200 2496 95206 2508
rect 102502 2496 102508 2508
rect 95200 2468 102508 2496
rect 95200 2456 95206 2468
rect 102502 2456 102508 2468
rect 102560 2456 102566 2508
rect 108114 2456 108120 2508
rect 108172 2496 108178 2508
rect 108393 2499 108451 2505
rect 108393 2496 108405 2499
rect 108172 2468 108405 2496
rect 108172 2456 108178 2468
rect 108393 2465 108405 2468
rect 108439 2465 108451 2499
rect 108393 2459 108451 2465
rect 110322 2456 110328 2508
rect 110380 2496 110386 2508
rect 111061 2499 111119 2505
rect 111061 2496 111073 2499
rect 110380 2468 111073 2496
rect 110380 2456 110386 2468
rect 111061 2465 111073 2468
rect 111107 2465 111119 2499
rect 111061 2459 111119 2465
rect 132678 2456 132684 2508
rect 132736 2496 132742 2508
rect 133785 2499 133843 2505
rect 133785 2496 133797 2499
rect 132736 2468 133797 2496
rect 132736 2456 132742 2468
rect 133785 2465 133797 2468
rect 133831 2465 133843 2499
rect 133785 2459 133843 2465
rect 151446 2456 151452 2508
rect 151504 2496 151510 2508
rect 152553 2499 152611 2505
rect 152553 2496 152565 2499
rect 151504 2468 152565 2496
rect 151504 2456 151510 2468
rect 152553 2465 152565 2468
rect 152599 2465 152611 2499
rect 152553 2459 152611 2465
rect 164694 2456 164700 2508
rect 164752 2496 164758 2508
rect 165801 2499 165859 2505
rect 165801 2496 165813 2499
rect 164752 2468 165813 2496
rect 164752 2456 164758 2468
rect 165801 2465 165813 2468
rect 165847 2465 165859 2499
rect 165801 2459 165859 2465
rect 95237 2431 95295 2437
rect 95237 2428 95249 2431
rect 92768 2400 95249 2428
rect 92569 2391 92627 2397
rect 95237 2397 95249 2400
rect 95283 2397 95295 2431
rect 95237 2391 95295 2397
rect 95602 2388 95608 2440
rect 95660 2428 95666 2440
rect 97905 2431 97963 2437
rect 97905 2428 97917 2431
rect 95660 2400 97917 2428
rect 95660 2388 95666 2400
rect 97905 2397 97917 2400
rect 97951 2397 97963 2431
rect 97905 2391 97963 2397
rect 97994 2388 98000 2440
rect 98052 2428 98058 2440
rect 99377 2431 99435 2437
rect 99377 2428 99389 2431
rect 98052 2400 99389 2428
rect 98052 2388 98058 2400
rect 99377 2397 99389 2400
rect 99423 2397 99435 2431
rect 99377 2391 99435 2397
rect 100018 2388 100024 2440
rect 100076 2428 100082 2440
rect 101309 2431 101367 2437
rect 101309 2428 101321 2431
rect 100076 2400 101321 2428
rect 100076 2388 100082 2400
rect 101309 2397 101321 2400
rect 101355 2397 101367 2431
rect 101309 2391 101367 2397
rect 107746 2388 107752 2440
rect 107804 2428 107810 2440
rect 109313 2431 109371 2437
rect 109313 2428 109325 2431
rect 107804 2400 109325 2428
rect 107804 2388 107810 2400
rect 109313 2397 109325 2400
rect 109359 2397 109371 2431
rect 109313 2391 109371 2397
rect 109954 2388 109960 2440
rect 110012 2428 110018 2440
rect 111981 2431 112039 2437
rect 111981 2428 111993 2431
rect 110012 2400 111993 2428
rect 110012 2388 110018 2400
rect 111981 2397 111993 2400
rect 112027 2397 112039 2431
rect 111981 2391 112039 2397
rect 90358 2360 90364 2372
rect 83056 2332 84884 2360
rect 85592 2332 87368 2360
rect 87432 2332 89116 2360
rect 89180 2332 90364 2360
rect 83056 2320 83062 2332
rect 76653 2295 76711 2301
rect 76653 2292 76665 2295
rect 75472 2264 76665 2292
rect 72476 2252 72482 2264
rect 76653 2261 76665 2264
rect 76699 2261 76711 2295
rect 76653 2255 76711 2261
rect 76837 2295 76895 2301
rect 76837 2261 76849 2295
rect 76883 2261 76895 2295
rect 76837 2255 76895 2261
rect 76926 2252 76932 2304
rect 76984 2292 76990 2304
rect 77849 2295 77907 2301
rect 77849 2292 77861 2295
rect 76984 2264 77861 2292
rect 76984 2252 76990 2264
rect 77849 2261 77861 2264
rect 77895 2261 77907 2295
rect 77849 2255 77907 2261
rect 80149 2295 80207 2301
rect 80149 2261 80161 2295
rect 80195 2292 80207 2295
rect 80238 2292 80244 2304
rect 80195 2264 80244 2292
rect 80195 2261 80207 2264
rect 80149 2255 80207 2261
rect 80238 2252 80244 2264
rect 80296 2252 80302 2304
rect 80330 2252 80336 2304
rect 80388 2292 80394 2304
rect 82446 2292 82452 2304
rect 80388 2264 82452 2292
rect 80388 2252 80394 2264
rect 82446 2252 82452 2264
rect 82504 2252 82510 2304
rect 82630 2252 82636 2304
rect 82688 2292 82694 2304
rect 84562 2292 84568 2304
rect 82688 2264 84568 2292
rect 82688 2252 82694 2264
rect 84562 2252 84568 2264
rect 84620 2292 84626 2304
rect 84749 2295 84807 2301
rect 84749 2292 84761 2295
rect 84620 2264 84761 2292
rect 84620 2252 84626 2264
rect 84749 2261 84761 2264
rect 84795 2261 84807 2295
rect 84856 2292 84884 2332
rect 85761 2295 85819 2301
rect 85761 2292 85773 2295
rect 84856 2264 85773 2292
rect 84749 2255 84807 2261
rect 85761 2261 85773 2264
rect 85807 2261 85819 2295
rect 86954 2292 86960 2304
rect 86915 2264 86960 2292
rect 85761 2255 85819 2261
rect 86954 2252 86960 2264
rect 87012 2252 87018 2304
rect 87046 2252 87052 2304
rect 87104 2292 87110 2304
rect 87141 2295 87199 2301
rect 87141 2292 87153 2295
rect 87104 2264 87153 2292
rect 87104 2252 87110 2264
rect 87141 2261 87153 2264
rect 87187 2261 87199 2295
rect 87340 2292 87368 2332
rect 87414 2292 87420 2304
rect 87340 2264 87420 2292
rect 87141 2255 87199 2261
rect 87414 2252 87420 2264
rect 87472 2252 87478 2304
rect 87966 2292 87972 2304
rect 87927 2264 87972 2292
rect 87966 2252 87972 2264
rect 88024 2252 88030 2304
rect 88058 2252 88064 2304
rect 88116 2292 88122 2304
rect 88153 2295 88211 2301
rect 88153 2292 88165 2295
rect 88116 2264 88165 2292
rect 88116 2252 88122 2264
rect 88153 2261 88165 2264
rect 88199 2261 88211 2295
rect 89088 2292 89116 2332
rect 90358 2320 90364 2332
rect 90416 2320 90422 2372
rect 90634 2360 90640 2372
rect 90595 2332 90640 2360
rect 90634 2320 90640 2332
rect 90692 2320 90698 2372
rect 91370 2320 91376 2372
rect 91428 2360 91434 2372
rect 94041 2363 94099 2369
rect 94041 2360 94053 2363
rect 91428 2332 94053 2360
rect 91428 2320 91434 2332
rect 94041 2329 94053 2332
rect 94087 2329 94099 2363
rect 94041 2323 94099 2329
rect 94498 2320 94504 2372
rect 94556 2360 94562 2372
rect 94556 2332 96660 2360
rect 94556 2320 94562 2332
rect 90266 2292 90272 2304
rect 89088 2264 90272 2292
rect 88153 2255 88211 2261
rect 90266 2252 90272 2264
rect 90324 2252 90330 2304
rect 91278 2292 91284 2304
rect 91239 2264 91284 2292
rect 91278 2252 91284 2264
rect 91336 2252 91342 2304
rect 92566 2252 92572 2304
rect 92624 2292 92630 2304
rect 96632 2301 96660 2332
rect 96706 2320 96712 2372
rect 96764 2360 96770 2372
rect 98641 2363 98699 2369
rect 98641 2360 98653 2363
rect 96764 2332 98653 2360
rect 96764 2320 96770 2332
rect 98641 2329 98653 2332
rect 98687 2329 98699 2363
rect 98641 2323 98699 2329
rect 98914 2320 98920 2372
rect 98972 2360 98978 2372
rect 100573 2363 100631 2369
rect 100573 2360 100585 2363
rect 98972 2332 100585 2360
rect 98972 2320 98978 2332
rect 100573 2329 100585 2332
rect 100619 2329 100631 2363
rect 100573 2323 100631 2329
rect 101122 2320 101128 2372
rect 101180 2360 101186 2372
rect 102045 2363 102103 2369
rect 102045 2360 102057 2363
rect 101180 2332 102057 2360
rect 101180 2320 101186 2332
rect 102045 2329 102057 2332
rect 102091 2329 102103 2363
rect 102045 2323 102103 2329
rect 108850 2320 108856 2372
rect 108908 2360 108914 2372
rect 110049 2363 110107 2369
rect 110049 2360 110061 2363
rect 108908 2332 110061 2360
rect 108908 2320 108914 2332
rect 110049 2329 110061 2332
rect 110095 2329 110107 2363
rect 110049 2323 110107 2329
rect 111058 2320 111064 2372
rect 111116 2360 111122 2372
rect 111116 2332 112024 2360
rect 111116 2320 111122 2332
rect 93213 2295 93271 2301
rect 93213 2292 93225 2295
rect 92624 2264 93225 2292
rect 92624 2252 92630 2264
rect 93213 2261 93225 2264
rect 93259 2261 93271 2295
rect 93213 2255 93271 2261
rect 96617 2295 96675 2301
rect 96617 2261 96629 2295
rect 96663 2261 96675 2295
rect 96617 2255 96675 2261
rect 102226 2252 102232 2304
rect 102284 2292 102290 2304
rect 103149 2295 103207 2301
rect 103149 2292 103161 2295
rect 102284 2264 103161 2292
rect 102284 2252 102290 2264
rect 103149 2261 103161 2264
rect 103195 2261 103207 2295
rect 103149 2255 103207 2261
rect 103330 2252 103336 2304
rect 103388 2292 103394 2304
rect 103885 2295 103943 2301
rect 103885 2292 103897 2295
rect 103388 2264 103897 2292
rect 103388 2252 103394 2264
rect 103885 2261 103897 2264
rect 103931 2261 103943 2295
rect 103885 2255 103943 2261
rect 104434 2252 104440 2304
rect 104492 2292 104498 2304
rect 104621 2295 104679 2301
rect 104621 2292 104633 2295
rect 104492 2264 104633 2292
rect 104492 2252 104498 2264
rect 104621 2261 104633 2264
rect 104667 2261 104679 2295
rect 104621 2255 104679 2261
rect 105538 2252 105544 2304
rect 105596 2292 105602 2304
rect 105817 2295 105875 2301
rect 105817 2292 105829 2295
rect 105596 2264 105829 2292
rect 105596 2252 105602 2264
rect 105817 2261 105829 2264
rect 105863 2261 105875 2295
rect 105817 2255 105875 2261
rect 106642 2252 106648 2304
rect 106700 2292 106706 2304
rect 106829 2295 106887 2301
rect 106829 2292 106841 2295
rect 106700 2264 106841 2292
rect 106700 2252 106706 2264
rect 106829 2261 106841 2264
rect 106875 2261 106887 2295
rect 106829 2255 106887 2261
rect 106918 2252 106924 2304
rect 106976 2292 106982 2304
rect 108485 2295 108543 2301
rect 108485 2292 108497 2295
rect 106976 2264 108497 2292
rect 106976 2252 106982 2264
rect 108485 2261 108497 2264
rect 108531 2261 108543 2295
rect 111996 2292 112024 2332
rect 112162 2320 112168 2372
rect 112220 2360 112226 2372
rect 113913 2363 113971 2369
rect 113913 2360 113925 2363
rect 112220 2332 113925 2360
rect 112220 2320 112226 2332
rect 113913 2329 113925 2332
rect 113959 2329 113971 2363
rect 113913 2323 113971 2329
rect 114370 2320 114376 2372
rect 114428 2360 114434 2372
rect 115385 2363 115443 2369
rect 115385 2360 115397 2363
rect 114428 2332 115397 2360
rect 114428 2320 114434 2332
rect 115385 2329 115397 2332
rect 115431 2329 115443 2363
rect 115385 2323 115443 2329
rect 116578 2320 116584 2372
rect 116636 2360 116642 2372
rect 117317 2363 117375 2369
rect 117317 2360 117329 2363
rect 116636 2332 117329 2360
rect 116636 2320 116642 2332
rect 117317 2329 117329 2332
rect 117363 2329 117375 2363
rect 117317 2323 117375 2329
rect 125318 2320 125324 2372
rect 125376 2360 125382 2372
rect 125597 2363 125655 2369
rect 125597 2360 125609 2363
rect 125376 2332 125609 2360
rect 125376 2320 125382 2332
rect 125597 2329 125609 2332
rect 125643 2329 125655 2363
rect 125597 2323 125655 2329
rect 130838 2320 130844 2372
rect 130896 2360 130902 2372
rect 131117 2363 131175 2369
rect 131117 2360 131129 2363
rect 130896 2332 131129 2360
rect 130896 2320 130902 2332
rect 131117 2329 131129 2332
rect 131163 2329 131175 2363
rect 147398 2360 147404 2372
rect 147359 2332 147404 2360
rect 131117 2323 131175 2329
rect 147398 2320 147404 2332
rect 147456 2320 147462 2372
rect 174998 2320 175004 2372
rect 175056 2360 175062 2372
rect 175277 2363 175335 2369
rect 175277 2360 175289 2363
rect 175056 2332 175289 2360
rect 175056 2320 175062 2332
rect 175277 2329 175289 2332
rect 175323 2329 175335 2363
rect 175277 2323 175335 2329
rect 112625 2295 112683 2301
rect 112625 2292 112637 2295
rect 111996 2264 112637 2292
rect 108485 2255 108543 2261
rect 112625 2261 112637 2264
rect 112671 2261 112683 2295
rect 112625 2255 112683 2261
rect 113266 2252 113272 2304
rect 113324 2292 113330 2304
rect 114557 2295 114615 2301
rect 114557 2292 114569 2295
rect 113324 2264 114569 2292
rect 113324 2252 113330 2264
rect 114557 2261 114569 2264
rect 114603 2261 114615 2295
rect 114557 2255 114615 2261
rect 115474 2252 115480 2304
rect 115532 2292 115538 2304
rect 116489 2295 116547 2301
rect 116489 2292 116501 2295
rect 115532 2264 116501 2292
rect 115532 2252 115538 2264
rect 116489 2261 116501 2264
rect 116535 2261 116547 2295
rect 116489 2255 116547 2261
rect 117682 2252 117688 2304
rect 117740 2292 117746 2304
rect 117961 2295 118019 2301
rect 117961 2292 117973 2295
rect 117740 2264 117973 2292
rect 117740 2252 117746 2264
rect 117961 2261 117973 2264
rect 118007 2261 118019 2295
rect 117961 2255 118019 2261
rect 118786 2252 118792 2304
rect 118844 2292 118850 2304
rect 119157 2295 119215 2301
rect 119157 2292 119169 2295
rect 118844 2264 119169 2292
rect 118844 2252 118850 2264
rect 119157 2261 119169 2264
rect 119203 2261 119215 2295
rect 119157 2255 119215 2261
rect 119890 2252 119896 2304
rect 119948 2292 119954 2304
rect 120077 2295 120135 2301
rect 120077 2292 120089 2295
rect 119948 2264 120089 2292
rect 119948 2252 119954 2264
rect 120077 2261 120089 2264
rect 120123 2261 120135 2295
rect 120077 2255 120135 2261
rect 120902 2252 120908 2304
rect 120960 2292 120966 2304
rect 121825 2295 121883 2301
rect 121825 2292 121837 2295
rect 120960 2264 121837 2292
rect 120960 2252 120966 2264
rect 121825 2261 121837 2264
rect 121871 2261 121883 2295
rect 121825 2255 121883 2261
rect 122006 2252 122012 2304
rect 122064 2292 122070 2304
rect 122561 2295 122619 2301
rect 122561 2292 122573 2295
rect 122064 2264 122573 2292
rect 122064 2252 122070 2264
rect 122561 2261 122573 2264
rect 122607 2261 122619 2295
rect 122561 2255 122619 2261
rect 123110 2252 123116 2304
rect 123168 2292 123174 2304
rect 123297 2295 123355 2301
rect 123297 2292 123309 2295
rect 123168 2264 123309 2292
rect 123168 2252 123174 2264
rect 123297 2261 123309 2264
rect 123343 2261 123355 2295
rect 123297 2255 123355 2261
rect 124214 2252 124220 2304
rect 124272 2292 124278 2304
rect 124493 2295 124551 2301
rect 124493 2292 124505 2295
rect 124272 2264 124505 2292
rect 124272 2252 124278 2264
rect 124493 2261 124505 2264
rect 124539 2261 124551 2295
rect 124493 2255 124551 2261
rect 126422 2252 126428 2304
rect 126480 2292 126486 2304
rect 127161 2295 127219 2301
rect 127161 2292 127173 2295
rect 126480 2264 127173 2292
rect 126480 2252 126486 2264
rect 127161 2261 127173 2264
rect 127207 2261 127219 2295
rect 127161 2255 127219 2261
rect 127526 2252 127532 2304
rect 127584 2292 127590 2304
rect 127897 2295 127955 2301
rect 127897 2292 127909 2295
rect 127584 2264 127909 2292
rect 127584 2252 127590 2264
rect 127897 2261 127909 2264
rect 127943 2261 127955 2295
rect 128630 2292 128636 2304
rect 128591 2264 128636 2292
rect 127897 2255 127955 2261
rect 128630 2252 128636 2264
rect 128688 2252 128694 2304
rect 129734 2252 129740 2304
rect 129792 2292 129798 2304
rect 129921 2295 129979 2301
rect 129921 2292 129933 2295
rect 129792 2264 129933 2292
rect 129792 2252 129798 2264
rect 129921 2261 129933 2264
rect 129967 2261 129979 2295
rect 129921 2255 129979 2261
rect 131942 2252 131948 2304
rect 132000 2292 132006 2304
rect 132497 2295 132555 2301
rect 132497 2292 132509 2295
rect 132000 2264 132509 2292
rect 132000 2252 132006 2264
rect 132497 2261 132509 2264
rect 132543 2261 132555 2295
rect 132497 2255 132555 2261
rect 133046 2252 133052 2304
rect 133104 2292 133110 2304
rect 133233 2295 133291 2301
rect 133233 2292 133245 2295
rect 133104 2264 133245 2292
rect 133104 2252 133110 2264
rect 133233 2261 133245 2264
rect 133279 2261 133291 2295
rect 133233 2255 133291 2261
rect 134150 2252 134156 2304
rect 134208 2292 134214 2304
rect 135165 2295 135223 2301
rect 135165 2292 135177 2295
rect 134208 2264 135177 2292
rect 134208 2252 134214 2264
rect 135165 2261 135177 2264
rect 135211 2261 135223 2295
rect 135165 2255 135223 2261
rect 135254 2252 135260 2304
rect 135312 2292 135318 2304
rect 135901 2295 135959 2301
rect 135901 2292 135913 2295
rect 135312 2264 135913 2292
rect 135312 2252 135318 2264
rect 135901 2261 135913 2264
rect 135947 2261 135959 2295
rect 135901 2255 135959 2261
rect 136358 2252 136364 2304
rect 136416 2292 136422 2304
rect 136637 2295 136695 2301
rect 136637 2292 136649 2295
rect 136416 2264 136649 2292
rect 136416 2252 136422 2264
rect 136637 2261 136649 2264
rect 136683 2261 136695 2295
rect 136637 2255 136695 2261
rect 137462 2252 137468 2304
rect 137520 2292 137526 2304
rect 137833 2295 137891 2301
rect 137833 2292 137845 2295
rect 137520 2264 137845 2292
rect 137520 2252 137526 2264
rect 137833 2261 137845 2264
rect 137879 2261 137891 2295
rect 137833 2255 137891 2261
rect 138566 2252 138572 2304
rect 138624 2292 138630 2304
rect 138753 2295 138811 2301
rect 138753 2292 138765 2295
rect 138624 2264 138765 2292
rect 138624 2252 138630 2264
rect 138753 2261 138765 2264
rect 138799 2261 138811 2295
rect 138753 2255 138811 2261
rect 139670 2252 139676 2304
rect 139728 2292 139734 2304
rect 140501 2295 140559 2301
rect 140501 2292 140513 2295
rect 139728 2264 140513 2292
rect 139728 2252 139734 2264
rect 140501 2261 140513 2264
rect 140547 2261 140559 2295
rect 140501 2255 140559 2261
rect 140774 2252 140780 2304
rect 140832 2292 140838 2304
rect 141237 2295 141295 2301
rect 141237 2292 141249 2295
rect 140832 2264 141249 2292
rect 140832 2252 140838 2264
rect 141237 2261 141249 2264
rect 141283 2261 141295 2295
rect 141237 2255 141295 2261
rect 141878 2252 141884 2304
rect 141936 2292 141942 2304
rect 141973 2295 142031 2301
rect 141973 2292 141985 2295
rect 141936 2264 141985 2292
rect 141936 2252 141942 2264
rect 141973 2261 141985 2264
rect 142019 2261 142031 2295
rect 141973 2255 142031 2261
rect 142982 2252 142988 2304
rect 143040 2292 143046 2304
rect 143169 2295 143227 2301
rect 143169 2292 143181 2295
rect 143040 2264 143181 2292
rect 143040 2252 143046 2264
rect 143169 2261 143181 2264
rect 143215 2261 143227 2295
rect 143169 2255 143227 2261
rect 144086 2252 144092 2304
rect 144144 2292 144150 2304
rect 144273 2295 144331 2301
rect 144273 2292 144285 2295
rect 144144 2264 144285 2292
rect 144144 2252 144150 2264
rect 144273 2261 144285 2264
rect 144319 2261 144331 2295
rect 144273 2255 144331 2261
rect 145190 2252 145196 2304
rect 145248 2292 145254 2304
rect 145837 2295 145895 2301
rect 145837 2292 145849 2295
rect 145248 2264 145849 2292
rect 145248 2252 145254 2264
rect 145837 2261 145849 2264
rect 145883 2261 145895 2295
rect 145837 2255 145895 2261
rect 146294 2252 146300 2304
rect 146352 2292 146358 2304
rect 146573 2295 146631 2301
rect 146573 2292 146585 2295
rect 146352 2264 146585 2292
rect 146352 2252 146358 2264
rect 146573 2261 146585 2264
rect 146619 2261 146631 2295
rect 146573 2255 146631 2261
rect 148502 2252 148508 2304
rect 148560 2292 148566 2304
rect 148689 2295 148747 2301
rect 148689 2292 148701 2295
rect 148560 2264 148701 2292
rect 148560 2252 148566 2264
rect 148689 2261 148701 2264
rect 148735 2261 148747 2295
rect 148689 2255 148747 2261
rect 149606 2252 149612 2304
rect 149664 2292 149670 2304
rect 149793 2295 149851 2301
rect 149793 2292 149805 2295
rect 149664 2264 149805 2292
rect 149664 2252 149670 2264
rect 149793 2261 149805 2264
rect 149839 2261 149851 2295
rect 149793 2255 149851 2261
rect 150710 2252 150716 2304
rect 150768 2292 150774 2304
rect 151173 2295 151231 2301
rect 151173 2292 151185 2295
rect 150768 2264 151185 2292
rect 150768 2252 150774 2264
rect 151173 2261 151185 2264
rect 151219 2261 151231 2295
rect 151173 2255 151231 2261
rect 151814 2252 151820 2304
rect 151872 2292 151878 2304
rect 152001 2295 152059 2301
rect 152001 2292 152013 2295
rect 151872 2264 152013 2292
rect 151872 2252 151878 2264
rect 152001 2261 152013 2264
rect 152047 2261 152059 2295
rect 152001 2255 152059 2261
rect 152918 2252 152924 2304
rect 152976 2292 152982 2304
rect 153841 2295 153899 2301
rect 153841 2292 153853 2295
rect 152976 2264 153853 2292
rect 152976 2252 152982 2264
rect 153841 2261 153853 2264
rect 153887 2261 153899 2295
rect 153841 2255 153899 2261
rect 154022 2252 154028 2304
rect 154080 2292 154086 2304
rect 154577 2295 154635 2301
rect 154577 2292 154589 2295
rect 154080 2264 154589 2292
rect 154080 2252 154086 2264
rect 154577 2261 154589 2264
rect 154623 2261 154635 2295
rect 154577 2255 154635 2261
rect 155126 2252 155132 2304
rect 155184 2292 155190 2304
rect 155313 2295 155371 2301
rect 155313 2292 155325 2295
rect 155184 2264 155325 2292
rect 155184 2252 155190 2264
rect 155313 2261 155325 2264
rect 155359 2261 155371 2295
rect 155313 2255 155371 2261
rect 156230 2252 156236 2304
rect 156288 2292 156294 2304
rect 156509 2295 156567 2301
rect 156509 2292 156521 2295
rect 156288 2264 156521 2292
rect 156288 2252 156294 2264
rect 156509 2261 156521 2264
rect 156555 2261 156567 2295
rect 156509 2255 156567 2261
rect 157334 2252 157340 2304
rect 157392 2292 157398 2304
rect 157521 2295 157579 2301
rect 157521 2292 157533 2295
rect 157392 2264 157533 2292
rect 157392 2252 157398 2264
rect 157521 2261 157533 2264
rect 157567 2261 157579 2295
rect 157521 2255 157579 2261
rect 158438 2252 158444 2304
rect 158496 2292 158502 2304
rect 159177 2295 159235 2301
rect 159177 2292 159189 2295
rect 158496 2264 159189 2292
rect 158496 2252 158502 2264
rect 159177 2261 159189 2264
rect 159223 2261 159235 2295
rect 159177 2255 159235 2261
rect 159542 2252 159548 2304
rect 159600 2292 159606 2304
rect 159913 2295 159971 2301
rect 159913 2292 159925 2295
rect 159600 2264 159925 2292
rect 159600 2252 159606 2264
rect 159913 2261 159925 2264
rect 159959 2261 159971 2295
rect 160646 2292 160652 2304
rect 160607 2264 160652 2292
rect 159913 2255 159971 2261
rect 160646 2252 160652 2264
rect 160704 2252 160710 2304
rect 161750 2252 161756 2304
rect 161808 2292 161814 2304
rect 161937 2295 161995 2301
rect 161937 2292 161949 2295
rect 161808 2264 161949 2292
rect 161808 2252 161814 2264
rect 161937 2261 161949 2264
rect 161983 2261 161995 2295
rect 161937 2255 161995 2261
rect 162854 2252 162860 2304
rect 162912 2292 162918 2304
rect 163041 2295 163099 2301
rect 163041 2292 163053 2295
rect 162912 2264 163053 2292
rect 162912 2252 162918 2264
rect 163041 2261 163053 2264
rect 163087 2261 163099 2295
rect 163041 2255 163099 2261
rect 163958 2252 163964 2304
rect 164016 2292 164022 2304
rect 164513 2295 164571 2301
rect 164513 2292 164525 2295
rect 164016 2264 164525 2292
rect 164016 2252 164022 2264
rect 164513 2261 164525 2264
rect 164559 2261 164571 2295
rect 164513 2255 164571 2261
rect 165062 2252 165068 2304
rect 165120 2292 165126 2304
rect 165249 2295 165307 2301
rect 165249 2292 165261 2295
rect 165120 2264 165261 2292
rect 165120 2252 165126 2264
rect 165249 2261 165261 2264
rect 165295 2261 165307 2295
rect 165249 2255 165307 2261
rect 166166 2252 166172 2304
rect 166224 2292 166230 2304
rect 167181 2295 167239 2301
rect 167181 2292 167193 2295
rect 166224 2264 167193 2292
rect 166224 2252 166230 2264
rect 167181 2261 167193 2264
rect 167227 2261 167239 2295
rect 167181 2255 167239 2261
rect 167270 2252 167276 2304
rect 167328 2292 167334 2304
rect 167917 2295 167975 2301
rect 167917 2292 167929 2295
rect 167328 2264 167929 2292
rect 167328 2252 167334 2264
rect 167917 2261 167929 2264
rect 167963 2261 167975 2295
rect 167917 2255 167975 2261
rect 168374 2252 168380 2304
rect 168432 2292 168438 2304
rect 168653 2295 168711 2301
rect 168653 2292 168665 2295
rect 168432 2264 168665 2292
rect 168432 2252 168438 2264
rect 168653 2261 168665 2264
rect 168699 2261 168711 2295
rect 168653 2255 168711 2261
rect 169478 2252 169484 2304
rect 169536 2292 169542 2304
rect 169849 2295 169907 2301
rect 169849 2292 169861 2295
rect 169536 2264 169861 2292
rect 169536 2252 169542 2264
rect 169849 2261 169861 2264
rect 169895 2261 169907 2295
rect 169849 2255 169907 2261
rect 170582 2252 170588 2304
rect 170640 2292 170646 2304
rect 170769 2295 170827 2301
rect 170769 2292 170781 2295
rect 170640 2264 170781 2292
rect 170640 2252 170646 2264
rect 170769 2261 170781 2264
rect 170815 2261 170827 2295
rect 170769 2255 170827 2261
rect 171686 2252 171692 2304
rect 171744 2292 171750 2304
rect 172517 2295 172575 2301
rect 172517 2292 172529 2295
rect 171744 2264 172529 2292
rect 171744 2252 171750 2264
rect 172517 2261 172529 2264
rect 172563 2261 172575 2295
rect 172517 2255 172575 2261
rect 172790 2252 172796 2304
rect 172848 2292 172854 2304
rect 173253 2295 173311 2301
rect 173253 2292 173265 2295
rect 172848 2264 173265 2292
rect 172848 2252 172854 2264
rect 173253 2261 173265 2264
rect 173299 2261 173311 2295
rect 173253 2255 173311 2261
rect 173894 2252 173900 2304
rect 173952 2292 173958 2304
rect 173989 2295 174047 2301
rect 173989 2292 174001 2295
rect 173952 2264 174001 2292
rect 173952 2252 173958 2264
rect 173989 2261 174001 2264
rect 174035 2261 174047 2295
rect 173989 2255 174047 2261
rect 176102 2252 176108 2304
rect 176160 2292 176166 2304
rect 176289 2295 176347 2301
rect 176289 2292 176301 2295
rect 176160 2264 176301 2292
rect 176160 2252 176166 2264
rect 176289 2261 176301 2264
rect 176335 2261 176347 2295
rect 176289 2255 176347 2261
rect 177206 2252 177212 2304
rect 177264 2292 177270 2304
rect 177853 2295 177911 2301
rect 177853 2292 177865 2295
rect 177264 2264 177865 2292
rect 177264 2252 177270 2264
rect 177853 2261 177865 2264
rect 177899 2261 177911 2295
rect 177853 2255 177911 2261
rect 1104 2202 178848 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 34966 2202
rect 35018 2150 35030 2202
rect 35082 2150 35094 2202
rect 35146 2150 35158 2202
rect 35210 2150 65686 2202
rect 65738 2150 65750 2202
rect 65802 2150 65814 2202
rect 65866 2150 65878 2202
rect 65930 2150 96406 2202
rect 96458 2150 96470 2202
rect 96522 2150 96534 2202
rect 96586 2150 96598 2202
rect 96650 2150 127126 2202
rect 127178 2150 127190 2202
rect 127242 2150 127254 2202
rect 127306 2150 127318 2202
rect 127370 2150 157846 2202
rect 157898 2150 157910 2202
rect 157962 2150 157974 2202
rect 158026 2150 158038 2202
rect 158090 2150 178848 2202
rect 1104 2128 178848 2150
rect 8570 2048 8576 2100
rect 8628 2088 8634 2100
rect 33410 2088 33416 2100
rect 8628 2060 33416 2088
rect 8628 2048 8634 2060
rect 33410 2048 33416 2060
rect 33468 2048 33474 2100
rect 39114 2048 39120 2100
rect 39172 2088 39178 2100
rect 61197 2091 61255 2097
rect 61197 2088 61209 2091
rect 39172 2060 61209 2088
rect 39172 2048 39178 2060
rect 61197 2057 61209 2060
rect 61243 2057 61255 2091
rect 61197 2051 61255 2057
rect 61286 2048 61292 2100
rect 61344 2088 61350 2100
rect 72970 2088 72976 2100
rect 61344 2060 72976 2088
rect 61344 2048 61350 2060
rect 72970 2048 72976 2060
rect 73028 2048 73034 2100
rect 77110 2088 77116 2100
rect 77071 2060 77116 2088
rect 77110 2048 77116 2060
rect 77168 2048 77174 2100
rect 78582 2048 78588 2100
rect 78640 2088 78646 2100
rect 82262 2088 82268 2100
rect 78640 2060 82268 2088
rect 78640 2048 78646 2060
rect 82262 2048 82268 2060
rect 82320 2048 82326 2100
rect 82814 2048 82820 2100
rect 82872 2088 82878 2100
rect 90269 2091 90327 2097
rect 90269 2088 90281 2091
rect 82872 2060 90281 2088
rect 82872 2048 82878 2060
rect 90269 2057 90281 2060
rect 90315 2057 90327 2091
rect 90269 2051 90327 2057
rect 90358 2048 90364 2100
rect 90416 2088 90422 2100
rect 95142 2088 95148 2100
rect 90416 2060 95148 2088
rect 90416 2048 90422 2060
rect 95142 2048 95148 2060
rect 95200 2048 95206 2100
rect 9674 1980 9680 2032
rect 9732 2020 9738 2032
rect 15378 2020 15384 2032
rect 9732 1992 15384 2020
rect 9732 1980 9738 1992
rect 15378 1980 15384 1992
rect 15436 1980 15442 2032
rect 33778 1980 33784 2032
rect 33836 2020 33842 2032
rect 46934 2020 46940 2032
rect 33836 1992 46940 2020
rect 33836 1980 33842 1992
rect 46934 1980 46940 1992
rect 46992 1980 46998 2032
rect 47026 1980 47032 2032
rect 47084 2020 47090 2032
rect 48593 2023 48651 2029
rect 47084 1992 48544 2020
rect 47084 1980 47090 1992
rect 2774 1912 2780 1964
rect 2832 1952 2838 1964
rect 38746 1952 38752 1964
rect 2832 1924 38752 1952
rect 2832 1912 2838 1924
rect 38746 1912 38752 1924
rect 38804 1912 38810 1964
rect 42610 1912 42616 1964
rect 42668 1952 42674 1964
rect 45186 1952 45192 1964
rect 42668 1924 45192 1952
rect 42668 1912 42674 1924
rect 45186 1912 45192 1924
rect 45244 1912 45250 1964
rect 45370 1912 45376 1964
rect 45428 1952 45434 1964
rect 48314 1952 48320 1964
rect 45428 1924 48320 1952
rect 45428 1912 45434 1924
rect 48314 1912 48320 1924
rect 48372 1912 48378 1964
rect 48516 1952 48544 1992
rect 48593 1989 48605 2023
rect 48639 2020 48651 2023
rect 71958 2020 71964 2032
rect 48639 1992 71964 2020
rect 48639 1989 48651 1992
rect 48593 1983 48651 1989
rect 71958 1980 71964 1992
rect 72016 1980 72022 2032
rect 74534 1980 74540 2032
rect 74592 2020 74598 2032
rect 80330 2020 80336 2032
rect 74592 1992 80336 2020
rect 74592 1980 74598 1992
rect 80330 1980 80336 1992
rect 80388 1980 80394 2032
rect 84194 1980 84200 2032
rect 84252 2020 84258 2032
rect 87690 2020 87696 2032
rect 84252 1992 87696 2020
rect 84252 1980 84258 1992
rect 87690 1980 87696 1992
rect 87748 1980 87754 2032
rect 88334 1980 88340 2032
rect 88392 2020 88398 2032
rect 89622 2020 89628 2032
rect 88392 1992 89628 2020
rect 88392 1980 88398 1992
rect 89622 1980 89628 1992
rect 89680 1980 89686 2032
rect 63678 1952 63684 1964
rect 48516 1924 63684 1952
rect 63678 1912 63684 1924
rect 63736 1912 63742 1964
rect 65150 1912 65156 1964
rect 65208 1952 65214 1964
rect 87966 1952 87972 1964
rect 65208 1924 87972 1952
rect 65208 1912 65214 1924
rect 87966 1912 87972 1924
rect 88024 1912 88030 1964
rect 88150 1912 88156 1964
rect 88208 1952 88214 1964
rect 103146 1952 103152 1964
rect 88208 1924 103152 1952
rect 88208 1912 88214 1924
rect 103146 1912 103152 1924
rect 103204 1912 103210 1964
rect 7190 1844 7196 1896
rect 7248 1884 7254 1896
rect 33318 1884 33324 1896
rect 7248 1856 33324 1884
rect 7248 1844 7254 1856
rect 33318 1844 33324 1856
rect 33376 1844 33382 1896
rect 34514 1844 34520 1896
rect 34572 1884 34578 1896
rect 62666 1884 62672 1896
rect 34572 1856 62672 1884
rect 34572 1844 34578 1856
rect 62666 1844 62672 1856
rect 62724 1844 62730 1896
rect 71590 1844 71596 1896
rect 71648 1884 71654 1896
rect 76374 1884 76380 1896
rect 71648 1856 76380 1884
rect 71648 1844 71654 1856
rect 76374 1844 76380 1856
rect 76432 1884 76438 1896
rect 84010 1884 84016 1896
rect 76432 1856 84016 1884
rect 76432 1844 76438 1856
rect 84010 1844 84016 1856
rect 84068 1844 84074 1896
rect 85390 1844 85396 1896
rect 85448 1884 85454 1896
rect 88518 1884 88524 1896
rect 85448 1856 88524 1884
rect 85448 1844 85454 1856
rect 88518 1844 88524 1856
rect 88576 1844 88582 1896
rect 88613 1887 88671 1893
rect 88613 1853 88625 1887
rect 88659 1884 88671 1887
rect 92750 1884 92756 1896
rect 88659 1856 92756 1884
rect 88659 1853 88671 1856
rect 88613 1847 88671 1853
rect 92750 1844 92756 1856
rect 92808 1844 92814 1896
rect 32490 1776 32496 1828
rect 32548 1816 32554 1828
rect 43254 1816 43260 1828
rect 32548 1788 43260 1816
rect 32548 1776 32554 1788
rect 43254 1776 43260 1788
rect 43312 1776 43318 1828
rect 44726 1776 44732 1828
rect 44784 1816 44790 1828
rect 45370 1816 45376 1828
rect 44784 1788 45376 1816
rect 44784 1776 44790 1788
rect 45370 1776 45376 1788
rect 45428 1776 45434 1828
rect 47946 1776 47952 1828
rect 48004 1816 48010 1828
rect 53282 1816 53288 1828
rect 48004 1788 53288 1816
rect 48004 1776 48010 1788
rect 53282 1776 53288 1788
rect 53340 1776 53346 1828
rect 57606 1776 57612 1828
rect 57664 1816 57670 1828
rect 80238 1816 80244 1828
rect 57664 1788 80244 1816
rect 57664 1776 57670 1788
rect 80238 1776 80244 1788
rect 80296 1776 80302 1828
rect 82170 1816 82176 1828
rect 80532 1788 82176 1816
rect 37274 1708 37280 1760
rect 37332 1748 37338 1760
rect 62574 1748 62580 1760
rect 37332 1720 62580 1748
rect 37332 1708 37338 1720
rect 62574 1708 62580 1720
rect 62632 1708 62638 1760
rect 80054 1708 80060 1760
rect 80112 1748 80118 1760
rect 80532 1748 80560 1788
rect 82170 1776 82176 1788
rect 82228 1776 82234 1828
rect 83182 1776 83188 1828
rect 83240 1816 83246 1828
rect 85850 1816 85856 1828
rect 83240 1788 85856 1816
rect 83240 1776 83246 1788
rect 85850 1776 85856 1788
rect 85908 1776 85914 1828
rect 87322 1776 87328 1828
rect 87380 1816 87386 1828
rect 103054 1816 103060 1828
rect 87380 1788 103060 1816
rect 87380 1776 87386 1788
rect 103054 1776 103060 1788
rect 103112 1776 103118 1828
rect 80112 1720 80560 1748
rect 80112 1708 80118 1720
rect 80606 1708 80612 1760
rect 80664 1748 80670 1760
rect 90177 1751 90235 1757
rect 90177 1748 90189 1751
rect 80664 1720 90189 1748
rect 80664 1708 80670 1720
rect 90177 1717 90189 1720
rect 90223 1717 90235 1751
rect 90177 1711 90235 1717
rect 90269 1751 90327 1757
rect 90269 1717 90281 1751
rect 90315 1748 90327 1751
rect 98362 1748 98368 1760
rect 90315 1720 98368 1748
rect 90315 1717 90327 1720
rect 90269 1711 90327 1717
rect 98362 1708 98368 1720
rect 98420 1708 98426 1760
rect 20530 1640 20536 1692
rect 20588 1680 20594 1692
rect 47578 1680 47584 1692
rect 20588 1652 47584 1680
rect 20588 1640 20594 1652
rect 47578 1640 47584 1652
rect 47636 1640 47642 1692
rect 61197 1683 61255 1689
rect 61197 1649 61209 1683
rect 61243 1680 61255 1683
rect 66070 1680 66076 1692
rect 61243 1652 66076 1680
rect 61243 1649 61255 1652
rect 61197 1643 61255 1649
rect 66070 1640 66076 1652
rect 66128 1640 66134 1692
rect 86954 1680 86960 1692
rect 70366 1652 86960 1680
rect 31110 1572 31116 1624
rect 31168 1612 31174 1624
rect 41414 1612 41420 1624
rect 31168 1584 41420 1612
rect 31168 1572 31174 1584
rect 41414 1572 41420 1584
rect 41472 1572 41478 1624
rect 45830 1572 45836 1624
rect 45888 1612 45894 1624
rect 48593 1615 48651 1621
rect 48593 1612 48605 1615
rect 45888 1584 48605 1612
rect 45888 1572 45894 1584
rect 48593 1581 48605 1584
rect 48639 1581 48651 1615
rect 48593 1575 48651 1581
rect 63034 1572 63040 1624
rect 63092 1612 63098 1624
rect 70366 1612 70394 1652
rect 86954 1640 86960 1652
rect 87012 1640 87018 1692
rect 87049 1683 87107 1689
rect 87049 1649 87061 1683
rect 87095 1680 87107 1683
rect 93486 1680 93492 1692
rect 87095 1652 93492 1680
rect 87095 1649 87107 1652
rect 87049 1643 87107 1649
rect 93486 1640 93492 1652
rect 93544 1640 93550 1692
rect 106918 1680 106924 1692
rect 99346 1652 106924 1680
rect 63092 1584 70394 1612
rect 63092 1572 63098 1584
rect 73430 1572 73436 1624
rect 73488 1612 73494 1624
rect 85114 1612 85120 1624
rect 73488 1584 85120 1612
rect 73488 1572 73494 1584
rect 85114 1572 85120 1584
rect 85172 1572 85178 1624
rect 85206 1572 85212 1624
rect 85264 1612 85270 1624
rect 85264 1584 87184 1612
rect 85264 1572 85270 1584
rect 71406 1504 71412 1556
rect 71464 1544 71470 1556
rect 81434 1544 81440 1556
rect 71464 1516 81440 1544
rect 71464 1504 71470 1516
rect 81434 1504 81440 1516
rect 81492 1504 81498 1556
rect 82078 1504 82084 1556
rect 82136 1544 82142 1556
rect 87049 1547 87107 1553
rect 87049 1544 87061 1547
rect 82136 1516 87061 1544
rect 82136 1504 82142 1516
rect 87049 1513 87061 1516
rect 87095 1513 87107 1547
rect 87156 1544 87184 1584
rect 87230 1572 87236 1624
rect 87288 1612 87294 1624
rect 87782 1612 87788 1624
rect 87288 1584 87788 1612
rect 87288 1572 87294 1584
rect 87782 1572 87788 1584
rect 87840 1612 87846 1624
rect 99346 1612 99374 1652
rect 106918 1640 106924 1652
rect 106976 1640 106982 1692
rect 87840 1584 99374 1612
rect 87840 1572 87846 1584
rect 88613 1547 88671 1553
rect 88613 1544 88625 1547
rect 87156 1516 88625 1544
rect 87049 1507 87107 1513
rect 88613 1513 88625 1516
rect 88659 1513 88671 1547
rect 88613 1507 88671 1513
rect 90177 1547 90235 1553
rect 90177 1513 90189 1547
rect 90223 1544 90235 1547
rect 97626 1544 97632 1556
rect 90223 1516 97632 1544
rect 90223 1513 90235 1516
rect 90177 1507 90235 1513
rect 97626 1504 97632 1516
rect 97684 1504 97690 1556
rect 75730 1436 75736 1488
rect 75788 1476 75794 1488
rect 77018 1476 77024 1488
rect 75788 1448 77024 1476
rect 75788 1436 75794 1448
rect 77018 1436 77024 1448
rect 77076 1436 77082 1488
rect 77113 1479 77171 1485
rect 77113 1445 77125 1479
rect 77159 1476 77171 1479
rect 91646 1476 91652 1488
rect 77159 1448 91652 1476
rect 77159 1445 77171 1448
rect 77113 1439 77171 1445
rect 91646 1436 91652 1448
rect 91704 1436 91710 1488
rect 74626 1368 74632 1420
rect 74684 1408 74690 1420
rect 76926 1408 76932 1420
rect 74684 1380 76932 1408
rect 74684 1368 74690 1380
rect 76926 1368 76932 1380
rect 76984 1368 76990 1420
rect 84562 1368 84568 1420
rect 84620 1408 84626 1420
rect 90634 1408 90640 1420
rect 84620 1380 90640 1408
rect 84620 1368 84626 1380
rect 90634 1368 90640 1380
rect 90692 1368 90698 1420
rect 35618 1300 35624 1352
rect 35676 1340 35682 1352
rect 70302 1340 70308 1352
rect 35676 1312 70308 1340
rect 35676 1300 35682 1312
rect 70302 1300 70308 1312
rect 70360 1300 70366 1352
rect 85666 1300 85672 1352
rect 85724 1340 85730 1352
rect 91278 1340 91284 1352
rect 85724 1312 91284 1340
rect 85724 1300 85730 1312
rect 91278 1300 91284 1312
rect 91336 1300 91342 1352
rect 36722 1232 36728 1284
rect 36780 1272 36786 1284
rect 71498 1272 71504 1284
rect 36780 1244 71504 1272
rect 36780 1232 36786 1244
rect 71498 1232 71504 1244
rect 71556 1232 71562 1284
rect 83458 1232 83464 1284
rect 83516 1272 83522 1284
rect 89806 1272 89812 1284
rect 83516 1244 89812 1272
rect 83516 1232 83522 1244
rect 89806 1232 89812 1244
rect 89864 1232 89870 1284
rect 32950 1164 32956 1216
rect 33008 1204 33014 1216
rect 66622 1204 66628 1216
rect 33008 1176 66628 1204
rect 33008 1164 33014 1176
rect 66622 1164 66628 1176
rect 66680 1164 66686 1216
rect 34422 1096 34428 1148
rect 34480 1136 34486 1148
rect 67726 1136 67732 1148
rect 34480 1108 67732 1136
rect 34480 1096 34486 1108
rect 67726 1096 67732 1108
rect 67784 1096 67790 1148
rect 68738 1096 68744 1148
rect 68796 1136 68802 1148
rect 69566 1136 69572 1148
rect 68796 1108 69572 1136
rect 68796 1096 68802 1108
rect 69566 1096 69572 1108
rect 69624 1096 69630 1148
rect 15286 1028 15292 1080
rect 15344 1068 15350 1080
rect 41506 1068 41512 1080
rect 15344 1040 41512 1068
rect 15344 1028 15350 1040
rect 41506 1028 41512 1040
rect 41564 1028 41570 1080
rect 43622 1028 43628 1080
rect 43680 1068 43686 1080
rect 75546 1068 75552 1080
rect 43680 1040 75552 1068
rect 43680 1028 43686 1040
rect 75546 1028 75552 1040
rect 75604 1028 75610 1080
rect 43898 960 43904 1012
rect 43956 1000 43962 1012
rect 75270 1000 75276 1012
rect 43956 972 75276 1000
rect 43956 960 43962 972
rect 75270 960 75276 972
rect 75328 960 75334 1012
rect 88610 960 88616 1012
rect 88668 1000 88674 1012
rect 90174 1000 90180 1012
rect 88668 972 90180 1000
rect 88668 960 88674 972
rect 90174 960 90180 972
rect 90232 960 90238 1012
rect 27338 892 27344 944
rect 27396 932 27402 944
rect 58250 932 58256 944
rect 27396 904 58256 932
rect 27396 892 27402 904
rect 58250 892 58256 904
rect 58308 892 58314 944
rect 24118 824 24124 876
rect 24176 864 24182 876
rect 54754 864 54760 876
rect 24176 836 54760 864
rect 24176 824 24182 836
rect 54754 824 54760 836
rect 54812 824 54818 876
rect 28626 756 28632 808
rect 28684 796 28690 808
rect 58066 796 58072 808
rect 28684 768 58072 796
rect 28684 756 28690 768
rect 58066 756 58072 768
rect 58124 756 58130 808
rect 26602 688 26608 740
rect 26660 728 26666 740
rect 57146 728 57152 740
rect 26660 700 57152 728
rect 26660 688 26666 700
rect 57146 688 57152 700
rect 57204 688 57210 740
rect 29730 620 29736 672
rect 29788 660 29794 672
rect 59814 660 59820 672
rect 29788 632 59820 660
rect 29788 620 29794 632
rect 59814 620 59820 632
rect 59872 620 59878 672
rect 39298 552 39304 604
rect 39356 592 39362 604
rect 68830 592 68836 604
rect 39356 564 68836 592
rect 39356 552 39362 564
rect 68830 552 68836 564
rect 68888 552 68894 604
rect 31570 484 31576 536
rect 31628 524 31634 536
rect 56962 524 56968 536
rect 31628 496 56968 524
rect 31628 484 31634 496
rect 56962 484 56968 496
rect 57020 484 57026 536
rect 23106 416 23112 468
rect 23164 456 23170 468
rect 52914 456 52920 468
rect 23164 428 52920 456
rect 23164 416 23170 428
rect 52914 416 52920 428
rect 52972 416 52978 468
rect 20898 348 20904 400
rect 20956 388 20962 400
rect 48406 388 48412 400
rect 20956 360 48412 388
rect 20956 348 20962 360
rect 48406 348 48412 360
rect 48464 348 48470 400
rect 21910 280 21916 332
rect 21968 320 21974 332
rect 52546 320 52552 332
rect 21968 292 52552 320
rect 21968 280 21974 292
rect 52546 280 52552 292
rect 52604 280 52610 332
rect 25958 212 25964 264
rect 26016 252 26022 264
rect 55766 252 55772 264
rect 26016 224 55772 252
rect 26016 212 26022 224
rect 55766 212 55772 224
rect 55824 212 55830 264
rect 17770 144 17776 196
rect 17828 184 17834 196
rect 44634 184 44640 196
rect 17828 156 44640 184
rect 17828 144 17834 156
rect 44634 144 44640 156
rect 44692 144 44698 196
rect 16390 76 16396 128
rect 16448 116 16454 128
rect 44358 116 44364 128
rect 16448 88 44364 116
rect 16448 76 16454 88
rect 44358 76 44364 88
rect 44416 76 44422 128
<< via1 >>
rect 4246 117478 4298 117530
rect 4310 117478 4362 117530
rect 4374 117478 4426 117530
rect 4438 117478 4490 117530
rect 34966 117478 35018 117530
rect 35030 117478 35082 117530
rect 35094 117478 35146 117530
rect 35158 117478 35210 117530
rect 65686 117478 65738 117530
rect 65750 117478 65802 117530
rect 65814 117478 65866 117530
rect 65878 117478 65930 117530
rect 96406 117478 96458 117530
rect 96470 117478 96522 117530
rect 96534 117478 96586 117530
rect 96598 117478 96650 117530
rect 127126 117478 127178 117530
rect 127190 117478 127242 117530
rect 127254 117478 127306 117530
rect 127318 117478 127370 117530
rect 157846 117478 157898 117530
rect 157910 117478 157962 117530
rect 157974 117478 158026 117530
rect 158038 117478 158090 117530
rect 2320 117240 2372 117292
rect 3884 117240 3936 117292
rect 7012 117240 7064 117292
rect 8576 117240 8628 117292
rect 11704 117240 11756 117292
rect 13268 117240 13320 117292
rect 16580 117240 16632 117292
rect 17960 117240 18012 117292
rect 21088 117240 21140 117292
rect 22652 117240 22704 117292
rect 25780 117240 25832 117292
rect 27344 117283 27396 117292
rect 27344 117249 27353 117283
rect 27353 117249 27387 117283
rect 27387 117249 27396 117283
rect 27344 117240 27396 117249
rect 30472 117240 30524 117292
rect 32036 117240 32088 117292
rect 35348 117283 35400 117292
rect 35348 117249 35357 117283
rect 35357 117249 35391 117283
rect 35391 117249 35400 117283
rect 35348 117240 35400 117249
rect 36728 117240 36780 117292
rect 40040 117240 40092 117292
rect 41420 117240 41472 117292
rect 44548 117240 44600 117292
rect 46112 117240 46164 117292
rect 49240 117240 49292 117292
rect 51080 117283 51132 117292
rect 51080 117249 51089 117283
rect 51089 117249 51123 117283
rect 51123 117249 51132 117283
rect 51080 117240 51132 117249
rect 53932 117240 53984 117292
rect 55496 117240 55548 117292
rect 58624 117240 58676 117292
rect 60188 117240 60240 117292
rect 63500 117240 63552 117292
rect 64880 117240 64932 117292
rect 68008 117240 68060 117292
rect 69572 117240 69624 117292
rect 72700 117283 72752 117292
rect 72700 117249 72709 117283
rect 72709 117249 72743 117283
rect 72743 117249 72752 117283
rect 72700 117240 72752 117249
rect 74264 117240 74316 117292
rect 77392 117240 77444 117292
rect 78956 117240 79008 117292
rect 756 117172 808 117224
rect 5448 117215 5500 117224
rect 5448 117181 5457 117215
rect 5457 117181 5491 117215
rect 5491 117181 5500 117215
rect 5448 117172 5500 117181
rect 10140 117215 10192 117224
rect 10140 117181 10149 117215
rect 10149 117181 10183 117215
rect 10183 117181 10192 117215
rect 10140 117172 10192 117181
rect 14832 117172 14884 117224
rect 19524 117172 19576 117224
rect 24216 117215 24268 117224
rect 24216 117181 24225 117215
rect 24225 117181 24259 117215
rect 24259 117181 24268 117215
rect 24216 117172 24268 117181
rect 28908 117215 28960 117224
rect 28908 117181 28917 117215
rect 28917 117181 28951 117215
rect 28951 117181 28960 117215
rect 28908 117172 28960 117181
rect 33600 117215 33652 117224
rect 33600 117181 33609 117215
rect 33609 117181 33643 117215
rect 33643 117181 33652 117215
rect 33600 117172 33652 117181
rect 35256 117172 35308 117224
rect 38292 117172 38344 117224
rect 42984 117215 43036 117224
rect 42984 117181 42993 117215
rect 42993 117181 43027 117215
rect 43027 117181 43036 117215
rect 42984 117172 43036 117181
rect 47676 117215 47728 117224
rect 47676 117181 47685 117215
rect 47685 117181 47719 117215
rect 47719 117181 47728 117215
rect 47676 117172 47728 117181
rect 52368 117215 52420 117224
rect 52368 117181 52377 117215
rect 52377 117181 52411 117215
rect 52411 117181 52420 117215
rect 52368 117172 52420 117181
rect 57060 117172 57112 117224
rect 61752 117215 61804 117224
rect 61752 117181 61761 117215
rect 61761 117181 61795 117215
rect 61795 117181 61804 117215
rect 61752 117172 61804 117181
rect 66444 117215 66496 117224
rect 66444 117181 66453 117215
rect 66453 117181 66487 117215
rect 66487 117181 66496 117215
rect 66444 117172 66496 117181
rect 71136 117215 71188 117224
rect 71136 117181 71145 117215
rect 71145 117181 71179 117215
rect 71179 117181 71188 117215
rect 71136 117172 71188 117181
rect 75828 117172 75880 117224
rect 76932 117172 76984 117224
rect 80520 117215 80572 117224
rect 80520 117181 80529 117215
rect 80529 117181 80563 117215
rect 80563 117181 80572 117215
rect 80520 117172 80572 117181
rect 82084 117240 82136 117292
rect 83648 117240 83700 117292
rect 86960 117240 87012 117292
rect 88340 117240 88392 117292
rect 91560 117240 91612 117292
rect 93124 117240 93176 117292
rect 96252 117240 96304 117292
rect 97816 117283 97868 117292
rect 97816 117249 97825 117283
rect 97825 117249 97859 117283
rect 97859 117249 97868 117283
rect 97816 117240 97868 117249
rect 100944 117240 100996 117292
rect 102508 117240 102560 117292
rect 105636 117240 105688 117292
rect 107200 117240 107252 117292
rect 110420 117240 110472 117292
rect 111892 117240 111944 117292
rect 115020 117240 115072 117292
rect 116584 117240 116636 117292
rect 119712 117240 119764 117292
rect 121460 117240 121512 117292
rect 124404 117240 124456 117292
rect 125968 117240 126020 117292
rect 129096 117240 129148 117292
rect 130660 117240 130712 117292
rect 133880 117240 133932 117292
rect 135352 117240 135404 117292
rect 138480 117240 138532 117292
rect 140044 117240 140096 117292
rect 143172 117240 143224 117292
rect 144736 117283 144788 117292
rect 144736 117249 144745 117283
rect 144745 117249 144779 117283
rect 144779 117249 144788 117283
rect 144736 117240 144788 117249
rect 147864 117240 147916 117292
rect 149428 117240 149480 117292
rect 152556 117240 152608 117292
rect 154120 117240 154172 117292
rect 157340 117240 157392 117292
rect 158812 117240 158864 117292
rect 161940 117240 161992 117292
rect 163504 117240 163556 117292
rect 166632 117240 166684 117292
rect 168380 117240 168432 117292
rect 171324 117240 171376 117292
rect 172888 117240 172940 117292
rect 176016 117240 176068 117292
rect 177580 117240 177632 117292
rect 85212 117215 85264 117224
rect 85212 117181 85221 117215
rect 85221 117181 85255 117215
rect 85255 117181 85264 117215
rect 85212 117172 85264 117181
rect 89904 117215 89956 117224
rect 89904 117181 89913 117215
rect 89913 117181 89947 117215
rect 89947 117181 89956 117215
rect 89904 117172 89956 117181
rect 94688 117172 94740 117224
rect 97632 117172 97684 117224
rect 99380 117172 99432 117224
rect 104072 117215 104124 117224
rect 104072 117181 104081 117215
rect 104081 117181 104115 117215
rect 104115 117181 104124 117215
rect 104072 117172 104124 117181
rect 108764 117215 108816 117224
rect 108764 117181 108773 117215
rect 108773 117181 108807 117215
rect 108807 117181 108816 117215
rect 108764 117172 108816 117181
rect 113456 117172 113508 117224
rect 118148 117172 118200 117224
rect 122840 117215 122892 117224
rect 122840 117181 122849 117215
rect 122849 117181 122883 117215
rect 122883 117181 122892 117215
rect 127532 117215 127584 117224
rect 122840 117172 122892 117181
rect 127532 117181 127541 117215
rect 127541 117181 127575 117215
rect 127575 117181 127584 117215
rect 127532 117172 127584 117181
rect 132224 117172 132276 117224
rect 136916 117172 136968 117224
rect 141608 117215 141660 117224
rect 141608 117181 141617 117215
rect 141617 117181 141651 117215
rect 141651 117181 141660 117215
rect 141608 117172 141660 117181
rect 146300 117215 146352 117224
rect 146300 117181 146309 117215
rect 146309 117181 146343 117215
rect 146343 117181 146352 117215
rect 146300 117172 146352 117181
rect 150992 117215 151044 117224
rect 150992 117181 151001 117215
rect 151001 117181 151035 117215
rect 151035 117181 151044 117215
rect 150992 117172 151044 117181
rect 155684 117172 155736 117224
rect 160376 117215 160428 117224
rect 160376 117181 160385 117215
rect 160385 117181 160419 117215
rect 160419 117181 160428 117215
rect 160376 117172 160428 117181
rect 165068 117215 165120 117224
rect 165068 117181 165077 117215
rect 165077 117181 165111 117215
rect 165111 117181 165120 117215
rect 165068 117172 165120 117181
rect 169760 117215 169812 117224
rect 169760 117181 169769 117215
rect 169769 117181 169803 117215
rect 169803 117181 169812 117215
rect 169760 117172 169812 117181
rect 174452 117172 174504 117224
rect 179144 117172 179196 117224
rect 2412 117147 2464 117156
rect 2412 117113 2421 117147
rect 2421 117113 2455 117147
rect 2455 117113 2464 117147
rect 2412 117104 2464 117113
rect 4344 117147 4396 117156
rect 4344 117113 4353 117147
rect 4353 117113 4387 117147
rect 4387 117113 4396 117147
rect 4344 117104 4396 117113
rect 8300 117104 8352 117156
rect 8484 117147 8536 117156
rect 8484 117113 8493 117147
rect 8493 117113 8527 117147
rect 8527 117113 8536 117147
rect 8484 117104 8536 117113
rect 12348 117147 12400 117156
rect 12348 117113 12357 117147
rect 12357 117113 12391 117147
rect 12391 117113 12400 117147
rect 12348 117104 12400 117113
rect 13360 117147 13412 117156
rect 13360 117113 13369 117147
rect 13369 117113 13403 117147
rect 13403 117113 13412 117147
rect 13360 117104 13412 117113
rect 16488 117147 16540 117156
rect 16488 117113 16497 117147
rect 16497 117113 16531 117147
rect 16531 117113 16540 117147
rect 16488 117104 16540 117113
rect 18052 117147 18104 117156
rect 18052 117113 18061 117147
rect 18061 117113 18095 117147
rect 18095 117113 18104 117147
rect 18052 117104 18104 117113
rect 22560 117104 22612 117156
rect 23020 117147 23072 117156
rect 23020 117113 23029 117147
rect 23029 117113 23063 117147
rect 23063 117113 23072 117147
rect 23020 117104 23072 117113
rect 26516 117104 26568 117156
rect 30840 117104 30892 117156
rect 32128 117147 32180 117156
rect 32128 117113 32137 117147
rect 32137 117113 32171 117147
rect 32171 117113 32180 117147
rect 32128 117104 32180 117113
rect 36820 117147 36872 117156
rect 36820 117113 36829 117147
rect 36829 117113 36863 117147
rect 36863 117113 36872 117147
rect 36820 117104 36872 117113
rect 39764 117104 39816 117156
rect 41696 117147 41748 117156
rect 41696 117113 41705 117147
rect 41705 117113 41739 117147
rect 41739 117113 41748 117147
rect 41696 117104 41748 117113
rect 44364 117104 44416 117156
rect 47032 117147 47084 117156
rect 47032 117113 47041 117147
rect 47041 117113 47075 117147
rect 47075 117113 47084 117147
rect 47032 117104 47084 117113
rect 48964 117104 49016 117156
rect 50896 117147 50948 117156
rect 50896 117113 50905 117147
rect 50905 117113 50939 117147
rect 50939 117113 50948 117147
rect 50896 117104 50948 117113
rect 54024 117104 54076 117156
rect 55588 117147 55640 117156
rect 55588 117113 55597 117147
rect 55597 117113 55631 117147
rect 55631 117113 55640 117147
rect 55588 117104 55640 117113
rect 58256 117104 58308 117156
rect 60372 117147 60424 117156
rect 60372 117113 60381 117147
rect 60381 117113 60415 117147
rect 60415 117113 60424 117147
rect 60372 117104 60424 117113
rect 62948 117104 63000 117156
rect 65524 117104 65576 117156
rect 67640 117104 67692 117156
rect 69664 117147 69716 117156
rect 69664 117113 69673 117147
rect 69673 117113 69707 117147
rect 69707 117113 69716 117147
rect 69664 117104 69716 117113
rect 72424 117104 72476 117156
rect 33416 117036 33468 117088
rect 69572 117036 69624 117088
rect 77116 117104 77168 117156
rect 79048 117147 79100 117156
rect 79048 117113 79057 117147
rect 79057 117113 79091 117147
rect 79091 117113 79100 117147
rect 79048 117104 79100 117113
rect 81808 117104 81860 117156
rect 86592 117104 86644 117156
rect 88432 117147 88484 117156
rect 88432 117113 88441 117147
rect 88441 117113 88475 117147
rect 88475 117113 88484 117147
rect 88432 117104 88484 117113
rect 91376 117104 91428 117156
rect 93216 117147 93268 117156
rect 93216 117113 93225 117147
rect 93225 117113 93259 117147
rect 93259 117113 93268 117147
rect 93216 117104 93268 117113
rect 96068 117104 96120 117156
rect 73068 117036 73120 117088
rect 97632 117079 97684 117088
rect 97632 117045 97641 117079
rect 97641 117045 97675 117079
rect 97675 117045 97684 117079
rect 101220 117104 101272 117156
rect 103060 117147 103112 117156
rect 103060 117113 103069 117147
rect 103069 117113 103103 117147
rect 103103 117113 103112 117147
rect 103060 117104 103112 117113
rect 105360 117104 105412 117156
rect 107200 117147 107252 117156
rect 107200 117113 107209 117147
rect 107209 117113 107243 117147
rect 107243 117113 107252 117147
rect 107200 117104 107252 117113
rect 110236 117104 110288 117156
rect 111156 117104 111208 117156
rect 114928 117104 114980 117156
rect 116676 117147 116728 117156
rect 116676 117113 116685 117147
rect 116685 117113 116719 117147
rect 116719 117113 116728 117147
rect 116676 117104 116728 117113
rect 119620 117104 119672 117156
rect 121736 117147 121788 117156
rect 121736 117113 121745 117147
rect 121745 117113 121779 117147
rect 121779 117113 121788 117147
rect 121736 117104 121788 117113
rect 124312 117104 124364 117156
rect 128912 117104 128964 117156
rect 130752 117147 130804 117156
rect 130752 117113 130761 117147
rect 130761 117113 130795 117147
rect 130795 117113 130804 117147
rect 130752 117104 130804 117113
rect 133512 117104 133564 117156
rect 135444 117147 135496 117156
rect 135444 117113 135453 117147
rect 135453 117113 135487 117147
rect 135487 117113 135496 117147
rect 135444 117104 135496 117113
rect 138020 117104 138072 117156
rect 140412 117147 140464 117156
rect 140412 117113 140421 117147
rect 140421 117113 140455 117147
rect 140455 117113 140464 117147
rect 140412 117104 140464 117113
rect 143172 117104 143224 117156
rect 144552 117147 144604 117156
rect 144552 117113 144561 117147
rect 144561 117113 144595 117147
rect 144595 117113 144604 117147
rect 144552 117104 144604 117113
rect 146760 117104 146812 117156
rect 149520 117147 149572 117156
rect 149520 117113 149529 117147
rect 149529 117113 149563 117147
rect 149563 117113 149572 117147
rect 149520 117104 149572 117113
rect 150900 117104 150952 117156
rect 154120 117104 154172 117156
rect 154856 117104 154908 117156
rect 159088 117147 159140 117156
rect 159088 117113 159097 117147
rect 159097 117113 159131 117147
rect 159131 117113 159140 117147
rect 159088 117104 159140 117113
rect 162032 117147 162084 117156
rect 162032 117113 162041 117147
rect 162041 117113 162075 117147
rect 162075 117113 162084 117147
rect 162032 117104 162084 117113
rect 164332 117104 164384 117156
rect 97632 117036 97684 117045
rect 162124 117036 162176 117088
rect 168196 117104 168248 117156
rect 171232 117147 171284 117156
rect 171232 117113 171241 117147
rect 171241 117113 171275 117147
rect 171275 117113 171284 117147
rect 171232 117104 171284 117113
rect 172888 117104 172940 117156
rect 176016 117104 176068 117156
rect 176936 117104 176988 117156
rect 177580 117036 177632 117088
rect 19606 116934 19658 116986
rect 19670 116934 19722 116986
rect 19734 116934 19786 116986
rect 19798 116934 19850 116986
rect 50326 116934 50378 116986
rect 50390 116934 50442 116986
rect 50454 116934 50506 116986
rect 50518 116934 50570 116986
rect 81046 116934 81098 116986
rect 81110 116934 81162 116986
rect 81174 116934 81226 116986
rect 81238 116934 81290 116986
rect 111766 116934 111818 116986
rect 111830 116934 111882 116986
rect 111894 116934 111946 116986
rect 111958 116934 112010 116986
rect 142486 116934 142538 116986
rect 142550 116934 142602 116986
rect 142614 116934 142666 116986
rect 142678 116934 142730 116986
rect 173206 116934 173258 116986
rect 173270 116934 173322 116986
rect 173334 116934 173386 116986
rect 173398 116934 173450 116986
rect 13360 116832 13412 116884
rect 29276 116832 29328 116884
rect 58256 116875 58308 116884
rect 58256 116841 58265 116875
rect 58265 116841 58299 116875
rect 58299 116841 58308 116875
rect 58256 116832 58308 116841
rect 68468 116832 68520 116884
rect 111156 116832 111208 116884
rect 162032 116832 162084 116884
rect 18052 116764 18104 116816
rect 29092 116764 29144 116816
rect 67824 116764 67876 116816
rect 107200 116764 107252 116816
rect 4344 116696 4396 116748
rect 26424 116696 26476 116748
rect 58440 116739 58492 116748
rect 58440 116705 58449 116739
rect 58449 116705 58483 116739
rect 58483 116705 58492 116739
rect 58440 116696 58492 116705
rect 66076 116696 66128 116748
rect 103060 116696 103112 116748
rect 158812 116739 158864 116748
rect 158812 116705 158821 116739
rect 158821 116705 158855 116739
rect 158855 116705 158864 116739
rect 158812 116696 158864 116705
rect 23020 116628 23072 116680
rect 31024 116628 31076 116680
rect 65248 116628 65300 116680
rect 97632 116628 97684 116680
rect 8484 116560 8536 116612
rect 26608 116560 26660 116612
rect 61016 116560 61068 116612
rect 93216 116560 93268 116612
rect 60188 116492 60240 116544
rect 88432 116492 88484 116544
rect 4246 116390 4298 116442
rect 4310 116390 4362 116442
rect 4374 116390 4426 116442
rect 4438 116390 4490 116442
rect 34966 116390 35018 116442
rect 35030 116390 35082 116442
rect 35094 116390 35146 116442
rect 35158 116390 35210 116442
rect 65686 116390 65738 116442
rect 65750 116390 65802 116442
rect 65814 116390 65866 116442
rect 65878 116390 65930 116442
rect 96406 116390 96458 116442
rect 96470 116390 96522 116442
rect 96534 116390 96586 116442
rect 96598 116390 96650 116442
rect 127126 116390 127178 116442
rect 127190 116390 127242 116442
rect 127254 116390 127306 116442
rect 127318 116390 127370 116442
rect 157846 116390 157898 116442
rect 157910 116390 157962 116442
rect 157974 116390 158026 116442
rect 158038 116390 158090 116442
rect 2412 116288 2464 116340
rect 8300 116288 8352 116340
rect 12348 116288 12400 116340
rect 16488 116288 16540 116340
rect 22560 116331 22612 116340
rect 22560 116297 22569 116331
rect 22569 116297 22603 116331
rect 22603 116297 22612 116331
rect 22560 116288 22612 116297
rect 26516 116288 26568 116340
rect 30840 116331 30892 116340
rect 30840 116297 30849 116331
rect 30849 116297 30883 116331
rect 30883 116297 30892 116331
rect 30840 116288 30892 116297
rect 35256 116331 35308 116340
rect 35256 116297 35265 116331
rect 35265 116297 35299 116331
rect 35299 116297 35308 116331
rect 35256 116288 35308 116297
rect 39764 116331 39816 116340
rect 39764 116297 39773 116331
rect 39773 116297 39807 116331
rect 39807 116297 39816 116331
rect 39764 116288 39816 116297
rect 44364 116331 44416 116340
rect 44364 116297 44373 116331
rect 44373 116297 44407 116331
rect 44407 116297 44416 116331
rect 44364 116288 44416 116297
rect 48964 116331 49016 116340
rect 48964 116297 48973 116331
rect 48973 116297 49007 116331
rect 49007 116297 49016 116331
rect 48964 116288 49016 116297
rect 54024 116331 54076 116340
rect 54024 116297 54033 116331
rect 54033 116297 54067 116331
rect 54067 116297 54076 116331
rect 54024 116288 54076 116297
rect 62948 116331 63000 116340
rect 62948 116297 62957 116331
rect 62957 116297 62991 116331
rect 62991 116297 63000 116331
rect 62948 116288 63000 116297
rect 59268 116220 59320 116272
rect 76932 116288 76984 116340
rect 77116 116331 77168 116340
rect 77116 116297 77125 116331
rect 77125 116297 77159 116331
rect 77159 116297 77168 116331
rect 77116 116288 77168 116297
rect 81808 116331 81860 116340
rect 81808 116297 81817 116331
rect 81817 116297 81851 116331
rect 81851 116297 81860 116331
rect 81808 116288 81860 116297
rect 86592 116331 86644 116340
rect 86592 116297 86601 116331
rect 86601 116297 86635 116331
rect 86635 116297 86644 116331
rect 86592 116288 86644 116297
rect 91376 116331 91428 116340
rect 91376 116297 91385 116331
rect 91385 116297 91419 116331
rect 91419 116297 91428 116331
rect 91376 116288 91428 116297
rect 96068 116331 96120 116340
rect 96068 116297 96077 116331
rect 96077 116297 96111 116331
rect 96111 116297 96120 116331
rect 96068 116288 96120 116297
rect 101220 116331 101272 116340
rect 101220 116297 101229 116331
rect 101229 116297 101263 116331
rect 101263 116297 101272 116331
rect 101220 116288 101272 116297
rect 105360 116331 105412 116340
rect 105360 116297 105369 116331
rect 105369 116297 105403 116331
rect 105403 116297 105412 116331
rect 105360 116288 105412 116297
rect 110236 116331 110288 116340
rect 110236 116297 110245 116331
rect 110245 116297 110279 116331
rect 110279 116297 110288 116331
rect 110236 116288 110288 116297
rect 114928 116331 114980 116340
rect 114928 116297 114937 116331
rect 114937 116297 114971 116331
rect 114971 116297 114980 116331
rect 114928 116288 114980 116297
rect 119620 116331 119672 116340
rect 119620 116297 119629 116331
rect 119629 116297 119663 116331
rect 119663 116297 119672 116331
rect 119620 116288 119672 116297
rect 124312 116331 124364 116340
rect 124312 116297 124321 116331
rect 124321 116297 124355 116331
rect 124355 116297 124364 116331
rect 124312 116288 124364 116297
rect 128912 116331 128964 116340
rect 128912 116297 128921 116331
rect 128921 116297 128955 116331
rect 128955 116297 128964 116331
rect 128912 116288 128964 116297
rect 133512 116331 133564 116340
rect 133512 116297 133521 116331
rect 133521 116297 133555 116331
rect 133555 116297 133564 116331
rect 133512 116288 133564 116297
rect 138020 116331 138072 116340
rect 138020 116297 138029 116331
rect 138029 116297 138063 116331
rect 138063 116297 138072 116331
rect 138020 116288 138072 116297
rect 143172 116331 143224 116340
rect 143172 116297 143181 116331
rect 143181 116297 143215 116331
rect 143215 116297 143224 116331
rect 143172 116288 143224 116297
rect 146760 116331 146812 116340
rect 146760 116297 146769 116331
rect 146769 116297 146803 116331
rect 146803 116297 146812 116331
rect 146760 116288 146812 116297
rect 150900 116331 150952 116340
rect 150900 116297 150909 116331
rect 150909 116297 150943 116331
rect 150943 116297 150952 116331
rect 150900 116288 150952 116297
rect 154120 116331 154172 116340
rect 154120 116297 154129 116331
rect 154129 116297 154163 116331
rect 154163 116297 154172 116331
rect 154120 116288 154172 116297
rect 154856 116331 154908 116340
rect 154856 116297 154865 116331
rect 154865 116297 154899 116331
rect 154899 116297 154908 116331
rect 154856 116288 154908 116297
rect 159088 116331 159140 116340
rect 159088 116297 159097 116331
rect 159097 116297 159131 116331
rect 159131 116297 159140 116331
rect 159088 116288 159140 116297
rect 162124 116331 162176 116340
rect 162124 116297 162133 116331
rect 162133 116297 162167 116331
rect 162167 116297 162176 116331
rect 162124 116288 162176 116297
rect 164332 116331 164384 116340
rect 164332 116297 164341 116331
rect 164341 116297 164375 116331
rect 164375 116297 164384 116331
rect 164332 116288 164384 116297
rect 168196 116331 168248 116340
rect 168196 116297 168205 116331
rect 168205 116297 168239 116331
rect 168239 116297 168248 116331
rect 168196 116288 168248 116297
rect 172888 116331 172940 116340
rect 172888 116297 172897 116331
rect 172897 116297 172931 116331
rect 172931 116297 172940 116331
rect 172888 116288 172940 116297
rect 176016 116331 176068 116340
rect 176016 116297 176025 116331
rect 176025 116297 176059 116331
rect 176059 116297 176068 116331
rect 176016 116288 176068 116297
rect 176936 116331 176988 116340
rect 176936 116297 176945 116331
rect 176945 116297 176979 116331
rect 176979 116297 176988 116331
rect 176936 116288 176988 116297
rect 177580 116331 177632 116340
rect 177580 116297 177589 116331
rect 177589 116297 177623 116331
rect 177623 116297 177632 116331
rect 177580 116288 177632 116297
rect 67640 116263 67692 116272
rect 67640 116229 67649 116263
rect 67649 116229 67683 116263
rect 67683 116229 67692 116263
rect 67640 116220 67692 116229
rect 72424 116263 72476 116272
rect 72424 116229 72433 116263
rect 72433 116229 72467 116263
rect 72467 116229 72476 116263
rect 72424 116220 72476 116229
rect 31760 116084 31812 116136
rect 57152 116152 57204 116204
rect 79048 116220 79100 116272
rect 58440 116084 58492 116136
rect 158812 116084 158864 116136
rect 171232 116084 171284 116136
rect 54208 115948 54260 116000
rect 69572 116016 69624 116068
rect 72424 116016 72476 116068
rect 116676 116016 116728 116068
rect 19606 115846 19658 115898
rect 19670 115846 19722 115898
rect 19734 115846 19786 115898
rect 19798 115846 19850 115898
rect 50326 115846 50378 115898
rect 50390 115846 50442 115898
rect 50454 115846 50506 115898
rect 50518 115846 50570 115898
rect 81046 115846 81098 115898
rect 81110 115846 81162 115898
rect 81174 115846 81226 115898
rect 81238 115846 81290 115898
rect 111766 115846 111818 115898
rect 111830 115846 111882 115898
rect 111894 115846 111946 115898
rect 111958 115846 112010 115898
rect 142486 115846 142538 115898
rect 142550 115846 142602 115898
rect 142614 115846 142666 115898
rect 142678 115846 142730 115898
rect 173206 115846 173258 115898
rect 173270 115846 173322 115898
rect 173334 115846 173386 115898
rect 173398 115846 173450 115898
rect 4246 115302 4298 115354
rect 4310 115302 4362 115354
rect 4374 115302 4426 115354
rect 4438 115302 4490 115354
rect 34966 115302 35018 115354
rect 35030 115302 35082 115354
rect 35094 115302 35146 115354
rect 35158 115302 35210 115354
rect 65686 115302 65738 115354
rect 65750 115302 65802 115354
rect 65814 115302 65866 115354
rect 65878 115302 65930 115354
rect 96406 115302 96458 115354
rect 96470 115302 96522 115354
rect 96534 115302 96586 115354
rect 96598 115302 96650 115354
rect 127126 115302 127178 115354
rect 127190 115302 127242 115354
rect 127254 115302 127306 115354
rect 127318 115302 127370 115354
rect 157846 115302 157898 115354
rect 157910 115302 157962 115354
rect 157974 115302 158026 115354
rect 158038 115302 158090 115354
rect 19606 114758 19658 114810
rect 19670 114758 19722 114810
rect 19734 114758 19786 114810
rect 19798 114758 19850 114810
rect 50326 114758 50378 114810
rect 50390 114758 50442 114810
rect 50454 114758 50506 114810
rect 50518 114758 50570 114810
rect 81046 114758 81098 114810
rect 81110 114758 81162 114810
rect 81174 114758 81226 114810
rect 81238 114758 81290 114810
rect 111766 114758 111818 114810
rect 111830 114758 111882 114810
rect 111894 114758 111946 114810
rect 111958 114758 112010 114810
rect 142486 114758 142538 114810
rect 142550 114758 142602 114810
rect 142614 114758 142666 114810
rect 142678 114758 142730 114810
rect 173206 114758 173258 114810
rect 173270 114758 173322 114810
rect 173334 114758 173386 114810
rect 173398 114758 173450 114810
rect 4246 114214 4298 114266
rect 4310 114214 4362 114266
rect 4374 114214 4426 114266
rect 4438 114214 4490 114266
rect 34966 114214 35018 114266
rect 35030 114214 35082 114266
rect 35094 114214 35146 114266
rect 35158 114214 35210 114266
rect 65686 114214 65738 114266
rect 65750 114214 65802 114266
rect 65814 114214 65866 114266
rect 65878 114214 65930 114266
rect 96406 114214 96458 114266
rect 96470 114214 96522 114266
rect 96534 114214 96586 114266
rect 96598 114214 96650 114266
rect 127126 114214 127178 114266
rect 127190 114214 127242 114266
rect 127254 114214 127306 114266
rect 127318 114214 127370 114266
rect 157846 114214 157898 114266
rect 157910 114214 157962 114266
rect 157974 114214 158026 114266
rect 158038 114214 158090 114266
rect 19606 113670 19658 113722
rect 19670 113670 19722 113722
rect 19734 113670 19786 113722
rect 19798 113670 19850 113722
rect 50326 113670 50378 113722
rect 50390 113670 50442 113722
rect 50454 113670 50506 113722
rect 50518 113670 50570 113722
rect 81046 113670 81098 113722
rect 81110 113670 81162 113722
rect 81174 113670 81226 113722
rect 81238 113670 81290 113722
rect 111766 113670 111818 113722
rect 111830 113670 111882 113722
rect 111894 113670 111946 113722
rect 111958 113670 112010 113722
rect 142486 113670 142538 113722
rect 142550 113670 142602 113722
rect 142614 113670 142666 113722
rect 142678 113670 142730 113722
rect 173206 113670 173258 113722
rect 173270 113670 173322 113722
rect 173334 113670 173386 113722
rect 173398 113670 173450 113722
rect 4246 113126 4298 113178
rect 4310 113126 4362 113178
rect 4374 113126 4426 113178
rect 4438 113126 4490 113178
rect 34966 113126 35018 113178
rect 35030 113126 35082 113178
rect 35094 113126 35146 113178
rect 35158 113126 35210 113178
rect 65686 113126 65738 113178
rect 65750 113126 65802 113178
rect 65814 113126 65866 113178
rect 65878 113126 65930 113178
rect 96406 113126 96458 113178
rect 96470 113126 96522 113178
rect 96534 113126 96586 113178
rect 96598 113126 96650 113178
rect 127126 113126 127178 113178
rect 127190 113126 127242 113178
rect 127254 113126 127306 113178
rect 127318 113126 127370 113178
rect 157846 113126 157898 113178
rect 157910 113126 157962 113178
rect 157974 113126 158026 113178
rect 158038 113126 158090 113178
rect 19606 112582 19658 112634
rect 19670 112582 19722 112634
rect 19734 112582 19786 112634
rect 19798 112582 19850 112634
rect 50326 112582 50378 112634
rect 50390 112582 50442 112634
rect 50454 112582 50506 112634
rect 50518 112582 50570 112634
rect 81046 112582 81098 112634
rect 81110 112582 81162 112634
rect 81174 112582 81226 112634
rect 81238 112582 81290 112634
rect 111766 112582 111818 112634
rect 111830 112582 111882 112634
rect 111894 112582 111946 112634
rect 111958 112582 112010 112634
rect 142486 112582 142538 112634
rect 142550 112582 142602 112634
rect 142614 112582 142666 112634
rect 142678 112582 142730 112634
rect 173206 112582 173258 112634
rect 173270 112582 173322 112634
rect 173334 112582 173386 112634
rect 173398 112582 173450 112634
rect 4246 112038 4298 112090
rect 4310 112038 4362 112090
rect 4374 112038 4426 112090
rect 4438 112038 4490 112090
rect 34966 112038 35018 112090
rect 35030 112038 35082 112090
rect 35094 112038 35146 112090
rect 35158 112038 35210 112090
rect 65686 112038 65738 112090
rect 65750 112038 65802 112090
rect 65814 112038 65866 112090
rect 65878 112038 65930 112090
rect 96406 112038 96458 112090
rect 96470 112038 96522 112090
rect 96534 112038 96586 112090
rect 96598 112038 96650 112090
rect 127126 112038 127178 112090
rect 127190 112038 127242 112090
rect 127254 112038 127306 112090
rect 127318 112038 127370 112090
rect 157846 112038 157898 112090
rect 157910 112038 157962 112090
rect 157974 112038 158026 112090
rect 158038 112038 158090 112090
rect 19606 111494 19658 111546
rect 19670 111494 19722 111546
rect 19734 111494 19786 111546
rect 19798 111494 19850 111546
rect 50326 111494 50378 111546
rect 50390 111494 50442 111546
rect 50454 111494 50506 111546
rect 50518 111494 50570 111546
rect 81046 111494 81098 111546
rect 81110 111494 81162 111546
rect 81174 111494 81226 111546
rect 81238 111494 81290 111546
rect 111766 111494 111818 111546
rect 111830 111494 111882 111546
rect 111894 111494 111946 111546
rect 111958 111494 112010 111546
rect 142486 111494 142538 111546
rect 142550 111494 142602 111546
rect 142614 111494 142666 111546
rect 142678 111494 142730 111546
rect 173206 111494 173258 111546
rect 173270 111494 173322 111546
rect 173334 111494 173386 111546
rect 173398 111494 173450 111546
rect 4246 110950 4298 111002
rect 4310 110950 4362 111002
rect 4374 110950 4426 111002
rect 4438 110950 4490 111002
rect 34966 110950 35018 111002
rect 35030 110950 35082 111002
rect 35094 110950 35146 111002
rect 35158 110950 35210 111002
rect 65686 110950 65738 111002
rect 65750 110950 65802 111002
rect 65814 110950 65866 111002
rect 65878 110950 65930 111002
rect 96406 110950 96458 111002
rect 96470 110950 96522 111002
rect 96534 110950 96586 111002
rect 96598 110950 96650 111002
rect 127126 110950 127178 111002
rect 127190 110950 127242 111002
rect 127254 110950 127306 111002
rect 127318 110950 127370 111002
rect 157846 110950 157898 111002
rect 157910 110950 157962 111002
rect 157974 110950 158026 111002
rect 158038 110950 158090 111002
rect 19606 110406 19658 110458
rect 19670 110406 19722 110458
rect 19734 110406 19786 110458
rect 19798 110406 19850 110458
rect 50326 110406 50378 110458
rect 50390 110406 50442 110458
rect 50454 110406 50506 110458
rect 50518 110406 50570 110458
rect 81046 110406 81098 110458
rect 81110 110406 81162 110458
rect 81174 110406 81226 110458
rect 81238 110406 81290 110458
rect 111766 110406 111818 110458
rect 111830 110406 111882 110458
rect 111894 110406 111946 110458
rect 111958 110406 112010 110458
rect 142486 110406 142538 110458
rect 142550 110406 142602 110458
rect 142614 110406 142666 110458
rect 142678 110406 142730 110458
rect 173206 110406 173258 110458
rect 173270 110406 173322 110458
rect 173334 110406 173386 110458
rect 173398 110406 173450 110458
rect 4246 109862 4298 109914
rect 4310 109862 4362 109914
rect 4374 109862 4426 109914
rect 4438 109862 4490 109914
rect 34966 109862 35018 109914
rect 35030 109862 35082 109914
rect 35094 109862 35146 109914
rect 35158 109862 35210 109914
rect 65686 109862 65738 109914
rect 65750 109862 65802 109914
rect 65814 109862 65866 109914
rect 65878 109862 65930 109914
rect 96406 109862 96458 109914
rect 96470 109862 96522 109914
rect 96534 109862 96586 109914
rect 96598 109862 96650 109914
rect 127126 109862 127178 109914
rect 127190 109862 127242 109914
rect 127254 109862 127306 109914
rect 127318 109862 127370 109914
rect 157846 109862 157898 109914
rect 157910 109862 157962 109914
rect 157974 109862 158026 109914
rect 158038 109862 158090 109914
rect 19606 109318 19658 109370
rect 19670 109318 19722 109370
rect 19734 109318 19786 109370
rect 19798 109318 19850 109370
rect 50326 109318 50378 109370
rect 50390 109318 50442 109370
rect 50454 109318 50506 109370
rect 50518 109318 50570 109370
rect 81046 109318 81098 109370
rect 81110 109318 81162 109370
rect 81174 109318 81226 109370
rect 81238 109318 81290 109370
rect 111766 109318 111818 109370
rect 111830 109318 111882 109370
rect 111894 109318 111946 109370
rect 111958 109318 112010 109370
rect 142486 109318 142538 109370
rect 142550 109318 142602 109370
rect 142614 109318 142666 109370
rect 142678 109318 142730 109370
rect 173206 109318 173258 109370
rect 173270 109318 173322 109370
rect 173334 109318 173386 109370
rect 173398 109318 173450 109370
rect 4246 108774 4298 108826
rect 4310 108774 4362 108826
rect 4374 108774 4426 108826
rect 4438 108774 4490 108826
rect 34966 108774 35018 108826
rect 35030 108774 35082 108826
rect 35094 108774 35146 108826
rect 35158 108774 35210 108826
rect 65686 108774 65738 108826
rect 65750 108774 65802 108826
rect 65814 108774 65866 108826
rect 65878 108774 65930 108826
rect 96406 108774 96458 108826
rect 96470 108774 96522 108826
rect 96534 108774 96586 108826
rect 96598 108774 96650 108826
rect 127126 108774 127178 108826
rect 127190 108774 127242 108826
rect 127254 108774 127306 108826
rect 127318 108774 127370 108826
rect 157846 108774 157898 108826
rect 157910 108774 157962 108826
rect 157974 108774 158026 108826
rect 158038 108774 158090 108826
rect 19606 108230 19658 108282
rect 19670 108230 19722 108282
rect 19734 108230 19786 108282
rect 19798 108230 19850 108282
rect 50326 108230 50378 108282
rect 50390 108230 50442 108282
rect 50454 108230 50506 108282
rect 50518 108230 50570 108282
rect 81046 108230 81098 108282
rect 81110 108230 81162 108282
rect 81174 108230 81226 108282
rect 81238 108230 81290 108282
rect 111766 108230 111818 108282
rect 111830 108230 111882 108282
rect 111894 108230 111946 108282
rect 111958 108230 112010 108282
rect 142486 108230 142538 108282
rect 142550 108230 142602 108282
rect 142614 108230 142666 108282
rect 142678 108230 142730 108282
rect 173206 108230 173258 108282
rect 173270 108230 173322 108282
rect 173334 108230 173386 108282
rect 173398 108230 173450 108282
rect 4246 107686 4298 107738
rect 4310 107686 4362 107738
rect 4374 107686 4426 107738
rect 4438 107686 4490 107738
rect 34966 107686 35018 107738
rect 35030 107686 35082 107738
rect 35094 107686 35146 107738
rect 35158 107686 35210 107738
rect 65686 107686 65738 107738
rect 65750 107686 65802 107738
rect 65814 107686 65866 107738
rect 65878 107686 65930 107738
rect 96406 107686 96458 107738
rect 96470 107686 96522 107738
rect 96534 107686 96586 107738
rect 96598 107686 96650 107738
rect 127126 107686 127178 107738
rect 127190 107686 127242 107738
rect 127254 107686 127306 107738
rect 127318 107686 127370 107738
rect 157846 107686 157898 107738
rect 157910 107686 157962 107738
rect 157974 107686 158026 107738
rect 158038 107686 158090 107738
rect 19606 107142 19658 107194
rect 19670 107142 19722 107194
rect 19734 107142 19786 107194
rect 19798 107142 19850 107194
rect 50326 107142 50378 107194
rect 50390 107142 50442 107194
rect 50454 107142 50506 107194
rect 50518 107142 50570 107194
rect 81046 107142 81098 107194
rect 81110 107142 81162 107194
rect 81174 107142 81226 107194
rect 81238 107142 81290 107194
rect 111766 107142 111818 107194
rect 111830 107142 111882 107194
rect 111894 107142 111946 107194
rect 111958 107142 112010 107194
rect 142486 107142 142538 107194
rect 142550 107142 142602 107194
rect 142614 107142 142666 107194
rect 142678 107142 142730 107194
rect 173206 107142 173258 107194
rect 173270 107142 173322 107194
rect 173334 107142 173386 107194
rect 173398 107142 173450 107194
rect 4246 106598 4298 106650
rect 4310 106598 4362 106650
rect 4374 106598 4426 106650
rect 4438 106598 4490 106650
rect 34966 106598 35018 106650
rect 35030 106598 35082 106650
rect 35094 106598 35146 106650
rect 35158 106598 35210 106650
rect 65686 106598 65738 106650
rect 65750 106598 65802 106650
rect 65814 106598 65866 106650
rect 65878 106598 65930 106650
rect 96406 106598 96458 106650
rect 96470 106598 96522 106650
rect 96534 106598 96586 106650
rect 96598 106598 96650 106650
rect 127126 106598 127178 106650
rect 127190 106598 127242 106650
rect 127254 106598 127306 106650
rect 127318 106598 127370 106650
rect 157846 106598 157898 106650
rect 157910 106598 157962 106650
rect 157974 106598 158026 106650
rect 158038 106598 158090 106650
rect 19606 106054 19658 106106
rect 19670 106054 19722 106106
rect 19734 106054 19786 106106
rect 19798 106054 19850 106106
rect 50326 106054 50378 106106
rect 50390 106054 50442 106106
rect 50454 106054 50506 106106
rect 50518 106054 50570 106106
rect 81046 106054 81098 106106
rect 81110 106054 81162 106106
rect 81174 106054 81226 106106
rect 81238 106054 81290 106106
rect 111766 106054 111818 106106
rect 111830 106054 111882 106106
rect 111894 106054 111946 106106
rect 111958 106054 112010 106106
rect 142486 106054 142538 106106
rect 142550 106054 142602 106106
rect 142614 106054 142666 106106
rect 142678 106054 142730 106106
rect 173206 106054 173258 106106
rect 173270 106054 173322 106106
rect 173334 106054 173386 106106
rect 173398 106054 173450 106106
rect 4246 105510 4298 105562
rect 4310 105510 4362 105562
rect 4374 105510 4426 105562
rect 4438 105510 4490 105562
rect 34966 105510 35018 105562
rect 35030 105510 35082 105562
rect 35094 105510 35146 105562
rect 35158 105510 35210 105562
rect 65686 105510 65738 105562
rect 65750 105510 65802 105562
rect 65814 105510 65866 105562
rect 65878 105510 65930 105562
rect 96406 105510 96458 105562
rect 96470 105510 96522 105562
rect 96534 105510 96586 105562
rect 96598 105510 96650 105562
rect 127126 105510 127178 105562
rect 127190 105510 127242 105562
rect 127254 105510 127306 105562
rect 127318 105510 127370 105562
rect 157846 105510 157898 105562
rect 157910 105510 157962 105562
rect 157974 105510 158026 105562
rect 158038 105510 158090 105562
rect 19606 104966 19658 105018
rect 19670 104966 19722 105018
rect 19734 104966 19786 105018
rect 19798 104966 19850 105018
rect 50326 104966 50378 105018
rect 50390 104966 50442 105018
rect 50454 104966 50506 105018
rect 50518 104966 50570 105018
rect 81046 104966 81098 105018
rect 81110 104966 81162 105018
rect 81174 104966 81226 105018
rect 81238 104966 81290 105018
rect 111766 104966 111818 105018
rect 111830 104966 111882 105018
rect 111894 104966 111946 105018
rect 111958 104966 112010 105018
rect 142486 104966 142538 105018
rect 142550 104966 142602 105018
rect 142614 104966 142666 105018
rect 142678 104966 142730 105018
rect 173206 104966 173258 105018
rect 173270 104966 173322 105018
rect 173334 104966 173386 105018
rect 173398 104966 173450 105018
rect 4246 104422 4298 104474
rect 4310 104422 4362 104474
rect 4374 104422 4426 104474
rect 4438 104422 4490 104474
rect 34966 104422 35018 104474
rect 35030 104422 35082 104474
rect 35094 104422 35146 104474
rect 35158 104422 35210 104474
rect 65686 104422 65738 104474
rect 65750 104422 65802 104474
rect 65814 104422 65866 104474
rect 65878 104422 65930 104474
rect 96406 104422 96458 104474
rect 96470 104422 96522 104474
rect 96534 104422 96586 104474
rect 96598 104422 96650 104474
rect 127126 104422 127178 104474
rect 127190 104422 127242 104474
rect 127254 104422 127306 104474
rect 127318 104422 127370 104474
rect 157846 104422 157898 104474
rect 157910 104422 157962 104474
rect 157974 104422 158026 104474
rect 158038 104422 158090 104474
rect 19606 103878 19658 103930
rect 19670 103878 19722 103930
rect 19734 103878 19786 103930
rect 19798 103878 19850 103930
rect 50326 103878 50378 103930
rect 50390 103878 50442 103930
rect 50454 103878 50506 103930
rect 50518 103878 50570 103930
rect 81046 103878 81098 103930
rect 81110 103878 81162 103930
rect 81174 103878 81226 103930
rect 81238 103878 81290 103930
rect 111766 103878 111818 103930
rect 111830 103878 111882 103930
rect 111894 103878 111946 103930
rect 111958 103878 112010 103930
rect 142486 103878 142538 103930
rect 142550 103878 142602 103930
rect 142614 103878 142666 103930
rect 142678 103878 142730 103930
rect 173206 103878 173258 103930
rect 173270 103878 173322 103930
rect 173334 103878 173386 103930
rect 173398 103878 173450 103930
rect 4246 103334 4298 103386
rect 4310 103334 4362 103386
rect 4374 103334 4426 103386
rect 4438 103334 4490 103386
rect 34966 103334 35018 103386
rect 35030 103334 35082 103386
rect 35094 103334 35146 103386
rect 35158 103334 35210 103386
rect 65686 103334 65738 103386
rect 65750 103334 65802 103386
rect 65814 103334 65866 103386
rect 65878 103334 65930 103386
rect 96406 103334 96458 103386
rect 96470 103334 96522 103386
rect 96534 103334 96586 103386
rect 96598 103334 96650 103386
rect 127126 103334 127178 103386
rect 127190 103334 127242 103386
rect 127254 103334 127306 103386
rect 127318 103334 127370 103386
rect 157846 103334 157898 103386
rect 157910 103334 157962 103386
rect 157974 103334 158026 103386
rect 158038 103334 158090 103386
rect 19606 102790 19658 102842
rect 19670 102790 19722 102842
rect 19734 102790 19786 102842
rect 19798 102790 19850 102842
rect 50326 102790 50378 102842
rect 50390 102790 50442 102842
rect 50454 102790 50506 102842
rect 50518 102790 50570 102842
rect 81046 102790 81098 102842
rect 81110 102790 81162 102842
rect 81174 102790 81226 102842
rect 81238 102790 81290 102842
rect 111766 102790 111818 102842
rect 111830 102790 111882 102842
rect 111894 102790 111946 102842
rect 111958 102790 112010 102842
rect 142486 102790 142538 102842
rect 142550 102790 142602 102842
rect 142614 102790 142666 102842
rect 142678 102790 142730 102842
rect 173206 102790 173258 102842
rect 173270 102790 173322 102842
rect 173334 102790 173386 102842
rect 173398 102790 173450 102842
rect 4246 102246 4298 102298
rect 4310 102246 4362 102298
rect 4374 102246 4426 102298
rect 4438 102246 4490 102298
rect 34966 102246 35018 102298
rect 35030 102246 35082 102298
rect 35094 102246 35146 102298
rect 35158 102246 35210 102298
rect 65686 102246 65738 102298
rect 65750 102246 65802 102298
rect 65814 102246 65866 102298
rect 65878 102246 65930 102298
rect 96406 102246 96458 102298
rect 96470 102246 96522 102298
rect 96534 102246 96586 102298
rect 96598 102246 96650 102298
rect 127126 102246 127178 102298
rect 127190 102246 127242 102298
rect 127254 102246 127306 102298
rect 127318 102246 127370 102298
rect 157846 102246 157898 102298
rect 157910 102246 157962 102298
rect 157974 102246 158026 102298
rect 158038 102246 158090 102298
rect 19606 101702 19658 101754
rect 19670 101702 19722 101754
rect 19734 101702 19786 101754
rect 19798 101702 19850 101754
rect 50326 101702 50378 101754
rect 50390 101702 50442 101754
rect 50454 101702 50506 101754
rect 50518 101702 50570 101754
rect 81046 101702 81098 101754
rect 81110 101702 81162 101754
rect 81174 101702 81226 101754
rect 81238 101702 81290 101754
rect 111766 101702 111818 101754
rect 111830 101702 111882 101754
rect 111894 101702 111946 101754
rect 111958 101702 112010 101754
rect 142486 101702 142538 101754
rect 142550 101702 142602 101754
rect 142614 101702 142666 101754
rect 142678 101702 142730 101754
rect 173206 101702 173258 101754
rect 173270 101702 173322 101754
rect 173334 101702 173386 101754
rect 173398 101702 173450 101754
rect 4246 101158 4298 101210
rect 4310 101158 4362 101210
rect 4374 101158 4426 101210
rect 4438 101158 4490 101210
rect 34966 101158 35018 101210
rect 35030 101158 35082 101210
rect 35094 101158 35146 101210
rect 35158 101158 35210 101210
rect 65686 101158 65738 101210
rect 65750 101158 65802 101210
rect 65814 101158 65866 101210
rect 65878 101158 65930 101210
rect 96406 101158 96458 101210
rect 96470 101158 96522 101210
rect 96534 101158 96586 101210
rect 96598 101158 96650 101210
rect 127126 101158 127178 101210
rect 127190 101158 127242 101210
rect 127254 101158 127306 101210
rect 127318 101158 127370 101210
rect 157846 101158 157898 101210
rect 157910 101158 157962 101210
rect 157974 101158 158026 101210
rect 158038 101158 158090 101210
rect 19606 100614 19658 100666
rect 19670 100614 19722 100666
rect 19734 100614 19786 100666
rect 19798 100614 19850 100666
rect 50326 100614 50378 100666
rect 50390 100614 50442 100666
rect 50454 100614 50506 100666
rect 50518 100614 50570 100666
rect 81046 100614 81098 100666
rect 81110 100614 81162 100666
rect 81174 100614 81226 100666
rect 81238 100614 81290 100666
rect 111766 100614 111818 100666
rect 111830 100614 111882 100666
rect 111894 100614 111946 100666
rect 111958 100614 112010 100666
rect 142486 100614 142538 100666
rect 142550 100614 142602 100666
rect 142614 100614 142666 100666
rect 142678 100614 142730 100666
rect 173206 100614 173258 100666
rect 173270 100614 173322 100666
rect 173334 100614 173386 100666
rect 173398 100614 173450 100666
rect 4246 100070 4298 100122
rect 4310 100070 4362 100122
rect 4374 100070 4426 100122
rect 4438 100070 4490 100122
rect 34966 100070 35018 100122
rect 35030 100070 35082 100122
rect 35094 100070 35146 100122
rect 35158 100070 35210 100122
rect 65686 100070 65738 100122
rect 65750 100070 65802 100122
rect 65814 100070 65866 100122
rect 65878 100070 65930 100122
rect 96406 100070 96458 100122
rect 96470 100070 96522 100122
rect 96534 100070 96586 100122
rect 96598 100070 96650 100122
rect 127126 100070 127178 100122
rect 127190 100070 127242 100122
rect 127254 100070 127306 100122
rect 127318 100070 127370 100122
rect 157846 100070 157898 100122
rect 157910 100070 157962 100122
rect 157974 100070 158026 100122
rect 158038 100070 158090 100122
rect 19606 99526 19658 99578
rect 19670 99526 19722 99578
rect 19734 99526 19786 99578
rect 19798 99526 19850 99578
rect 50326 99526 50378 99578
rect 50390 99526 50442 99578
rect 50454 99526 50506 99578
rect 50518 99526 50570 99578
rect 81046 99526 81098 99578
rect 81110 99526 81162 99578
rect 81174 99526 81226 99578
rect 81238 99526 81290 99578
rect 111766 99526 111818 99578
rect 111830 99526 111882 99578
rect 111894 99526 111946 99578
rect 111958 99526 112010 99578
rect 142486 99526 142538 99578
rect 142550 99526 142602 99578
rect 142614 99526 142666 99578
rect 142678 99526 142730 99578
rect 173206 99526 173258 99578
rect 173270 99526 173322 99578
rect 173334 99526 173386 99578
rect 173398 99526 173450 99578
rect 4246 98982 4298 99034
rect 4310 98982 4362 99034
rect 4374 98982 4426 99034
rect 4438 98982 4490 99034
rect 34966 98982 35018 99034
rect 35030 98982 35082 99034
rect 35094 98982 35146 99034
rect 35158 98982 35210 99034
rect 65686 98982 65738 99034
rect 65750 98982 65802 99034
rect 65814 98982 65866 99034
rect 65878 98982 65930 99034
rect 96406 98982 96458 99034
rect 96470 98982 96522 99034
rect 96534 98982 96586 99034
rect 96598 98982 96650 99034
rect 127126 98982 127178 99034
rect 127190 98982 127242 99034
rect 127254 98982 127306 99034
rect 127318 98982 127370 99034
rect 157846 98982 157898 99034
rect 157910 98982 157962 99034
rect 157974 98982 158026 99034
rect 158038 98982 158090 99034
rect 19606 98438 19658 98490
rect 19670 98438 19722 98490
rect 19734 98438 19786 98490
rect 19798 98438 19850 98490
rect 50326 98438 50378 98490
rect 50390 98438 50442 98490
rect 50454 98438 50506 98490
rect 50518 98438 50570 98490
rect 81046 98438 81098 98490
rect 81110 98438 81162 98490
rect 81174 98438 81226 98490
rect 81238 98438 81290 98490
rect 111766 98438 111818 98490
rect 111830 98438 111882 98490
rect 111894 98438 111946 98490
rect 111958 98438 112010 98490
rect 142486 98438 142538 98490
rect 142550 98438 142602 98490
rect 142614 98438 142666 98490
rect 142678 98438 142730 98490
rect 173206 98438 173258 98490
rect 173270 98438 173322 98490
rect 173334 98438 173386 98490
rect 173398 98438 173450 98490
rect 4246 97894 4298 97946
rect 4310 97894 4362 97946
rect 4374 97894 4426 97946
rect 4438 97894 4490 97946
rect 34966 97894 35018 97946
rect 35030 97894 35082 97946
rect 35094 97894 35146 97946
rect 35158 97894 35210 97946
rect 65686 97894 65738 97946
rect 65750 97894 65802 97946
rect 65814 97894 65866 97946
rect 65878 97894 65930 97946
rect 96406 97894 96458 97946
rect 96470 97894 96522 97946
rect 96534 97894 96586 97946
rect 96598 97894 96650 97946
rect 127126 97894 127178 97946
rect 127190 97894 127242 97946
rect 127254 97894 127306 97946
rect 127318 97894 127370 97946
rect 157846 97894 157898 97946
rect 157910 97894 157962 97946
rect 157974 97894 158026 97946
rect 158038 97894 158090 97946
rect 19606 97350 19658 97402
rect 19670 97350 19722 97402
rect 19734 97350 19786 97402
rect 19798 97350 19850 97402
rect 50326 97350 50378 97402
rect 50390 97350 50442 97402
rect 50454 97350 50506 97402
rect 50518 97350 50570 97402
rect 81046 97350 81098 97402
rect 81110 97350 81162 97402
rect 81174 97350 81226 97402
rect 81238 97350 81290 97402
rect 111766 97350 111818 97402
rect 111830 97350 111882 97402
rect 111894 97350 111946 97402
rect 111958 97350 112010 97402
rect 142486 97350 142538 97402
rect 142550 97350 142602 97402
rect 142614 97350 142666 97402
rect 142678 97350 142730 97402
rect 173206 97350 173258 97402
rect 173270 97350 173322 97402
rect 173334 97350 173386 97402
rect 173398 97350 173450 97402
rect 4246 96806 4298 96858
rect 4310 96806 4362 96858
rect 4374 96806 4426 96858
rect 4438 96806 4490 96858
rect 34966 96806 35018 96858
rect 35030 96806 35082 96858
rect 35094 96806 35146 96858
rect 35158 96806 35210 96858
rect 65686 96806 65738 96858
rect 65750 96806 65802 96858
rect 65814 96806 65866 96858
rect 65878 96806 65930 96858
rect 96406 96806 96458 96858
rect 96470 96806 96522 96858
rect 96534 96806 96586 96858
rect 96598 96806 96650 96858
rect 127126 96806 127178 96858
rect 127190 96806 127242 96858
rect 127254 96806 127306 96858
rect 127318 96806 127370 96858
rect 157846 96806 157898 96858
rect 157910 96806 157962 96858
rect 157974 96806 158026 96858
rect 158038 96806 158090 96858
rect 19606 96262 19658 96314
rect 19670 96262 19722 96314
rect 19734 96262 19786 96314
rect 19798 96262 19850 96314
rect 50326 96262 50378 96314
rect 50390 96262 50442 96314
rect 50454 96262 50506 96314
rect 50518 96262 50570 96314
rect 81046 96262 81098 96314
rect 81110 96262 81162 96314
rect 81174 96262 81226 96314
rect 81238 96262 81290 96314
rect 111766 96262 111818 96314
rect 111830 96262 111882 96314
rect 111894 96262 111946 96314
rect 111958 96262 112010 96314
rect 142486 96262 142538 96314
rect 142550 96262 142602 96314
rect 142614 96262 142666 96314
rect 142678 96262 142730 96314
rect 173206 96262 173258 96314
rect 173270 96262 173322 96314
rect 173334 96262 173386 96314
rect 173398 96262 173450 96314
rect 4246 95718 4298 95770
rect 4310 95718 4362 95770
rect 4374 95718 4426 95770
rect 4438 95718 4490 95770
rect 34966 95718 35018 95770
rect 35030 95718 35082 95770
rect 35094 95718 35146 95770
rect 35158 95718 35210 95770
rect 65686 95718 65738 95770
rect 65750 95718 65802 95770
rect 65814 95718 65866 95770
rect 65878 95718 65930 95770
rect 96406 95718 96458 95770
rect 96470 95718 96522 95770
rect 96534 95718 96586 95770
rect 96598 95718 96650 95770
rect 127126 95718 127178 95770
rect 127190 95718 127242 95770
rect 127254 95718 127306 95770
rect 127318 95718 127370 95770
rect 157846 95718 157898 95770
rect 157910 95718 157962 95770
rect 157974 95718 158026 95770
rect 158038 95718 158090 95770
rect 19606 95174 19658 95226
rect 19670 95174 19722 95226
rect 19734 95174 19786 95226
rect 19798 95174 19850 95226
rect 50326 95174 50378 95226
rect 50390 95174 50442 95226
rect 50454 95174 50506 95226
rect 50518 95174 50570 95226
rect 81046 95174 81098 95226
rect 81110 95174 81162 95226
rect 81174 95174 81226 95226
rect 81238 95174 81290 95226
rect 111766 95174 111818 95226
rect 111830 95174 111882 95226
rect 111894 95174 111946 95226
rect 111958 95174 112010 95226
rect 142486 95174 142538 95226
rect 142550 95174 142602 95226
rect 142614 95174 142666 95226
rect 142678 95174 142730 95226
rect 173206 95174 173258 95226
rect 173270 95174 173322 95226
rect 173334 95174 173386 95226
rect 173398 95174 173450 95226
rect 4246 94630 4298 94682
rect 4310 94630 4362 94682
rect 4374 94630 4426 94682
rect 4438 94630 4490 94682
rect 34966 94630 35018 94682
rect 35030 94630 35082 94682
rect 35094 94630 35146 94682
rect 35158 94630 35210 94682
rect 65686 94630 65738 94682
rect 65750 94630 65802 94682
rect 65814 94630 65866 94682
rect 65878 94630 65930 94682
rect 96406 94630 96458 94682
rect 96470 94630 96522 94682
rect 96534 94630 96586 94682
rect 96598 94630 96650 94682
rect 127126 94630 127178 94682
rect 127190 94630 127242 94682
rect 127254 94630 127306 94682
rect 127318 94630 127370 94682
rect 157846 94630 157898 94682
rect 157910 94630 157962 94682
rect 157974 94630 158026 94682
rect 158038 94630 158090 94682
rect 19606 94086 19658 94138
rect 19670 94086 19722 94138
rect 19734 94086 19786 94138
rect 19798 94086 19850 94138
rect 50326 94086 50378 94138
rect 50390 94086 50442 94138
rect 50454 94086 50506 94138
rect 50518 94086 50570 94138
rect 81046 94086 81098 94138
rect 81110 94086 81162 94138
rect 81174 94086 81226 94138
rect 81238 94086 81290 94138
rect 111766 94086 111818 94138
rect 111830 94086 111882 94138
rect 111894 94086 111946 94138
rect 111958 94086 112010 94138
rect 142486 94086 142538 94138
rect 142550 94086 142602 94138
rect 142614 94086 142666 94138
rect 142678 94086 142730 94138
rect 173206 94086 173258 94138
rect 173270 94086 173322 94138
rect 173334 94086 173386 94138
rect 173398 94086 173450 94138
rect 4246 93542 4298 93594
rect 4310 93542 4362 93594
rect 4374 93542 4426 93594
rect 4438 93542 4490 93594
rect 34966 93542 35018 93594
rect 35030 93542 35082 93594
rect 35094 93542 35146 93594
rect 35158 93542 35210 93594
rect 65686 93542 65738 93594
rect 65750 93542 65802 93594
rect 65814 93542 65866 93594
rect 65878 93542 65930 93594
rect 96406 93542 96458 93594
rect 96470 93542 96522 93594
rect 96534 93542 96586 93594
rect 96598 93542 96650 93594
rect 127126 93542 127178 93594
rect 127190 93542 127242 93594
rect 127254 93542 127306 93594
rect 127318 93542 127370 93594
rect 157846 93542 157898 93594
rect 157910 93542 157962 93594
rect 157974 93542 158026 93594
rect 158038 93542 158090 93594
rect 19606 92998 19658 93050
rect 19670 92998 19722 93050
rect 19734 92998 19786 93050
rect 19798 92998 19850 93050
rect 50326 92998 50378 93050
rect 50390 92998 50442 93050
rect 50454 92998 50506 93050
rect 50518 92998 50570 93050
rect 81046 92998 81098 93050
rect 81110 92998 81162 93050
rect 81174 92998 81226 93050
rect 81238 92998 81290 93050
rect 111766 92998 111818 93050
rect 111830 92998 111882 93050
rect 111894 92998 111946 93050
rect 111958 92998 112010 93050
rect 142486 92998 142538 93050
rect 142550 92998 142602 93050
rect 142614 92998 142666 93050
rect 142678 92998 142730 93050
rect 173206 92998 173258 93050
rect 173270 92998 173322 93050
rect 173334 92998 173386 93050
rect 173398 92998 173450 93050
rect 4246 92454 4298 92506
rect 4310 92454 4362 92506
rect 4374 92454 4426 92506
rect 4438 92454 4490 92506
rect 34966 92454 35018 92506
rect 35030 92454 35082 92506
rect 35094 92454 35146 92506
rect 35158 92454 35210 92506
rect 65686 92454 65738 92506
rect 65750 92454 65802 92506
rect 65814 92454 65866 92506
rect 65878 92454 65930 92506
rect 96406 92454 96458 92506
rect 96470 92454 96522 92506
rect 96534 92454 96586 92506
rect 96598 92454 96650 92506
rect 127126 92454 127178 92506
rect 127190 92454 127242 92506
rect 127254 92454 127306 92506
rect 127318 92454 127370 92506
rect 157846 92454 157898 92506
rect 157910 92454 157962 92506
rect 157974 92454 158026 92506
rect 158038 92454 158090 92506
rect 19606 91910 19658 91962
rect 19670 91910 19722 91962
rect 19734 91910 19786 91962
rect 19798 91910 19850 91962
rect 50326 91910 50378 91962
rect 50390 91910 50442 91962
rect 50454 91910 50506 91962
rect 50518 91910 50570 91962
rect 81046 91910 81098 91962
rect 81110 91910 81162 91962
rect 81174 91910 81226 91962
rect 81238 91910 81290 91962
rect 111766 91910 111818 91962
rect 111830 91910 111882 91962
rect 111894 91910 111946 91962
rect 111958 91910 112010 91962
rect 142486 91910 142538 91962
rect 142550 91910 142602 91962
rect 142614 91910 142666 91962
rect 142678 91910 142730 91962
rect 173206 91910 173258 91962
rect 173270 91910 173322 91962
rect 173334 91910 173386 91962
rect 173398 91910 173450 91962
rect 4246 91366 4298 91418
rect 4310 91366 4362 91418
rect 4374 91366 4426 91418
rect 4438 91366 4490 91418
rect 34966 91366 35018 91418
rect 35030 91366 35082 91418
rect 35094 91366 35146 91418
rect 35158 91366 35210 91418
rect 65686 91366 65738 91418
rect 65750 91366 65802 91418
rect 65814 91366 65866 91418
rect 65878 91366 65930 91418
rect 96406 91366 96458 91418
rect 96470 91366 96522 91418
rect 96534 91366 96586 91418
rect 96598 91366 96650 91418
rect 127126 91366 127178 91418
rect 127190 91366 127242 91418
rect 127254 91366 127306 91418
rect 127318 91366 127370 91418
rect 157846 91366 157898 91418
rect 157910 91366 157962 91418
rect 157974 91366 158026 91418
rect 158038 91366 158090 91418
rect 19606 90822 19658 90874
rect 19670 90822 19722 90874
rect 19734 90822 19786 90874
rect 19798 90822 19850 90874
rect 50326 90822 50378 90874
rect 50390 90822 50442 90874
rect 50454 90822 50506 90874
rect 50518 90822 50570 90874
rect 81046 90822 81098 90874
rect 81110 90822 81162 90874
rect 81174 90822 81226 90874
rect 81238 90822 81290 90874
rect 111766 90822 111818 90874
rect 111830 90822 111882 90874
rect 111894 90822 111946 90874
rect 111958 90822 112010 90874
rect 142486 90822 142538 90874
rect 142550 90822 142602 90874
rect 142614 90822 142666 90874
rect 142678 90822 142730 90874
rect 173206 90822 173258 90874
rect 173270 90822 173322 90874
rect 173334 90822 173386 90874
rect 173398 90822 173450 90874
rect 4246 90278 4298 90330
rect 4310 90278 4362 90330
rect 4374 90278 4426 90330
rect 4438 90278 4490 90330
rect 34966 90278 35018 90330
rect 35030 90278 35082 90330
rect 35094 90278 35146 90330
rect 35158 90278 35210 90330
rect 65686 90278 65738 90330
rect 65750 90278 65802 90330
rect 65814 90278 65866 90330
rect 65878 90278 65930 90330
rect 96406 90278 96458 90330
rect 96470 90278 96522 90330
rect 96534 90278 96586 90330
rect 96598 90278 96650 90330
rect 127126 90278 127178 90330
rect 127190 90278 127242 90330
rect 127254 90278 127306 90330
rect 127318 90278 127370 90330
rect 157846 90278 157898 90330
rect 157910 90278 157962 90330
rect 157974 90278 158026 90330
rect 158038 90278 158090 90330
rect 19606 89734 19658 89786
rect 19670 89734 19722 89786
rect 19734 89734 19786 89786
rect 19798 89734 19850 89786
rect 50326 89734 50378 89786
rect 50390 89734 50442 89786
rect 50454 89734 50506 89786
rect 50518 89734 50570 89786
rect 81046 89734 81098 89786
rect 81110 89734 81162 89786
rect 81174 89734 81226 89786
rect 81238 89734 81290 89786
rect 111766 89734 111818 89786
rect 111830 89734 111882 89786
rect 111894 89734 111946 89786
rect 111958 89734 112010 89786
rect 142486 89734 142538 89786
rect 142550 89734 142602 89786
rect 142614 89734 142666 89786
rect 142678 89734 142730 89786
rect 173206 89734 173258 89786
rect 173270 89734 173322 89786
rect 173334 89734 173386 89786
rect 173398 89734 173450 89786
rect 4246 89190 4298 89242
rect 4310 89190 4362 89242
rect 4374 89190 4426 89242
rect 4438 89190 4490 89242
rect 34966 89190 35018 89242
rect 35030 89190 35082 89242
rect 35094 89190 35146 89242
rect 35158 89190 35210 89242
rect 65686 89190 65738 89242
rect 65750 89190 65802 89242
rect 65814 89190 65866 89242
rect 65878 89190 65930 89242
rect 96406 89190 96458 89242
rect 96470 89190 96522 89242
rect 96534 89190 96586 89242
rect 96598 89190 96650 89242
rect 127126 89190 127178 89242
rect 127190 89190 127242 89242
rect 127254 89190 127306 89242
rect 127318 89190 127370 89242
rect 157846 89190 157898 89242
rect 157910 89190 157962 89242
rect 157974 89190 158026 89242
rect 158038 89190 158090 89242
rect 19606 88646 19658 88698
rect 19670 88646 19722 88698
rect 19734 88646 19786 88698
rect 19798 88646 19850 88698
rect 50326 88646 50378 88698
rect 50390 88646 50442 88698
rect 50454 88646 50506 88698
rect 50518 88646 50570 88698
rect 81046 88646 81098 88698
rect 81110 88646 81162 88698
rect 81174 88646 81226 88698
rect 81238 88646 81290 88698
rect 111766 88646 111818 88698
rect 111830 88646 111882 88698
rect 111894 88646 111946 88698
rect 111958 88646 112010 88698
rect 142486 88646 142538 88698
rect 142550 88646 142602 88698
rect 142614 88646 142666 88698
rect 142678 88646 142730 88698
rect 173206 88646 173258 88698
rect 173270 88646 173322 88698
rect 173334 88646 173386 88698
rect 173398 88646 173450 88698
rect 4246 88102 4298 88154
rect 4310 88102 4362 88154
rect 4374 88102 4426 88154
rect 4438 88102 4490 88154
rect 34966 88102 35018 88154
rect 35030 88102 35082 88154
rect 35094 88102 35146 88154
rect 35158 88102 35210 88154
rect 65686 88102 65738 88154
rect 65750 88102 65802 88154
rect 65814 88102 65866 88154
rect 65878 88102 65930 88154
rect 96406 88102 96458 88154
rect 96470 88102 96522 88154
rect 96534 88102 96586 88154
rect 96598 88102 96650 88154
rect 127126 88102 127178 88154
rect 127190 88102 127242 88154
rect 127254 88102 127306 88154
rect 127318 88102 127370 88154
rect 157846 88102 157898 88154
rect 157910 88102 157962 88154
rect 157974 88102 158026 88154
rect 158038 88102 158090 88154
rect 19606 87558 19658 87610
rect 19670 87558 19722 87610
rect 19734 87558 19786 87610
rect 19798 87558 19850 87610
rect 50326 87558 50378 87610
rect 50390 87558 50442 87610
rect 50454 87558 50506 87610
rect 50518 87558 50570 87610
rect 81046 87558 81098 87610
rect 81110 87558 81162 87610
rect 81174 87558 81226 87610
rect 81238 87558 81290 87610
rect 111766 87558 111818 87610
rect 111830 87558 111882 87610
rect 111894 87558 111946 87610
rect 111958 87558 112010 87610
rect 142486 87558 142538 87610
rect 142550 87558 142602 87610
rect 142614 87558 142666 87610
rect 142678 87558 142730 87610
rect 173206 87558 173258 87610
rect 173270 87558 173322 87610
rect 173334 87558 173386 87610
rect 173398 87558 173450 87610
rect 4246 87014 4298 87066
rect 4310 87014 4362 87066
rect 4374 87014 4426 87066
rect 4438 87014 4490 87066
rect 34966 87014 35018 87066
rect 35030 87014 35082 87066
rect 35094 87014 35146 87066
rect 35158 87014 35210 87066
rect 65686 87014 65738 87066
rect 65750 87014 65802 87066
rect 65814 87014 65866 87066
rect 65878 87014 65930 87066
rect 96406 87014 96458 87066
rect 96470 87014 96522 87066
rect 96534 87014 96586 87066
rect 96598 87014 96650 87066
rect 127126 87014 127178 87066
rect 127190 87014 127242 87066
rect 127254 87014 127306 87066
rect 127318 87014 127370 87066
rect 157846 87014 157898 87066
rect 157910 87014 157962 87066
rect 157974 87014 158026 87066
rect 158038 87014 158090 87066
rect 19606 86470 19658 86522
rect 19670 86470 19722 86522
rect 19734 86470 19786 86522
rect 19798 86470 19850 86522
rect 50326 86470 50378 86522
rect 50390 86470 50442 86522
rect 50454 86470 50506 86522
rect 50518 86470 50570 86522
rect 81046 86470 81098 86522
rect 81110 86470 81162 86522
rect 81174 86470 81226 86522
rect 81238 86470 81290 86522
rect 111766 86470 111818 86522
rect 111830 86470 111882 86522
rect 111894 86470 111946 86522
rect 111958 86470 112010 86522
rect 142486 86470 142538 86522
rect 142550 86470 142602 86522
rect 142614 86470 142666 86522
rect 142678 86470 142730 86522
rect 173206 86470 173258 86522
rect 173270 86470 173322 86522
rect 173334 86470 173386 86522
rect 173398 86470 173450 86522
rect 4246 85926 4298 85978
rect 4310 85926 4362 85978
rect 4374 85926 4426 85978
rect 4438 85926 4490 85978
rect 34966 85926 35018 85978
rect 35030 85926 35082 85978
rect 35094 85926 35146 85978
rect 35158 85926 35210 85978
rect 65686 85926 65738 85978
rect 65750 85926 65802 85978
rect 65814 85926 65866 85978
rect 65878 85926 65930 85978
rect 96406 85926 96458 85978
rect 96470 85926 96522 85978
rect 96534 85926 96586 85978
rect 96598 85926 96650 85978
rect 127126 85926 127178 85978
rect 127190 85926 127242 85978
rect 127254 85926 127306 85978
rect 127318 85926 127370 85978
rect 157846 85926 157898 85978
rect 157910 85926 157962 85978
rect 157974 85926 158026 85978
rect 158038 85926 158090 85978
rect 19606 85382 19658 85434
rect 19670 85382 19722 85434
rect 19734 85382 19786 85434
rect 19798 85382 19850 85434
rect 50326 85382 50378 85434
rect 50390 85382 50442 85434
rect 50454 85382 50506 85434
rect 50518 85382 50570 85434
rect 81046 85382 81098 85434
rect 81110 85382 81162 85434
rect 81174 85382 81226 85434
rect 81238 85382 81290 85434
rect 111766 85382 111818 85434
rect 111830 85382 111882 85434
rect 111894 85382 111946 85434
rect 111958 85382 112010 85434
rect 142486 85382 142538 85434
rect 142550 85382 142602 85434
rect 142614 85382 142666 85434
rect 142678 85382 142730 85434
rect 173206 85382 173258 85434
rect 173270 85382 173322 85434
rect 173334 85382 173386 85434
rect 173398 85382 173450 85434
rect 4246 84838 4298 84890
rect 4310 84838 4362 84890
rect 4374 84838 4426 84890
rect 4438 84838 4490 84890
rect 34966 84838 35018 84890
rect 35030 84838 35082 84890
rect 35094 84838 35146 84890
rect 35158 84838 35210 84890
rect 65686 84838 65738 84890
rect 65750 84838 65802 84890
rect 65814 84838 65866 84890
rect 65878 84838 65930 84890
rect 96406 84838 96458 84890
rect 96470 84838 96522 84890
rect 96534 84838 96586 84890
rect 96598 84838 96650 84890
rect 127126 84838 127178 84890
rect 127190 84838 127242 84890
rect 127254 84838 127306 84890
rect 127318 84838 127370 84890
rect 157846 84838 157898 84890
rect 157910 84838 157962 84890
rect 157974 84838 158026 84890
rect 158038 84838 158090 84890
rect 19606 84294 19658 84346
rect 19670 84294 19722 84346
rect 19734 84294 19786 84346
rect 19798 84294 19850 84346
rect 50326 84294 50378 84346
rect 50390 84294 50442 84346
rect 50454 84294 50506 84346
rect 50518 84294 50570 84346
rect 81046 84294 81098 84346
rect 81110 84294 81162 84346
rect 81174 84294 81226 84346
rect 81238 84294 81290 84346
rect 111766 84294 111818 84346
rect 111830 84294 111882 84346
rect 111894 84294 111946 84346
rect 111958 84294 112010 84346
rect 142486 84294 142538 84346
rect 142550 84294 142602 84346
rect 142614 84294 142666 84346
rect 142678 84294 142730 84346
rect 173206 84294 173258 84346
rect 173270 84294 173322 84346
rect 173334 84294 173386 84346
rect 173398 84294 173450 84346
rect 4246 83750 4298 83802
rect 4310 83750 4362 83802
rect 4374 83750 4426 83802
rect 4438 83750 4490 83802
rect 34966 83750 35018 83802
rect 35030 83750 35082 83802
rect 35094 83750 35146 83802
rect 35158 83750 35210 83802
rect 65686 83750 65738 83802
rect 65750 83750 65802 83802
rect 65814 83750 65866 83802
rect 65878 83750 65930 83802
rect 96406 83750 96458 83802
rect 96470 83750 96522 83802
rect 96534 83750 96586 83802
rect 96598 83750 96650 83802
rect 127126 83750 127178 83802
rect 127190 83750 127242 83802
rect 127254 83750 127306 83802
rect 127318 83750 127370 83802
rect 157846 83750 157898 83802
rect 157910 83750 157962 83802
rect 157974 83750 158026 83802
rect 158038 83750 158090 83802
rect 19606 83206 19658 83258
rect 19670 83206 19722 83258
rect 19734 83206 19786 83258
rect 19798 83206 19850 83258
rect 50326 83206 50378 83258
rect 50390 83206 50442 83258
rect 50454 83206 50506 83258
rect 50518 83206 50570 83258
rect 81046 83206 81098 83258
rect 81110 83206 81162 83258
rect 81174 83206 81226 83258
rect 81238 83206 81290 83258
rect 111766 83206 111818 83258
rect 111830 83206 111882 83258
rect 111894 83206 111946 83258
rect 111958 83206 112010 83258
rect 142486 83206 142538 83258
rect 142550 83206 142602 83258
rect 142614 83206 142666 83258
rect 142678 83206 142730 83258
rect 173206 83206 173258 83258
rect 173270 83206 173322 83258
rect 173334 83206 173386 83258
rect 173398 83206 173450 83258
rect 4246 82662 4298 82714
rect 4310 82662 4362 82714
rect 4374 82662 4426 82714
rect 4438 82662 4490 82714
rect 34966 82662 35018 82714
rect 35030 82662 35082 82714
rect 35094 82662 35146 82714
rect 35158 82662 35210 82714
rect 65686 82662 65738 82714
rect 65750 82662 65802 82714
rect 65814 82662 65866 82714
rect 65878 82662 65930 82714
rect 96406 82662 96458 82714
rect 96470 82662 96522 82714
rect 96534 82662 96586 82714
rect 96598 82662 96650 82714
rect 127126 82662 127178 82714
rect 127190 82662 127242 82714
rect 127254 82662 127306 82714
rect 127318 82662 127370 82714
rect 157846 82662 157898 82714
rect 157910 82662 157962 82714
rect 157974 82662 158026 82714
rect 158038 82662 158090 82714
rect 19606 82118 19658 82170
rect 19670 82118 19722 82170
rect 19734 82118 19786 82170
rect 19798 82118 19850 82170
rect 50326 82118 50378 82170
rect 50390 82118 50442 82170
rect 50454 82118 50506 82170
rect 50518 82118 50570 82170
rect 81046 82118 81098 82170
rect 81110 82118 81162 82170
rect 81174 82118 81226 82170
rect 81238 82118 81290 82170
rect 111766 82118 111818 82170
rect 111830 82118 111882 82170
rect 111894 82118 111946 82170
rect 111958 82118 112010 82170
rect 142486 82118 142538 82170
rect 142550 82118 142602 82170
rect 142614 82118 142666 82170
rect 142678 82118 142730 82170
rect 173206 82118 173258 82170
rect 173270 82118 173322 82170
rect 173334 82118 173386 82170
rect 173398 82118 173450 82170
rect 4246 81574 4298 81626
rect 4310 81574 4362 81626
rect 4374 81574 4426 81626
rect 4438 81574 4490 81626
rect 34966 81574 35018 81626
rect 35030 81574 35082 81626
rect 35094 81574 35146 81626
rect 35158 81574 35210 81626
rect 65686 81574 65738 81626
rect 65750 81574 65802 81626
rect 65814 81574 65866 81626
rect 65878 81574 65930 81626
rect 96406 81574 96458 81626
rect 96470 81574 96522 81626
rect 96534 81574 96586 81626
rect 96598 81574 96650 81626
rect 127126 81574 127178 81626
rect 127190 81574 127242 81626
rect 127254 81574 127306 81626
rect 127318 81574 127370 81626
rect 157846 81574 157898 81626
rect 157910 81574 157962 81626
rect 157974 81574 158026 81626
rect 158038 81574 158090 81626
rect 19606 81030 19658 81082
rect 19670 81030 19722 81082
rect 19734 81030 19786 81082
rect 19798 81030 19850 81082
rect 50326 81030 50378 81082
rect 50390 81030 50442 81082
rect 50454 81030 50506 81082
rect 50518 81030 50570 81082
rect 81046 81030 81098 81082
rect 81110 81030 81162 81082
rect 81174 81030 81226 81082
rect 81238 81030 81290 81082
rect 111766 81030 111818 81082
rect 111830 81030 111882 81082
rect 111894 81030 111946 81082
rect 111958 81030 112010 81082
rect 142486 81030 142538 81082
rect 142550 81030 142602 81082
rect 142614 81030 142666 81082
rect 142678 81030 142730 81082
rect 173206 81030 173258 81082
rect 173270 81030 173322 81082
rect 173334 81030 173386 81082
rect 173398 81030 173450 81082
rect 4246 80486 4298 80538
rect 4310 80486 4362 80538
rect 4374 80486 4426 80538
rect 4438 80486 4490 80538
rect 34966 80486 35018 80538
rect 35030 80486 35082 80538
rect 35094 80486 35146 80538
rect 35158 80486 35210 80538
rect 65686 80486 65738 80538
rect 65750 80486 65802 80538
rect 65814 80486 65866 80538
rect 65878 80486 65930 80538
rect 96406 80486 96458 80538
rect 96470 80486 96522 80538
rect 96534 80486 96586 80538
rect 96598 80486 96650 80538
rect 127126 80486 127178 80538
rect 127190 80486 127242 80538
rect 127254 80486 127306 80538
rect 127318 80486 127370 80538
rect 157846 80486 157898 80538
rect 157910 80486 157962 80538
rect 157974 80486 158026 80538
rect 158038 80486 158090 80538
rect 19606 79942 19658 79994
rect 19670 79942 19722 79994
rect 19734 79942 19786 79994
rect 19798 79942 19850 79994
rect 50326 79942 50378 79994
rect 50390 79942 50442 79994
rect 50454 79942 50506 79994
rect 50518 79942 50570 79994
rect 81046 79942 81098 79994
rect 81110 79942 81162 79994
rect 81174 79942 81226 79994
rect 81238 79942 81290 79994
rect 111766 79942 111818 79994
rect 111830 79942 111882 79994
rect 111894 79942 111946 79994
rect 111958 79942 112010 79994
rect 142486 79942 142538 79994
rect 142550 79942 142602 79994
rect 142614 79942 142666 79994
rect 142678 79942 142730 79994
rect 173206 79942 173258 79994
rect 173270 79942 173322 79994
rect 173334 79942 173386 79994
rect 173398 79942 173450 79994
rect 4246 79398 4298 79450
rect 4310 79398 4362 79450
rect 4374 79398 4426 79450
rect 4438 79398 4490 79450
rect 34966 79398 35018 79450
rect 35030 79398 35082 79450
rect 35094 79398 35146 79450
rect 35158 79398 35210 79450
rect 65686 79398 65738 79450
rect 65750 79398 65802 79450
rect 65814 79398 65866 79450
rect 65878 79398 65930 79450
rect 96406 79398 96458 79450
rect 96470 79398 96522 79450
rect 96534 79398 96586 79450
rect 96598 79398 96650 79450
rect 127126 79398 127178 79450
rect 127190 79398 127242 79450
rect 127254 79398 127306 79450
rect 127318 79398 127370 79450
rect 157846 79398 157898 79450
rect 157910 79398 157962 79450
rect 157974 79398 158026 79450
rect 158038 79398 158090 79450
rect 19606 78854 19658 78906
rect 19670 78854 19722 78906
rect 19734 78854 19786 78906
rect 19798 78854 19850 78906
rect 50326 78854 50378 78906
rect 50390 78854 50442 78906
rect 50454 78854 50506 78906
rect 50518 78854 50570 78906
rect 81046 78854 81098 78906
rect 81110 78854 81162 78906
rect 81174 78854 81226 78906
rect 81238 78854 81290 78906
rect 111766 78854 111818 78906
rect 111830 78854 111882 78906
rect 111894 78854 111946 78906
rect 111958 78854 112010 78906
rect 142486 78854 142538 78906
rect 142550 78854 142602 78906
rect 142614 78854 142666 78906
rect 142678 78854 142730 78906
rect 173206 78854 173258 78906
rect 173270 78854 173322 78906
rect 173334 78854 173386 78906
rect 173398 78854 173450 78906
rect 4246 78310 4298 78362
rect 4310 78310 4362 78362
rect 4374 78310 4426 78362
rect 4438 78310 4490 78362
rect 34966 78310 35018 78362
rect 35030 78310 35082 78362
rect 35094 78310 35146 78362
rect 35158 78310 35210 78362
rect 65686 78310 65738 78362
rect 65750 78310 65802 78362
rect 65814 78310 65866 78362
rect 65878 78310 65930 78362
rect 96406 78310 96458 78362
rect 96470 78310 96522 78362
rect 96534 78310 96586 78362
rect 96598 78310 96650 78362
rect 127126 78310 127178 78362
rect 127190 78310 127242 78362
rect 127254 78310 127306 78362
rect 127318 78310 127370 78362
rect 157846 78310 157898 78362
rect 157910 78310 157962 78362
rect 157974 78310 158026 78362
rect 158038 78310 158090 78362
rect 19606 77766 19658 77818
rect 19670 77766 19722 77818
rect 19734 77766 19786 77818
rect 19798 77766 19850 77818
rect 50326 77766 50378 77818
rect 50390 77766 50442 77818
rect 50454 77766 50506 77818
rect 50518 77766 50570 77818
rect 81046 77766 81098 77818
rect 81110 77766 81162 77818
rect 81174 77766 81226 77818
rect 81238 77766 81290 77818
rect 111766 77766 111818 77818
rect 111830 77766 111882 77818
rect 111894 77766 111946 77818
rect 111958 77766 112010 77818
rect 142486 77766 142538 77818
rect 142550 77766 142602 77818
rect 142614 77766 142666 77818
rect 142678 77766 142730 77818
rect 173206 77766 173258 77818
rect 173270 77766 173322 77818
rect 173334 77766 173386 77818
rect 173398 77766 173450 77818
rect 4246 77222 4298 77274
rect 4310 77222 4362 77274
rect 4374 77222 4426 77274
rect 4438 77222 4490 77274
rect 34966 77222 35018 77274
rect 35030 77222 35082 77274
rect 35094 77222 35146 77274
rect 35158 77222 35210 77274
rect 65686 77222 65738 77274
rect 65750 77222 65802 77274
rect 65814 77222 65866 77274
rect 65878 77222 65930 77274
rect 96406 77222 96458 77274
rect 96470 77222 96522 77274
rect 96534 77222 96586 77274
rect 96598 77222 96650 77274
rect 127126 77222 127178 77274
rect 127190 77222 127242 77274
rect 127254 77222 127306 77274
rect 127318 77222 127370 77274
rect 157846 77222 157898 77274
rect 157910 77222 157962 77274
rect 157974 77222 158026 77274
rect 158038 77222 158090 77274
rect 19606 76678 19658 76730
rect 19670 76678 19722 76730
rect 19734 76678 19786 76730
rect 19798 76678 19850 76730
rect 50326 76678 50378 76730
rect 50390 76678 50442 76730
rect 50454 76678 50506 76730
rect 50518 76678 50570 76730
rect 81046 76678 81098 76730
rect 81110 76678 81162 76730
rect 81174 76678 81226 76730
rect 81238 76678 81290 76730
rect 111766 76678 111818 76730
rect 111830 76678 111882 76730
rect 111894 76678 111946 76730
rect 111958 76678 112010 76730
rect 142486 76678 142538 76730
rect 142550 76678 142602 76730
rect 142614 76678 142666 76730
rect 142678 76678 142730 76730
rect 173206 76678 173258 76730
rect 173270 76678 173322 76730
rect 173334 76678 173386 76730
rect 173398 76678 173450 76730
rect 4246 76134 4298 76186
rect 4310 76134 4362 76186
rect 4374 76134 4426 76186
rect 4438 76134 4490 76186
rect 34966 76134 35018 76186
rect 35030 76134 35082 76186
rect 35094 76134 35146 76186
rect 35158 76134 35210 76186
rect 65686 76134 65738 76186
rect 65750 76134 65802 76186
rect 65814 76134 65866 76186
rect 65878 76134 65930 76186
rect 96406 76134 96458 76186
rect 96470 76134 96522 76186
rect 96534 76134 96586 76186
rect 96598 76134 96650 76186
rect 127126 76134 127178 76186
rect 127190 76134 127242 76186
rect 127254 76134 127306 76186
rect 127318 76134 127370 76186
rect 157846 76134 157898 76186
rect 157910 76134 157962 76186
rect 157974 76134 158026 76186
rect 158038 76134 158090 76186
rect 19606 75590 19658 75642
rect 19670 75590 19722 75642
rect 19734 75590 19786 75642
rect 19798 75590 19850 75642
rect 50326 75590 50378 75642
rect 50390 75590 50442 75642
rect 50454 75590 50506 75642
rect 50518 75590 50570 75642
rect 81046 75590 81098 75642
rect 81110 75590 81162 75642
rect 81174 75590 81226 75642
rect 81238 75590 81290 75642
rect 111766 75590 111818 75642
rect 111830 75590 111882 75642
rect 111894 75590 111946 75642
rect 111958 75590 112010 75642
rect 142486 75590 142538 75642
rect 142550 75590 142602 75642
rect 142614 75590 142666 75642
rect 142678 75590 142730 75642
rect 173206 75590 173258 75642
rect 173270 75590 173322 75642
rect 173334 75590 173386 75642
rect 173398 75590 173450 75642
rect 4246 75046 4298 75098
rect 4310 75046 4362 75098
rect 4374 75046 4426 75098
rect 4438 75046 4490 75098
rect 34966 75046 35018 75098
rect 35030 75046 35082 75098
rect 35094 75046 35146 75098
rect 35158 75046 35210 75098
rect 65686 75046 65738 75098
rect 65750 75046 65802 75098
rect 65814 75046 65866 75098
rect 65878 75046 65930 75098
rect 96406 75046 96458 75098
rect 96470 75046 96522 75098
rect 96534 75046 96586 75098
rect 96598 75046 96650 75098
rect 127126 75046 127178 75098
rect 127190 75046 127242 75098
rect 127254 75046 127306 75098
rect 127318 75046 127370 75098
rect 157846 75046 157898 75098
rect 157910 75046 157962 75098
rect 157974 75046 158026 75098
rect 158038 75046 158090 75098
rect 19606 74502 19658 74554
rect 19670 74502 19722 74554
rect 19734 74502 19786 74554
rect 19798 74502 19850 74554
rect 50326 74502 50378 74554
rect 50390 74502 50442 74554
rect 50454 74502 50506 74554
rect 50518 74502 50570 74554
rect 81046 74502 81098 74554
rect 81110 74502 81162 74554
rect 81174 74502 81226 74554
rect 81238 74502 81290 74554
rect 111766 74502 111818 74554
rect 111830 74502 111882 74554
rect 111894 74502 111946 74554
rect 111958 74502 112010 74554
rect 142486 74502 142538 74554
rect 142550 74502 142602 74554
rect 142614 74502 142666 74554
rect 142678 74502 142730 74554
rect 173206 74502 173258 74554
rect 173270 74502 173322 74554
rect 173334 74502 173386 74554
rect 173398 74502 173450 74554
rect 4246 73958 4298 74010
rect 4310 73958 4362 74010
rect 4374 73958 4426 74010
rect 4438 73958 4490 74010
rect 34966 73958 35018 74010
rect 35030 73958 35082 74010
rect 35094 73958 35146 74010
rect 35158 73958 35210 74010
rect 65686 73958 65738 74010
rect 65750 73958 65802 74010
rect 65814 73958 65866 74010
rect 65878 73958 65930 74010
rect 96406 73958 96458 74010
rect 96470 73958 96522 74010
rect 96534 73958 96586 74010
rect 96598 73958 96650 74010
rect 127126 73958 127178 74010
rect 127190 73958 127242 74010
rect 127254 73958 127306 74010
rect 127318 73958 127370 74010
rect 157846 73958 157898 74010
rect 157910 73958 157962 74010
rect 157974 73958 158026 74010
rect 158038 73958 158090 74010
rect 19606 73414 19658 73466
rect 19670 73414 19722 73466
rect 19734 73414 19786 73466
rect 19798 73414 19850 73466
rect 50326 73414 50378 73466
rect 50390 73414 50442 73466
rect 50454 73414 50506 73466
rect 50518 73414 50570 73466
rect 81046 73414 81098 73466
rect 81110 73414 81162 73466
rect 81174 73414 81226 73466
rect 81238 73414 81290 73466
rect 111766 73414 111818 73466
rect 111830 73414 111882 73466
rect 111894 73414 111946 73466
rect 111958 73414 112010 73466
rect 142486 73414 142538 73466
rect 142550 73414 142602 73466
rect 142614 73414 142666 73466
rect 142678 73414 142730 73466
rect 173206 73414 173258 73466
rect 173270 73414 173322 73466
rect 173334 73414 173386 73466
rect 173398 73414 173450 73466
rect 4246 72870 4298 72922
rect 4310 72870 4362 72922
rect 4374 72870 4426 72922
rect 4438 72870 4490 72922
rect 34966 72870 35018 72922
rect 35030 72870 35082 72922
rect 35094 72870 35146 72922
rect 35158 72870 35210 72922
rect 65686 72870 65738 72922
rect 65750 72870 65802 72922
rect 65814 72870 65866 72922
rect 65878 72870 65930 72922
rect 96406 72870 96458 72922
rect 96470 72870 96522 72922
rect 96534 72870 96586 72922
rect 96598 72870 96650 72922
rect 127126 72870 127178 72922
rect 127190 72870 127242 72922
rect 127254 72870 127306 72922
rect 127318 72870 127370 72922
rect 157846 72870 157898 72922
rect 157910 72870 157962 72922
rect 157974 72870 158026 72922
rect 158038 72870 158090 72922
rect 19606 72326 19658 72378
rect 19670 72326 19722 72378
rect 19734 72326 19786 72378
rect 19798 72326 19850 72378
rect 50326 72326 50378 72378
rect 50390 72326 50442 72378
rect 50454 72326 50506 72378
rect 50518 72326 50570 72378
rect 81046 72326 81098 72378
rect 81110 72326 81162 72378
rect 81174 72326 81226 72378
rect 81238 72326 81290 72378
rect 111766 72326 111818 72378
rect 111830 72326 111882 72378
rect 111894 72326 111946 72378
rect 111958 72326 112010 72378
rect 142486 72326 142538 72378
rect 142550 72326 142602 72378
rect 142614 72326 142666 72378
rect 142678 72326 142730 72378
rect 173206 72326 173258 72378
rect 173270 72326 173322 72378
rect 173334 72326 173386 72378
rect 173398 72326 173450 72378
rect 4246 71782 4298 71834
rect 4310 71782 4362 71834
rect 4374 71782 4426 71834
rect 4438 71782 4490 71834
rect 34966 71782 35018 71834
rect 35030 71782 35082 71834
rect 35094 71782 35146 71834
rect 35158 71782 35210 71834
rect 65686 71782 65738 71834
rect 65750 71782 65802 71834
rect 65814 71782 65866 71834
rect 65878 71782 65930 71834
rect 96406 71782 96458 71834
rect 96470 71782 96522 71834
rect 96534 71782 96586 71834
rect 96598 71782 96650 71834
rect 127126 71782 127178 71834
rect 127190 71782 127242 71834
rect 127254 71782 127306 71834
rect 127318 71782 127370 71834
rect 157846 71782 157898 71834
rect 157910 71782 157962 71834
rect 157974 71782 158026 71834
rect 158038 71782 158090 71834
rect 19606 71238 19658 71290
rect 19670 71238 19722 71290
rect 19734 71238 19786 71290
rect 19798 71238 19850 71290
rect 50326 71238 50378 71290
rect 50390 71238 50442 71290
rect 50454 71238 50506 71290
rect 50518 71238 50570 71290
rect 81046 71238 81098 71290
rect 81110 71238 81162 71290
rect 81174 71238 81226 71290
rect 81238 71238 81290 71290
rect 111766 71238 111818 71290
rect 111830 71238 111882 71290
rect 111894 71238 111946 71290
rect 111958 71238 112010 71290
rect 142486 71238 142538 71290
rect 142550 71238 142602 71290
rect 142614 71238 142666 71290
rect 142678 71238 142730 71290
rect 173206 71238 173258 71290
rect 173270 71238 173322 71290
rect 173334 71238 173386 71290
rect 173398 71238 173450 71290
rect 4246 70694 4298 70746
rect 4310 70694 4362 70746
rect 4374 70694 4426 70746
rect 4438 70694 4490 70746
rect 34966 70694 35018 70746
rect 35030 70694 35082 70746
rect 35094 70694 35146 70746
rect 35158 70694 35210 70746
rect 65686 70694 65738 70746
rect 65750 70694 65802 70746
rect 65814 70694 65866 70746
rect 65878 70694 65930 70746
rect 96406 70694 96458 70746
rect 96470 70694 96522 70746
rect 96534 70694 96586 70746
rect 96598 70694 96650 70746
rect 127126 70694 127178 70746
rect 127190 70694 127242 70746
rect 127254 70694 127306 70746
rect 127318 70694 127370 70746
rect 157846 70694 157898 70746
rect 157910 70694 157962 70746
rect 157974 70694 158026 70746
rect 158038 70694 158090 70746
rect 19606 70150 19658 70202
rect 19670 70150 19722 70202
rect 19734 70150 19786 70202
rect 19798 70150 19850 70202
rect 50326 70150 50378 70202
rect 50390 70150 50442 70202
rect 50454 70150 50506 70202
rect 50518 70150 50570 70202
rect 81046 70150 81098 70202
rect 81110 70150 81162 70202
rect 81174 70150 81226 70202
rect 81238 70150 81290 70202
rect 111766 70150 111818 70202
rect 111830 70150 111882 70202
rect 111894 70150 111946 70202
rect 111958 70150 112010 70202
rect 142486 70150 142538 70202
rect 142550 70150 142602 70202
rect 142614 70150 142666 70202
rect 142678 70150 142730 70202
rect 173206 70150 173258 70202
rect 173270 70150 173322 70202
rect 173334 70150 173386 70202
rect 173398 70150 173450 70202
rect 4246 69606 4298 69658
rect 4310 69606 4362 69658
rect 4374 69606 4426 69658
rect 4438 69606 4490 69658
rect 34966 69606 35018 69658
rect 35030 69606 35082 69658
rect 35094 69606 35146 69658
rect 35158 69606 35210 69658
rect 65686 69606 65738 69658
rect 65750 69606 65802 69658
rect 65814 69606 65866 69658
rect 65878 69606 65930 69658
rect 96406 69606 96458 69658
rect 96470 69606 96522 69658
rect 96534 69606 96586 69658
rect 96598 69606 96650 69658
rect 127126 69606 127178 69658
rect 127190 69606 127242 69658
rect 127254 69606 127306 69658
rect 127318 69606 127370 69658
rect 157846 69606 157898 69658
rect 157910 69606 157962 69658
rect 157974 69606 158026 69658
rect 158038 69606 158090 69658
rect 19606 69062 19658 69114
rect 19670 69062 19722 69114
rect 19734 69062 19786 69114
rect 19798 69062 19850 69114
rect 50326 69062 50378 69114
rect 50390 69062 50442 69114
rect 50454 69062 50506 69114
rect 50518 69062 50570 69114
rect 81046 69062 81098 69114
rect 81110 69062 81162 69114
rect 81174 69062 81226 69114
rect 81238 69062 81290 69114
rect 111766 69062 111818 69114
rect 111830 69062 111882 69114
rect 111894 69062 111946 69114
rect 111958 69062 112010 69114
rect 142486 69062 142538 69114
rect 142550 69062 142602 69114
rect 142614 69062 142666 69114
rect 142678 69062 142730 69114
rect 173206 69062 173258 69114
rect 173270 69062 173322 69114
rect 173334 69062 173386 69114
rect 173398 69062 173450 69114
rect 4246 68518 4298 68570
rect 4310 68518 4362 68570
rect 4374 68518 4426 68570
rect 4438 68518 4490 68570
rect 34966 68518 35018 68570
rect 35030 68518 35082 68570
rect 35094 68518 35146 68570
rect 35158 68518 35210 68570
rect 65686 68518 65738 68570
rect 65750 68518 65802 68570
rect 65814 68518 65866 68570
rect 65878 68518 65930 68570
rect 96406 68518 96458 68570
rect 96470 68518 96522 68570
rect 96534 68518 96586 68570
rect 96598 68518 96650 68570
rect 127126 68518 127178 68570
rect 127190 68518 127242 68570
rect 127254 68518 127306 68570
rect 127318 68518 127370 68570
rect 157846 68518 157898 68570
rect 157910 68518 157962 68570
rect 157974 68518 158026 68570
rect 158038 68518 158090 68570
rect 19606 67974 19658 68026
rect 19670 67974 19722 68026
rect 19734 67974 19786 68026
rect 19798 67974 19850 68026
rect 50326 67974 50378 68026
rect 50390 67974 50442 68026
rect 50454 67974 50506 68026
rect 50518 67974 50570 68026
rect 81046 67974 81098 68026
rect 81110 67974 81162 68026
rect 81174 67974 81226 68026
rect 81238 67974 81290 68026
rect 111766 67974 111818 68026
rect 111830 67974 111882 68026
rect 111894 67974 111946 68026
rect 111958 67974 112010 68026
rect 142486 67974 142538 68026
rect 142550 67974 142602 68026
rect 142614 67974 142666 68026
rect 142678 67974 142730 68026
rect 173206 67974 173258 68026
rect 173270 67974 173322 68026
rect 173334 67974 173386 68026
rect 173398 67974 173450 68026
rect 4246 67430 4298 67482
rect 4310 67430 4362 67482
rect 4374 67430 4426 67482
rect 4438 67430 4490 67482
rect 34966 67430 35018 67482
rect 35030 67430 35082 67482
rect 35094 67430 35146 67482
rect 35158 67430 35210 67482
rect 65686 67430 65738 67482
rect 65750 67430 65802 67482
rect 65814 67430 65866 67482
rect 65878 67430 65930 67482
rect 96406 67430 96458 67482
rect 96470 67430 96522 67482
rect 96534 67430 96586 67482
rect 96598 67430 96650 67482
rect 127126 67430 127178 67482
rect 127190 67430 127242 67482
rect 127254 67430 127306 67482
rect 127318 67430 127370 67482
rect 157846 67430 157898 67482
rect 157910 67430 157962 67482
rect 157974 67430 158026 67482
rect 158038 67430 158090 67482
rect 19606 66886 19658 66938
rect 19670 66886 19722 66938
rect 19734 66886 19786 66938
rect 19798 66886 19850 66938
rect 50326 66886 50378 66938
rect 50390 66886 50442 66938
rect 50454 66886 50506 66938
rect 50518 66886 50570 66938
rect 81046 66886 81098 66938
rect 81110 66886 81162 66938
rect 81174 66886 81226 66938
rect 81238 66886 81290 66938
rect 111766 66886 111818 66938
rect 111830 66886 111882 66938
rect 111894 66886 111946 66938
rect 111958 66886 112010 66938
rect 142486 66886 142538 66938
rect 142550 66886 142602 66938
rect 142614 66886 142666 66938
rect 142678 66886 142730 66938
rect 173206 66886 173258 66938
rect 173270 66886 173322 66938
rect 173334 66886 173386 66938
rect 173398 66886 173450 66938
rect 4246 66342 4298 66394
rect 4310 66342 4362 66394
rect 4374 66342 4426 66394
rect 4438 66342 4490 66394
rect 34966 66342 35018 66394
rect 35030 66342 35082 66394
rect 35094 66342 35146 66394
rect 35158 66342 35210 66394
rect 65686 66342 65738 66394
rect 65750 66342 65802 66394
rect 65814 66342 65866 66394
rect 65878 66342 65930 66394
rect 96406 66342 96458 66394
rect 96470 66342 96522 66394
rect 96534 66342 96586 66394
rect 96598 66342 96650 66394
rect 127126 66342 127178 66394
rect 127190 66342 127242 66394
rect 127254 66342 127306 66394
rect 127318 66342 127370 66394
rect 157846 66342 157898 66394
rect 157910 66342 157962 66394
rect 157974 66342 158026 66394
rect 158038 66342 158090 66394
rect 19606 65798 19658 65850
rect 19670 65798 19722 65850
rect 19734 65798 19786 65850
rect 19798 65798 19850 65850
rect 50326 65798 50378 65850
rect 50390 65798 50442 65850
rect 50454 65798 50506 65850
rect 50518 65798 50570 65850
rect 81046 65798 81098 65850
rect 81110 65798 81162 65850
rect 81174 65798 81226 65850
rect 81238 65798 81290 65850
rect 111766 65798 111818 65850
rect 111830 65798 111882 65850
rect 111894 65798 111946 65850
rect 111958 65798 112010 65850
rect 142486 65798 142538 65850
rect 142550 65798 142602 65850
rect 142614 65798 142666 65850
rect 142678 65798 142730 65850
rect 173206 65798 173258 65850
rect 173270 65798 173322 65850
rect 173334 65798 173386 65850
rect 173398 65798 173450 65850
rect 4246 65254 4298 65306
rect 4310 65254 4362 65306
rect 4374 65254 4426 65306
rect 4438 65254 4490 65306
rect 34966 65254 35018 65306
rect 35030 65254 35082 65306
rect 35094 65254 35146 65306
rect 35158 65254 35210 65306
rect 65686 65254 65738 65306
rect 65750 65254 65802 65306
rect 65814 65254 65866 65306
rect 65878 65254 65930 65306
rect 96406 65254 96458 65306
rect 96470 65254 96522 65306
rect 96534 65254 96586 65306
rect 96598 65254 96650 65306
rect 127126 65254 127178 65306
rect 127190 65254 127242 65306
rect 127254 65254 127306 65306
rect 127318 65254 127370 65306
rect 157846 65254 157898 65306
rect 157910 65254 157962 65306
rect 157974 65254 158026 65306
rect 158038 65254 158090 65306
rect 19606 64710 19658 64762
rect 19670 64710 19722 64762
rect 19734 64710 19786 64762
rect 19798 64710 19850 64762
rect 50326 64710 50378 64762
rect 50390 64710 50442 64762
rect 50454 64710 50506 64762
rect 50518 64710 50570 64762
rect 81046 64710 81098 64762
rect 81110 64710 81162 64762
rect 81174 64710 81226 64762
rect 81238 64710 81290 64762
rect 111766 64710 111818 64762
rect 111830 64710 111882 64762
rect 111894 64710 111946 64762
rect 111958 64710 112010 64762
rect 142486 64710 142538 64762
rect 142550 64710 142602 64762
rect 142614 64710 142666 64762
rect 142678 64710 142730 64762
rect 173206 64710 173258 64762
rect 173270 64710 173322 64762
rect 173334 64710 173386 64762
rect 173398 64710 173450 64762
rect 4246 64166 4298 64218
rect 4310 64166 4362 64218
rect 4374 64166 4426 64218
rect 4438 64166 4490 64218
rect 34966 64166 35018 64218
rect 35030 64166 35082 64218
rect 35094 64166 35146 64218
rect 35158 64166 35210 64218
rect 65686 64166 65738 64218
rect 65750 64166 65802 64218
rect 65814 64166 65866 64218
rect 65878 64166 65930 64218
rect 96406 64166 96458 64218
rect 96470 64166 96522 64218
rect 96534 64166 96586 64218
rect 96598 64166 96650 64218
rect 127126 64166 127178 64218
rect 127190 64166 127242 64218
rect 127254 64166 127306 64218
rect 127318 64166 127370 64218
rect 157846 64166 157898 64218
rect 157910 64166 157962 64218
rect 157974 64166 158026 64218
rect 158038 64166 158090 64218
rect 19606 63622 19658 63674
rect 19670 63622 19722 63674
rect 19734 63622 19786 63674
rect 19798 63622 19850 63674
rect 50326 63622 50378 63674
rect 50390 63622 50442 63674
rect 50454 63622 50506 63674
rect 50518 63622 50570 63674
rect 81046 63622 81098 63674
rect 81110 63622 81162 63674
rect 81174 63622 81226 63674
rect 81238 63622 81290 63674
rect 111766 63622 111818 63674
rect 111830 63622 111882 63674
rect 111894 63622 111946 63674
rect 111958 63622 112010 63674
rect 142486 63622 142538 63674
rect 142550 63622 142602 63674
rect 142614 63622 142666 63674
rect 142678 63622 142730 63674
rect 173206 63622 173258 63674
rect 173270 63622 173322 63674
rect 173334 63622 173386 63674
rect 173398 63622 173450 63674
rect 4246 63078 4298 63130
rect 4310 63078 4362 63130
rect 4374 63078 4426 63130
rect 4438 63078 4490 63130
rect 34966 63078 35018 63130
rect 35030 63078 35082 63130
rect 35094 63078 35146 63130
rect 35158 63078 35210 63130
rect 65686 63078 65738 63130
rect 65750 63078 65802 63130
rect 65814 63078 65866 63130
rect 65878 63078 65930 63130
rect 96406 63078 96458 63130
rect 96470 63078 96522 63130
rect 96534 63078 96586 63130
rect 96598 63078 96650 63130
rect 127126 63078 127178 63130
rect 127190 63078 127242 63130
rect 127254 63078 127306 63130
rect 127318 63078 127370 63130
rect 157846 63078 157898 63130
rect 157910 63078 157962 63130
rect 157974 63078 158026 63130
rect 158038 63078 158090 63130
rect 19606 62534 19658 62586
rect 19670 62534 19722 62586
rect 19734 62534 19786 62586
rect 19798 62534 19850 62586
rect 50326 62534 50378 62586
rect 50390 62534 50442 62586
rect 50454 62534 50506 62586
rect 50518 62534 50570 62586
rect 81046 62534 81098 62586
rect 81110 62534 81162 62586
rect 81174 62534 81226 62586
rect 81238 62534 81290 62586
rect 111766 62534 111818 62586
rect 111830 62534 111882 62586
rect 111894 62534 111946 62586
rect 111958 62534 112010 62586
rect 142486 62534 142538 62586
rect 142550 62534 142602 62586
rect 142614 62534 142666 62586
rect 142678 62534 142730 62586
rect 173206 62534 173258 62586
rect 173270 62534 173322 62586
rect 173334 62534 173386 62586
rect 173398 62534 173450 62586
rect 4246 61990 4298 62042
rect 4310 61990 4362 62042
rect 4374 61990 4426 62042
rect 4438 61990 4490 62042
rect 34966 61990 35018 62042
rect 35030 61990 35082 62042
rect 35094 61990 35146 62042
rect 35158 61990 35210 62042
rect 65686 61990 65738 62042
rect 65750 61990 65802 62042
rect 65814 61990 65866 62042
rect 65878 61990 65930 62042
rect 96406 61990 96458 62042
rect 96470 61990 96522 62042
rect 96534 61990 96586 62042
rect 96598 61990 96650 62042
rect 127126 61990 127178 62042
rect 127190 61990 127242 62042
rect 127254 61990 127306 62042
rect 127318 61990 127370 62042
rect 157846 61990 157898 62042
rect 157910 61990 157962 62042
rect 157974 61990 158026 62042
rect 158038 61990 158090 62042
rect 19606 61446 19658 61498
rect 19670 61446 19722 61498
rect 19734 61446 19786 61498
rect 19798 61446 19850 61498
rect 50326 61446 50378 61498
rect 50390 61446 50442 61498
rect 50454 61446 50506 61498
rect 50518 61446 50570 61498
rect 81046 61446 81098 61498
rect 81110 61446 81162 61498
rect 81174 61446 81226 61498
rect 81238 61446 81290 61498
rect 111766 61446 111818 61498
rect 111830 61446 111882 61498
rect 111894 61446 111946 61498
rect 111958 61446 112010 61498
rect 142486 61446 142538 61498
rect 142550 61446 142602 61498
rect 142614 61446 142666 61498
rect 142678 61446 142730 61498
rect 173206 61446 173258 61498
rect 173270 61446 173322 61498
rect 173334 61446 173386 61498
rect 173398 61446 173450 61498
rect 4246 60902 4298 60954
rect 4310 60902 4362 60954
rect 4374 60902 4426 60954
rect 4438 60902 4490 60954
rect 34966 60902 35018 60954
rect 35030 60902 35082 60954
rect 35094 60902 35146 60954
rect 35158 60902 35210 60954
rect 65686 60902 65738 60954
rect 65750 60902 65802 60954
rect 65814 60902 65866 60954
rect 65878 60902 65930 60954
rect 96406 60902 96458 60954
rect 96470 60902 96522 60954
rect 96534 60902 96586 60954
rect 96598 60902 96650 60954
rect 127126 60902 127178 60954
rect 127190 60902 127242 60954
rect 127254 60902 127306 60954
rect 127318 60902 127370 60954
rect 157846 60902 157898 60954
rect 157910 60902 157962 60954
rect 157974 60902 158026 60954
rect 158038 60902 158090 60954
rect 19606 60358 19658 60410
rect 19670 60358 19722 60410
rect 19734 60358 19786 60410
rect 19798 60358 19850 60410
rect 50326 60358 50378 60410
rect 50390 60358 50442 60410
rect 50454 60358 50506 60410
rect 50518 60358 50570 60410
rect 81046 60358 81098 60410
rect 81110 60358 81162 60410
rect 81174 60358 81226 60410
rect 81238 60358 81290 60410
rect 111766 60358 111818 60410
rect 111830 60358 111882 60410
rect 111894 60358 111946 60410
rect 111958 60358 112010 60410
rect 142486 60358 142538 60410
rect 142550 60358 142602 60410
rect 142614 60358 142666 60410
rect 142678 60358 142730 60410
rect 173206 60358 173258 60410
rect 173270 60358 173322 60410
rect 173334 60358 173386 60410
rect 173398 60358 173450 60410
rect 3056 60120 3108 60172
rect 176936 60120 176988 60172
rect 2044 60027 2096 60036
rect 2044 59993 2053 60027
rect 2053 59993 2087 60027
rect 2087 59993 2096 60027
rect 2044 59984 2096 59993
rect 178132 60027 178184 60036
rect 178132 59993 178141 60027
rect 178141 59993 178175 60027
rect 178175 59993 178184 60027
rect 178132 59984 178184 59993
rect 4246 59814 4298 59866
rect 4310 59814 4362 59866
rect 4374 59814 4426 59866
rect 4438 59814 4490 59866
rect 34966 59814 35018 59866
rect 35030 59814 35082 59866
rect 35094 59814 35146 59866
rect 35158 59814 35210 59866
rect 65686 59814 65738 59866
rect 65750 59814 65802 59866
rect 65814 59814 65866 59866
rect 65878 59814 65930 59866
rect 96406 59814 96458 59866
rect 96470 59814 96522 59866
rect 96534 59814 96586 59866
rect 96598 59814 96650 59866
rect 127126 59814 127178 59866
rect 127190 59814 127242 59866
rect 127254 59814 127306 59866
rect 127318 59814 127370 59866
rect 157846 59814 157898 59866
rect 157910 59814 157962 59866
rect 157974 59814 158026 59866
rect 158038 59814 158090 59866
rect 3056 59755 3108 59764
rect 3056 59721 3065 59755
rect 3065 59721 3099 59755
rect 3099 59721 3108 59755
rect 3056 59712 3108 59721
rect 176936 59755 176988 59764
rect 176936 59721 176945 59755
rect 176945 59721 176979 59755
rect 176979 59721 176988 59755
rect 176936 59712 176988 59721
rect 19606 59270 19658 59322
rect 19670 59270 19722 59322
rect 19734 59270 19786 59322
rect 19798 59270 19850 59322
rect 50326 59270 50378 59322
rect 50390 59270 50442 59322
rect 50454 59270 50506 59322
rect 50518 59270 50570 59322
rect 81046 59270 81098 59322
rect 81110 59270 81162 59322
rect 81174 59270 81226 59322
rect 81238 59270 81290 59322
rect 111766 59270 111818 59322
rect 111830 59270 111882 59322
rect 111894 59270 111946 59322
rect 111958 59270 112010 59322
rect 142486 59270 142538 59322
rect 142550 59270 142602 59322
rect 142614 59270 142666 59322
rect 142678 59270 142730 59322
rect 173206 59270 173258 59322
rect 173270 59270 173322 59322
rect 173334 59270 173386 59322
rect 173398 59270 173450 59322
rect 4246 58726 4298 58778
rect 4310 58726 4362 58778
rect 4374 58726 4426 58778
rect 4438 58726 4490 58778
rect 34966 58726 35018 58778
rect 35030 58726 35082 58778
rect 35094 58726 35146 58778
rect 35158 58726 35210 58778
rect 65686 58726 65738 58778
rect 65750 58726 65802 58778
rect 65814 58726 65866 58778
rect 65878 58726 65930 58778
rect 96406 58726 96458 58778
rect 96470 58726 96522 58778
rect 96534 58726 96586 58778
rect 96598 58726 96650 58778
rect 127126 58726 127178 58778
rect 127190 58726 127242 58778
rect 127254 58726 127306 58778
rect 127318 58726 127370 58778
rect 157846 58726 157898 58778
rect 157910 58726 157962 58778
rect 157974 58726 158026 58778
rect 158038 58726 158090 58778
rect 19606 58182 19658 58234
rect 19670 58182 19722 58234
rect 19734 58182 19786 58234
rect 19798 58182 19850 58234
rect 50326 58182 50378 58234
rect 50390 58182 50442 58234
rect 50454 58182 50506 58234
rect 50518 58182 50570 58234
rect 81046 58182 81098 58234
rect 81110 58182 81162 58234
rect 81174 58182 81226 58234
rect 81238 58182 81290 58234
rect 111766 58182 111818 58234
rect 111830 58182 111882 58234
rect 111894 58182 111946 58234
rect 111958 58182 112010 58234
rect 142486 58182 142538 58234
rect 142550 58182 142602 58234
rect 142614 58182 142666 58234
rect 142678 58182 142730 58234
rect 173206 58182 173258 58234
rect 173270 58182 173322 58234
rect 173334 58182 173386 58234
rect 173398 58182 173450 58234
rect 4246 57638 4298 57690
rect 4310 57638 4362 57690
rect 4374 57638 4426 57690
rect 4438 57638 4490 57690
rect 34966 57638 35018 57690
rect 35030 57638 35082 57690
rect 35094 57638 35146 57690
rect 35158 57638 35210 57690
rect 65686 57638 65738 57690
rect 65750 57638 65802 57690
rect 65814 57638 65866 57690
rect 65878 57638 65930 57690
rect 96406 57638 96458 57690
rect 96470 57638 96522 57690
rect 96534 57638 96586 57690
rect 96598 57638 96650 57690
rect 127126 57638 127178 57690
rect 127190 57638 127242 57690
rect 127254 57638 127306 57690
rect 127318 57638 127370 57690
rect 157846 57638 157898 57690
rect 157910 57638 157962 57690
rect 157974 57638 158026 57690
rect 158038 57638 158090 57690
rect 19606 57094 19658 57146
rect 19670 57094 19722 57146
rect 19734 57094 19786 57146
rect 19798 57094 19850 57146
rect 50326 57094 50378 57146
rect 50390 57094 50442 57146
rect 50454 57094 50506 57146
rect 50518 57094 50570 57146
rect 81046 57094 81098 57146
rect 81110 57094 81162 57146
rect 81174 57094 81226 57146
rect 81238 57094 81290 57146
rect 111766 57094 111818 57146
rect 111830 57094 111882 57146
rect 111894 57094 111946 57146
rect 111958 57094 112010 57146
rect 142486 57094 142538 57146
rect 142550 57094 142602 57146
rect 142614 57094 142666 57146
rect 142678 57094 142730 57146
rect 173206 57094 173258 57146
rect 173270 57094 173322 57146
rect 173334 57094 173386 57146
rect 173398 57094 173450 57146
rect 4246 56550 4298 56602
rect 4310 56550 4362 56602
rect 4374 56550 4426 56602
rect 4438 56550 4490 56602
rect 34966 56550 35018 56602
rect 35030 56550 35082 56602
rect 35094 56550 35146 56602
rect 35158 56550 35210 56602
rect 65686 56550 65738 56602
rect 65750 56550 65802 56602
rect 65814 56550 65866 56602
rect 65878 56550 65930 56602
rect 96406 56550 96458 56602
rect 96470 56550 96522 56602
rect 96534 56550 96586 56602
rect 96598 56550 96650 56602
rect 127126 56550 127178 56602
rect 127190 56550 127242 56602
rect 127254 56550 127306 56602
rect 127318 56550 127370 56602
rect 157846 56550 157898 56602
rect 157910 56550 157962 56602
rect 157974 56550 158026 56602
rect 158038 56550 158090 56602
rect 19606 56006 19658 56058
rect 19670 56006 19722 56058
rect 19734 56006 19786 56058
rect 19798 56006 19850 56058
rect 50326 56006 50378 56058
rect 50390 56006 50442 56058
rect 50454 56006 50506 56058
rect 50518 56006 50570 56058
rect 81046 56006 81098 56058
rect 81110 56006 81162 56058
rect 81174 56006 81226 56058
rect 81238 56006 81290 56058
rect 111766 56006 111818 56058
rect 111830 56006 111882 56058
rect 111894 56006 111946 56058
rect 111958 56006 112010 56058
rect 142486 56006 142538 56058
rect 142550 56006 142602 56058
rect 142614 56006 142666 56058
rect 142678 56006 142730 56058
rect 173206 56006 173258 56058
rect 173270 56006 173322 56058
rect 173334 56006 173386 56058
rect 173398 56006 173450 56058
rect 4246 55462 4298 55514
rect 4310 55462 4362 55514
rect 4374 55462 4426 55514
rect 4438 55462 4490 55514
rect 34966 55462 35018 55514
rect 35030 55462 35082 55514
rect 35094 55462 35146 55514
rect 35158 55462 35210 55514
rect 65686 55462 65738 55514
rect 65750 55462 65802 55514
rect 65814 55462 65866 55514
rect 65878 55462 65930 55514
rect 96406 55462 96458 55514
rect 96470 55462 96522 55514
rect 96534 55462 96586 55514
rect 96598 55462 96650 55514
rect 127126 55462 127178 55514
rect 127190 55462 127242 55514
rect 127254 55462 127306 55514
rect 127318 55462 127370 55514
rect 157846 55462 157898 55514
rect 157910 55462 157962 55514
rect 157974 55462 158026 55514
rect 158038 55462 158090 55514
rect 19606 54918 19658 54970
rect 19670 54918 19722 54970
rect 19734 54918 19786 54970
rect 19798 54918 19850 54970
rect 50326 54918 50378 54970
rect 50390 54918 50442 54970
rect 50454 54918 50506 54970
rect 50518 54918 50570 54970
rect 81046 54918 81098 54970
rect 81110 54918 81162 54970
rect 81174 54918 81226 54970
rect 81238 54918 81290 54970
rect 111766 54918 111818 54970
rect 111830 54918 111882 54970
rect 111894 54918 111946 54970
rect 111958 54918 112010 54970
rect 142486 54918 142538 54970
rect 142550 54918 142602 54970
rect 142614 54918 142666 54970
rect 142678 54918 142730 54970
rect 173206 54918 173258 54970
rect 173270 54918 173322 54970
rect 173334 54918 173386 54970
rect 173398 54918 173450 54970
rect 4246 54374 4298 54426
rect 4310 54374 4362 54426
rect 4374 54374 4426 54426
rect 4438 54374 4490 54426
rect 34966 54374 35018 54426
rect 35030 54374 35082 54426
rect 35094 54374 35146 54426
rect 35158 54374 35210 54426
rect 65686 54374 65738 54426
rect 65750 54374 65802 54426
rect 65814 54374 65866 54426
rect 65878 54374 65930 54426
rect 96406 54374 96458 54426
rect 96470 54374 96522 54426
rect 96534 54374 96586 54426
rect 96598 54374 96650 54426
rect 127126 54374 127178 54426
rect 127190 54374 127242 54426
rect 127254 54374 127306 54426
rect 127318 54374 127370 54426
rect 157846 54374 157898 54426
rect 157910 54374 157962 54426
rect 157974 54374 158026 54426
rect 158038 54374 158090 54426
rect 19606 53830 19658 53882
rect 19670 53830 19722 53882
rect 19734 53830 19786 53882
rect 19798 53830 19850 53882
rect 50326 53830 50378 53882
rect 50390 53830 50442 53882
rect 50454 53830 50506 53882
rect 50518 53830 50570 53882
rect 81046 53830 81098 53882
rect 81110 53830 81162 53882
rect 81174 53830 81226 53882
rect 81238 53830 81290 53882
rect 111766 53830 111818 53882
rect 111830 53830 111882 53882
rect 111894 53830 111946 53882
rect 111958 53830 112010 53882
rect 142486 53830 142538 53882
rect 142550 53830 142602 53882
rect 142614 53830 142666 53882
rect 142678 53830 142730 53882
rect 173206 53830 173258 53882
rect 173270 53830 173322 53882
rect 173334 53830 173386 53882
rect 173398 53830 173450 53882
rect 4246 53286 4298 53338
rect 4310 53286 4362 53338
rect 4374 53286 4426 53338
rect 4438 53286 4490 53338
rect 34966 53286 35018 53338
rect 35030 53286 35082 53338
rect 35094 53286 35146 53338
rect 35158 53286 35210 53338
rect 65686 53286 65738 53338
rect 65750 53286 65802 53338
rect 65814 53286 65866 53338
rect 65878 53286 65930 53338
rect 96406 53286 96458 53338
rect 96470 53286 96522 53338
rect 96534 53286 96586 53338
rect 96598 53286 96650 53338
rect 127126 53286 127178 53338
rect 127190 53286 127242 53338
rect 127254 53286 127306 53338
rect 127318 53286 127370 53338
rect 157846 53286 157898 53338
rect 157910 53286 157962 53338
rect 157974 53286 158026 53338
rect 158038 53286 158090 53338
rect 19606 52742 19658 52794
rect 19670 52742 19722 52794
rect 19734 52742 19786 52794
rect 19798 52742 19850 52794
rect 50326 52742 50378 52794
rect 50390 52742 50442 52794
rect 50454 52742 50506 52794
rect 50518 52742 50570 52794
rect 81046 52742 81098 52794
rect 81110 52742 81162 52794
rect 81174 52742 81226 52794
rect 81238 52742 81290 52794
rect 111766 52742 111818 52794
rect 111830 52742 111882 52794
rect 111894 52742 111946 52794
rect 111958 52742 112010 52794
rect 142486 52742 142538 52794
rect 142550 52742 142602 52794
rect 142614 52742 142666 52794
rect 142678 52742 142730 52794
rect 173206 52742 173258 52794
rect 173270 52742 173322 52794
rect 173334 52742 173386 52794
rect 173398 52742 173450 52794
rect 4246 52198 4298 52250
rect 4310 52198 4362 52250
rect 4374 52198 4426 52250
rect 4438 52198 4490 52250
rect 34966 52198 35018 52250
rect 35030 52198 35082 52250
rect 35094 52198 35146 52250
rect 35158 52198 35210 52250
rect 65686 52198 65738 52250
rect 65750 52198 65802 52250
rect 65814 52198 65866 52250
rect 65878 52198 65930 52250
rect 96406 52198 96458 52250
rect 96470 52198 96522 52250
rect 96534 52198 96586 52250
rect 96598 52198 96650 52250
rect 127126 52198 127178 52250
rect 127190 52198 127242 52250
rect 127254 52198 127306 52250
rect 127318 52198 127370 52250
rect 157846 52198 157898 52250
rect 157910 52198 157962 52250
rect 157974 52198 158026 52250
rect 158038 52198 158090 52250
rect 19606 51654 19658 51706
rect 19670 51654 19722 51706
rect 19734 51654 19786 51706
rect 19798 51654 19850 51706
rect 50326 51654 50378 51706
rect 50390 51654 50442 51706
rect 50454 51654 50506 51706
rect 50518 51654 50570 51706
rect 81046 51654 81098 51706
rect 81110 51654 81162 51706
rect 81174 51654 81226 51706
rect 81238 51654 81290 51706
rect 111766 51654 111818 51706
rect 111830 51654 111882 51706
rect 111894 51654 111946 51706
rect 111958 51654 112010 51706
rect 142486 51654 142538 51706
rect 142550 51654 142602 51706
rect 142614 51654 142666 51706
rect 142678 51654 142730 51706
rect 173206 51654 173258 51706
rect 173270 51654 173322 51706
rect 173334 51654 173386 51706
rect 173398 51654 173450 51706
rect 4246 51110 4298 51162
rect 4310 51110 4362 51162
rect 4374 51110 4426 51162
rect 4438 51110 4490 51162
rect 34966 51110 35018 51162
rect 35030 51110 35082 51162
rect 35094 51110 35146 51162
rect 35158 51110 35210 51162
rect 65686 51110 65738 51162
rect 65750 51110 65802 51162
rect 65814 51110 65866 51162
rect 65878 51110 65930 51162
rect 96406 51110 96458 51162
rect 96470 51110 96522 51162
rect 96534 51110 96586 51162
rect 96598 51110 96650 51162
rect 127126 51110 127178 51162
rect 127190 51110 127242 51162
rect 127254 51110 127306 51162
rect 127318 51110 127370 51162
rect 157846 51110 157898 51162
rect 157910 51110 157962 51162
rect 157974 51110 158026 51162
rect 158038 51110 158090 51162
rect 19606 50566 19658 50618
rect 19670 50566 19722 50618
rect 19734 50566 19786 50618
rect 19798 50566 19850 50618
rect 50326 50566 50378 50618
rect 50390 50566 50442 50618
rect 50454 50566 50506 50618
rect 50518 50566 50570 50618
rect 81046 50566 81098 50618
rect 81110 50566 81162 50618
rect 81174 50566 81226 50618
rect 81238 50566 81290 50618
rect 111766 50566 111818 50618
rect 111830 50566 111882 50618
rect 111894 50566 111946 50618
rect 111958 50566 112010 50618
rect 142486 50566 142538 50618
rect 142550 50566 142602 50618
rect 142614 50566 142666 50618
rect 142678 50566 142730 50618
rect 173206 50566 173258 50618
rect 173270 50566 173322 50618
rect 173334 50566 173386 50618
rect 173398 50566 173450 50618
rect 4246 50022 4298 50074
rect 4310 50022 4362 50074
rect 4374 50022 4426 50074
rect 4438 50022 4490 50074
rect 34966 50022 35018 50074
rect 35030 50022 35082 50074
rect 35094 50022 35146 50074
rect 35158 50022 35210 50074
rect 65686 50022 65738 50074
rect 65750 50022 65802 50074
rect 65814 50022 65866 50074
rect 65878 50022 65930 50074
rect 96406 50022 96458 50074
rect 96470 50022 96522 50074
rect 96534 50022 96586 50074
rect 96598 50022 96650 50074
rect 127126 50022 127178 50074
rect 127190 50022 127242 50074
rect 127254 50022 127306 50074
rect 127318 50022 127370 50074
rect 157846 50022 157898 50074
rect 157910 50022 157962 50074
rect 157974 50022 158026 50074
rect 158038 50022 158090 50074
rect 19606 49478 19658 49530
rect 19670 49478 19722 49530
rect 19734 49478 19786 49530
rect 19798 49478 19850 49530
rect 50326 49478 50378 49530
rect 50390 49478 50442 49530
rect 50454 49478 50506 49530
rect 50518 49478 50570 49530
rect 81046 49478 81098 49530
rect 81110 49478 81162 49530
rect 81174 49478 81226 49530
rect 81238 49478 81290 49530
rect 111766 49478 111818 49530
rect 111830 49478 111882 49530
rect 111894 49478 111946 49530
rect 111958 49478 112010 49530
rect 142486 49478 142538 49530
rect 142550 49478 142602 49530
rect 142614 49478 142666 49530
rect 142678 49478 142730 49530
rect 173206 49478 173258 49530
rect 173270 49478 173322 49530
rect 173334 49478 173386 49530
rect 173398 49478 173450 49530
rect 4246 48934 4298 48986
rect 4310 48934 4362 48986
rect 4374 48934 4426 48986
rect 4438 48934 4490 48986
rect 34966 48934 35018 48986
rect 35030 48934 35082 48986
rect 35094 48934 35146 48986
rect 35158 48934 35210 48986
rect 65686 48934 65738 48986
rect 65750 48934 65802 48986
rect 65814 48934 65866 48986
rect 65878 48934 65930 48986
rect 96406 48934 96458 48986
rect 96470 48934 96522 48986
rect 96534 48934 96586 48986
rect 96598 48934 96650 48986
rect 127126 48934 127178 48986
rect 127190 48934 127242 48986
rect 127254 48934 127306 48986
rect 127318 48934 127370 48986
rect 157846 48934 157898 48986
rect 157910 48934 157962 48986
rect 157974 48934 158026 48986
rect 158038 48934 158090 48986
rect 19606 48390 19658 48442
rect 19670 48390 19722 48442
rect 19734 48390 19786 48442
rect 19798 48390 19850 48442
rect 50326 48390 50378 48442
rect 50390 48390 50442 48442
rect 50454 48390 50506 48442
rect 50518 48390 50570 48442
rect 81046 48390 81098 48442
rect 81110 48390 81162 48442
rect 81174 48390 81226 48442
rect 81238 48390 81290 48442
rect 111766 48390 111818 48442
rect 111830 48390 111882 48442
rect 111894 48390 111946 48442
rect 111958 48390 112010 48442
rect 142486 48390 142538 48442
rect 142550 48390 142602 48442
rect 142614 48390 142666 48442
rect 142678 48390 142730 48442
rect 173206 48390 173258 48442
rect 173270 48390 173322 48442
rect 173334 48390 173386 48442
rect 173398 48390 173450 48442
rect 4246 47846 4298 47898
rect 4310 47846 4362 47898
rect 4374 47846 4426 47898
rect 4438 47846 4490 47898
rect 34966 47846 35018 47898
rect 35030 47846 35082 47898
rect 35094 47846 35146 47898
rect 35158 47846 35210 47898
rect 65686 47846 65738 47898
rect 65750 47846 65802 47898
rect 65814 47846 65866 47898
rect 65878 47846 65930 47898
rect 96406 47846 96458 47898
rect 96470 47846 96522 47898
rect 96534 47846 96586 47898
rect 96598 47846 96650 47898
rect 127126 47846 127178 47898
rect 127190 47846 127242 47898
rect 127254 47846 127306 47898
rect 127318 47846 127370 47898
rect 157846 47846 157898 47898
rect 157910 47846 157962 47898
rect 157974 47846 158026 47898
rect 158038 47846 158090 47898
rect 19606 47302 19658 47354
rect 19670 47302 19722 47354
rect 19734 47302 19786 47354
rect 19798 47302 19850 47354
rect 50326 47302 50378 47354
rect 50390 47302 50442 47354
rect 50454 47302 50506 47354
rect 50518 47302 50570 47354
rect 81046 47302 81098 47354
rect 81110 47302 81162 47354
rect 81174 47302 81226 47354
rect 81238 47302 81290 47354
rect 111766 47302 111818 47354
rect 111830 47302 111882 47354
rect 111894 47302 111946 47354
rect 111958 47302 112010 47354
rect 142486 47302 142538 47354
rect 142550 47302 142602 47354
rect 142614 47302 142666 47354
rect 142678 47302 142730 47354
rect 173206 47302 173258 47354
rect 173270 47302 173322 47354
rect 173334 47302 173386 47354
rect 173398 47302 173450 47354
rect 4246 46758 4298 46810
rect 4310 46758 4362 46810
rect 4374 46758 4426 46810
rect 4438 46758 4490 46810
rect 34966 46758 35018 46810
rect 35030 46758 35082 46810
rect 35094 46758 35146 46810
rect 35158 46758 35210 46810
rect 65686 46758 65738 46810
rect 65750 46758 65802 46810
rect 65814 46758 65866 46810
rect 65878 46758 65930 46810
rect 96406 46758 96458 46810
rect 96470 46758 96522 46810
rect 96534 46758 96586 46810
rect 96598 46758 96650 46810
rect 127126 46758 127178 46810
rect 127190 46758 127242 46810
rect 127254 46758 127306 46810
rect 127318 46758 127370 46810
rect 157846 46758 157898 46810
rect 157910 46758 157962 46810
rect 157974 46758 158026 46810
rect 158038 46758 158090 46810
rect 19606 46214 19658 46266
rect 19670 46214 19722 46266
rect 19734 46214 19786 46266
rect 19798 46214 19850 46266
rect 50326 46214 50378 46266
rect 50390 46214 50442 46266
rect 50454 46214 50506 46266
rect 50518 46214 50570 46266
rect 81046 46214 81098 46266
rect 81110 46214 81162 46266
rect 81174 46214 81226 46266
rect 81238 46214 81290 46266
rect 111766 46214 111818 46266
rect 111830 46214 111882 46266
rect 111894 46214 111946 46266
rect 111958 46214 112010 46266
rect 142486 46214 142538 46266
rect 142550 46214 142602 46266
rect 142614 46214 142666 46266
rect 142678 46214 142730 46266
rect 173206 46214 173258 46266
rect 173270 46214 173322 46266
rect 173334 46214 173386 46266
rect 173398 46214 173450 46266
rect 4246 45670 4298 45722
rect 4310 45670 4362 45722
rect 4374 45670 4426 45722
rect 4438 45670 4490 45722
rect 34966 45670 35018 45722
rect 35030 45670 35082 45722
rect 35094 45670 35146 45722
rect 35158 45670 35210 45722
rect 65686 45670 65738 45722
rect 65750 45670 65802 45722
rect 65814 45670 65866 45722
rect 65878 45670 65930 45722
rect 96406 45670 96458 45722
rect 96470 45670 96522 45722
rect 96534 45670 96586 45722
rect 96598 45670 96650 45722
rect 127126 45670 127178 45722
rect 127190 45670 127242 45722
rect 127254 45670 127306 45722
rect 127318 45670 127370 45722
rect 157846 45670 157898 45722
rect 157910 45670 157962 45722
rect 157974 45670 158026 45722
rect 158038 45670 158090 45722
rect 19606 45126 19658 45178
rect 19670 45126 19722 45178
rect 19734 45126 19786 45178
rect 19798 45126 19850 45178
rect 50326 45126 50378 45178
rect 50390 45126 50442 45178
rect 50454 45126 50506 45178
rect 50518 45126 50570 45178
rect 81046 45126 81098 45178
rect 81110 45126 81162 45178
rect 81174 45126 81226 45178
rect 81238 45126 81290 45178
rect 111766 45126 111818 45178
rect 111830 45126 111882 45178
rect 111894 45126 111946 45178
rect 111958 45126 112010 45178
rect 142486 45126 142538 45178
rect 142550 45126 142602 45178
rect 142614 45126 142666 45178
rect 142678 45126 142730 45178
rect 173206 45126 173258 45178
rect 173270 45126 173322 45178
rect 173334 45126 173386 45178
rect 173398 45126 173450 45178
rect 4246 44582 4298 44634
rect 4310 44582 4362 44634
rect 4374 44582 4426 44634
rect 4438 44582 4490 44634
rect 34966 44582 35018 44634
rect 35030 44582 35082 44634
rect 35094 44582 35146 44634
rect 35158 44582 35210 44634
rect 65686 44582 65738 44634
rect 65750 44582 65802 44634
rect 65814 44582 65866 44634
rect 65878 44582 65930 44634
rect 96406 44582 96458 44634
rect 96470 44582 96522 44634
rect 96534 44582 96586 44634
rect 96598 44582 96650 44634
rect 127126 44582 127178 44634
rect 127190 44582 127242 44634
rect 127254 44582 127306 44634
rect 127318 44582 127370 44634
rect 157846 44582 157898 44634
rect 157910 44582 157962 44634
rect 157974 44582 158026 44634
rect 158038 44582 158090 44634
rect 19606 44038 19658 44090
rect 19670 44038 19722 44090
rect 19734 44038 19786 44090
rect 19798 44038 19850 44090
rect 50326 44038 50378 44090
rect 50390 44038 50442 44090
rect 50454 44038 50506 44090
rect 50518 44038 50570 44090
rect 81046 44038 81098 44090
rect 81110 44038 81162 44090
rect 81174 44038 81226 44090
rect 81238 44038 81290 44090
rect 111766 44038 111818 44090
rect 111830 44038 111882 44090
rect 111894 44038 111946 44090
rect 111958 44038 112010 44090
rect 142486 44038 142538 44090
rect 142550 44038 142602 44090
rect 142614 44038 142666 44090
rect 142678 44038 142730 44090
rect 173206 44038 173258 44090
rect 173270 44038 173322 44090
rect 173334 44038 173386 44090
rect 173398 44038 173450 44090
rect 4246 43494 4298 43546
rect 4310 43494 4362 43546
rect 4374 43494 4426 43546
rect 4438 43494 4490 43546
rect 34966 43494 35018 43546
rect 35030 43494 35082 43546
rect 35094 43494 35146 43546
rect 35158 43494 35210 43546
rect 65686 43494 65738 43546
rect 65750 43494 65802 43546
rect 65814 43494 65866 43546
rect 65878 43494 65930 43546
rect 96406 43494 96458 43546
rect 96470 43494 96522 43546
rect 96534 43494 96586 43546
rect 96598 43494 96650 43546
rect 127126 43494 127178 43546
rect 127190 43494 127242 43546
rect 127254 43494 127306 43546
rect 127318 43494 127370 43546
rect 157846 43494 157898 43546
rect 157910 43494 157962 43546
rect 157974 43494 158026 43546
rect 158038 43494 158090 43546
rect 19606 42950 19658 43002
rect 19670 42950 19722 43002
rect 19734 42950 19786 43002
rect 19798 42950 19850 43002
rect 50326 42950 50378 43002
rect 50390 42950 50442 43002
rect 50454 42950 50506 43002
rect 50518 42950 50570 43002
rect 81046 42950 81098 43002
rect 81110 42950 81162 43002
rect 81174 42950 81226 43002
rect 81238 42950 81290 43002
rect 111766 42950 111818 43002
rect 111830 42950 111882 43002
rect 111894 42950 111946 43002
rect 111958 42950 112010 43002
rect 142486 42950 142538 43002
rect 142550 42950 142602 43002
rect 142614 42950 142666 43002
rect 142678 42950 142730 43002
rect 173206 42950 173258 43002
rect 173270 42950 173322 43002
rect 173334 42950 173386 43002
rect 173398 42950 173450 43002
rect 4246 42406 4298 42458
rect 4310 42406 4362 42458
rect 4374 42406 4426 42458
rect 4438 42406 4490 42458
rect 34966 42406 35018 42458
rect 35030 42406 35082 42458
rect 35094 42406 35146 42458
rect 35158 42406 35210 42458
rect 65686 42406 65738 42458
rect 65750 42406 65802 42458
rect 65814 42406 65866 42458
rect 65878 42406 65930 42458
rect 96406 42406 96458 42458
rect 96470 42406 96522 42458
rect 96534 42406 96586 42458
rect 96598 42406 96650 42458
rect 127126 42406 127178 42458
rect 127190 42406 127242 42458
rect 127254 42406 127306 42458
rect 127318 42406 127370 42458
rect 157846 42406 157898 42458
rect 157910 42406 157962 42458
rect 157974 42406 158026 42458
rect 158038 42406 158090 42458
rect 19606 41862 19658 41914
rect 19670 41862 19722 41914
rect 19734 41862 19786 41914
rect 19798 41862 19850 41914
rect 50326 41862 50378 41914
rect 50390 41862 50442 41914
rect 50454 41862 50506 41914
rect 50518 41862 50570 41914
rect 81046 41862 81098 41914
rect 81110 41862 81162 41914
rect 81174 41862 81226 41914
rect 81238 41862 81290 41914
rect 111766 41862 111818 41914
rect 111830 41862 111882 41914
rect 111894 41862 111946 41914
rect 111958 41862 112010 41914
rect 142486 41862 142538 41914
rect 142550 41862 142602 41914
rect 142614 41862 142666 41914
rect 142678 41862 142730 41914
rect 173206 41862 173258 41914
rect 173270 41862 173322 41914
rect 173334 41862 173386 41914
rect 173398 41862 173450 41914
rect 4246 41318 4298 41370
rect 4310 41318 4362 41370
rect 4374 41318 4426 41370
rect 4438 41318 4490 41370
rect 34966 41318 35018 41370
rect 35030 41318 35082 41370
rect 35094 41318 35146 41370
rect 35158 41318 35210 41370
rect 65686 41318 65738 41370
rect 65750 41318 65802 41370
rect 65814 41318 65866 41370
rect 65878 41318 65930 41370
rect 96406 41318 96458 41370
rect 96470 41318 96522 41370
rect 96534 41318 96586 41370
rect 96598 41318 96650 41370
rect 127126 41318 127178 41370
rect 127190 41318 127242 41370
rect 127254 41318 127306 41370
rect 127318 41318 127370 41370
rect 157846 41318 157898 41370
rect 157910 41318 157962 41370
rect 157974 41318 158026 41370
rect 158038 41318 158090 41370
rect 19606 40774 19658 40826
rect 19670 40774 19722 40826
rect 19734 40774 19786 40826
rect 19798 40774 19850 40826
rect 50326 40774 50378 40826
rect 50390 40774 50442 40826
rect 50454 40774 50506 40826
rect 50518 40774 50570 40826
rect 81046 40774 81098 40826
rect 81110 40774 81162 40826
rect 81174 40774 81226 40826
rect 81238 40774 81290 40826
rect 111766 40774 111818 40826
rect 111830 40774 111882 40826
rect 111894 40774 111946 40826
rect 111958 40774 112010 40826
rect 142486 40774 142538 40826
rect 142550 40774 142602 40826
rect 142614 40774 142666 40826
rect 142678 40774 142730 40826
rect 173206 40774 173258 40826
rect 173270 40774 173322 40826
rect 173334 40774 173386 40826
rect 173398 40774 173450 40826
rect 4246 40230 4298 40282
rect 4310 40230 4362 40282
rect 4374 40230 4426 40282
rect 4438 40230 4490 40282
rect 34966 40230 35018 40282
rect 35030 40230 35082 40282
rect 35094 40230 35146 40282
rect 35158 40230 35210 40282
rect 65686 40230 65738 40282
rect 65750 40230 65802 40282
rect 65814 40230 65866 40282
rect 65878 40230 65930 40282
rect 96406 40230 96458 40282
rect 96470 40230 96522 40282
rect 96534 40230 96586 40282
rect 96598 40230 96650 40282
rect 127126 40230 127178 40282
rect 127190 40230 127242 40282
rect 127254 40230 127306 40282
rect 127318 40230 127370 40282
rect 157846 40230 157898 40282
rect 157910 40230 157962 40282
rect 157974 40230 158026 40282
rect 158038 40230 158090 40282
rect 19606 39686 19658 39738
rect 19670 39686 19722 39738
rect 19734 39686 19786 39738
rect 19798 39686 19850 39738
rect 50326 39686 50378 39738
rect 50390 39686 50442 39738
rect 50454 39686 50506 39738
rect 50518 39686 50570 39738
rect 81046 39686 81098 39738
rect 81110 39686 81162 39738
rect 81174 39686 81226 39738
rect 81238 39686 81290 39738
rect 111766 39686 111818 39738
rect 111830 39686 111882 39738
rect 111894 39686 111946 39738
rect 111958 39686 112010 39738
rect 142486 39686 142538 39738
rect 142550 39686 142602 39738
rect 142614 39686 142666 39738
rect 142678 39686 142730 39738
rect 173206 39686 173258 39738
rect 173270 39686 173322 39738
rect 173334 39686 173386 39738
rect 173398 39686 173450 39738
rect 4246 39142 4298 39194
rect 4310 39142 4362 39194
rect 4374 39142 4426 39194
rect 4438 39142 4490 39194
rect 34966 39142 35018 39194
rect 35030 39142 35082 39194
rect 35094 39142 35146 39194
rect 35158 39142 35210 39194
rect 65686 39142 65738 39194
rect 65750 39142 65802 39194
rect 65814 39142 65866 39194
rect 65878 39142 65930 39194
rect 96406 39142 96458 39194
rect 96470 39142 96522 39194
rect 96534 39142 96586 39194
rect 96598 39142 96650 39194
rect 127126 39142 127178 39194
rect 127190 39142 127242 39194
rect 127254 39142 127306 39194
rect 127318 39142 127370 39194
rect 157846 39142 157898 39194
rect 157910 39142 157962 39194
rect 157974 39142 158026 39194
rect 158038 39142 158090 39194
rect 19606 38598 19658 38650
rect 19670 38598 19722 38650
rect 19734 38598 19786 38650
rect 19798 38598 19850 38650
rect 50326 38598 50378 38650
rect 50390 38598 50442 38650
rect 50454 38598 50506 38650
rect 50518 38598 50570 38650
rect 81046 38598 81098 38650
rect 81110 38598 81162 38650
rect 81174 38598 81226 38650
rect 81238 38598 81290 38650
rect 111766 38598 111818 38650
rect 111830 38598 111882 38650
rect 111894 38598 111946 38650
rect 111958 38598 112010 38650
rect 142486 38598 142538 38650
rect 142550 38598 142602 38650
rect 142614 38598 142666 38650
rect 142678 38598 142730 38650
rect 173206 38598 173258 38650
rect 173270 38598 173322 38650
rect 173334 38598 173386 38650
rect 173398 38598 173450 38650
rect 4246 38054 4298 38106
rect 4310 38054 4362 38106
rect 4374 38054 4426 38106
rect 4438 38054 4490 38106
rect 34966 38054 35018 38106
rect 35030 38054 35082 38106
rect 35094 38054 35146 38106
rect 35158 38054 35210 38106
rect 65686 38054 65738 38106
rect 65750 38054 65802 38106
rect 65814 38054 65866 38106
rect 65878 38054 65930 38106
rect 96406 38054 96458 38106
rect 96470 38054 96522 38106
rect 96534 38054 96586 38106
rect 96598 38054 96650 38106
rect 127126 38054 127178 38106
rect 127190 38054 127242 38106
rect 127254 38054 127306 38106
rect 127318 38054 127370 38106
rect 157846 38054 157898 38106
rect 157910 38054 157962 38106
rect 157974 38054 158026 38106
rect 158038 38054 158090 38106
rect 19606 37510 19658 37562
rect 19670 37510 19722 37562
rect 19734 37510 19786 37562
rect 19798 37510 19850 37562
rect 50326 37510 50378 37562
rect 50390 37510 50442 37562
rect 50454 37510 50506 37562
rect 50518 37510 50570 37562
rect 81046 37510 81098 37562
rect 81110 37510 81162 37562
rect 81174 37510 81226 37562
rect 81238 37510 81290 37562
rect 111766 37510 111818 37562
rect 111830 37510 111882 37562
rect 111894 37510 111946 37562
rect 111958 37510 112010 37562
rect 142486 37510 142538 37562
rect 142550 37510 142602 37562
rect 142614 37510 142666 37562
rect 142678 37510 142730 37562
rect 173206 37510 173258 37562
rect 173270 37510 173322 37562
rect 173334 37510 173386 37562
rect 173398 37510 173450 37562
rect 4246 36966 4298 37018
rect 4310 36966 4362 37018
rect 4374 36966 4426 37018
rect 4438 36966 4490 37018
rect 34966 36966 35018 37018
rect 35030 36966 35082 37018
rect 35094 36966 35146 37018
rect 35158 36966 35210 37018
rect 65686 36966 65738 37018
rect 65750 36966 65802 37018
rect 65814 36966 65866 37018
rect 65878 36966 65930 37018
rect 96406 36966 96458 37018
rect 96470 36966 96522 37018
rect 96534 36966 96586 37018
rect 96598 36966 96650 37018
rect 127126 36966 127178 37018
rect 127190 36966 127242 37018
rect 127254 36966 127306 37018
rect 127318 36966 127370 37018
rect 157846 36966 157898 37018
rect 157910 36966 157962 37018
rect 157974 36966 158026 37018
rect 158038 36966 158090 37018
rect 19606 36422 19658 36474
rect 19670 36422 19722 36474
rect 19734 36422 19786 36474
rect 19798 36422 19850 36474
rect 50326 36422 50378 36474
rect 50390 36422 50442 36474
rect 50454 36422 50506 36474
rect 50518 36422 50570 36474
rect 81046 36422 81098 36474
rect 81110 36422 81162 36474
rect 81174 36422 81226 36474
rect 81238 36422 81290 36474
rect 111766 36422 111818 36474
rect 111830 36422 111882 36474
rect 111894 36422 111946 36474
rect 111958 36422 112010 36474
rect 142486 36422 142538 36474
rect 142550 36422 142602 36474
rect 142614 36422 142666 36474
rect 142678 36422 142730 36474
rect 173206 36422 173258 36474
rect 173270 36422 173322 36474
rect 173334 36422 173386 36474
rect 173398 36422 173450 36474
rect 4246 35878 4298 35930
rect 4310 35878 4362 35930
rect 4374 35878 4426 35930
rect 4438 35878 4490 35930
rect 34966 35878 35018 35930
rect 35030 35878 35082 35930
rect 35094 35878 35146 35930
rect 35158 35878 35210 35930
rect 65686 35878 65738 35930
rect 65750 35878 65802 35930
rect 65814 35878 65866 35930
rect 65878 35878 65930 35930
rect 96406 35878 96458 35930
rect 96470 35878 96522 35930
rect 96534 35878 96586 35930
rect 96598 35878 96650 35930
rect 127126 35878 127178 35930
rect 127190 35878 127242 35930
rect 127254 35878 127306 35930
rect 127318 35878 127370 35930
rect 157846 35878 157898 35930
rect 157910 35878 157962 35930
rect 157974 35878 158026 35930
rect 158038 35878 158090 35930
rect 19606 35334 19658 35386
rect 19670 35334 19722 35386
rect 19734 35334 19786 35386
rect 19798 35334 19850 35386
rect 50326 35334 50378 35386
rect 50390 35334 50442 35386
rect 50454 35334 50506 35386
rect 50518 35334 50570 35386
rect 81046 35334 81098 35386
rect 81110 35334 81162 35386
rect 81174 35334 81226 35386
rect 81238 35334 81290 35386
rect 111766 35334 111818 35386
rect 111830 35334 111882 35386
rect 111894 35334 111946 35386
rect 111958 35334 112010 35386
rect 142486 35334 142538 35386
rect 142550 35334 142602 35386
rect 142614 35334 142666 35386
rect 142678 35334 142730 35386
rect 173206 35334 173258 35386
rect 173270 35334 173322 35386
rect 173334 35334 173386 35386
rect 173398 35334 173450 35386
rect 4246 34790 4298 34842
rect 4310 34790 4362 34842
rect 4374 34790 4426 34842
rect 4438 34790 4490 34842
rect 34966 34790 35018 34842
rect 35030 34790 35082 34842
rect 35094 34790 35146 34842
rect 35158 34790 35210 34842
rect 65686 34790 65738 34842
rect 65750 34790 65802 34842
rect 65814 34790 65866 34842
rect 65878 34790 65930 34842
rect 96406 34790 96458 34842
rect 96470 34790 96522 34842
rect 96534 34790 96586 34842
rect 96598 34790 96650 34842
rect 127126 34790 127178 34842
rect 127190 34790 127242 34842
rect 127254 34790 127306 34842
rect 127318 34790 127370 34842
rect 157846 34790 157898 34842
rect 157910 34790 157962 34842
rect 157974 34790 158026 34842
rect 158038 34790 158090 34842
rect 19606 34246 19658 34298
rect 19670 34246 19722 34298
rect 19734 34246 19786 34298
rect 19798 34246 19850 34298
rect 50326 34246 50378 34298
rect 50390 34246 50442 34298
rect 50454 34246 50506 34298
rect 50518 34246 50570 34298
rect 81046 34246 81098 34298
rect 81110 34246 81162 34298
rect 81174 34246 81226 34298
rect 81238 34246 81290 34298
rect 111766 34246 111818 34298
rect 111830 34246 111882 34298
rect 111894 34246 111946 34298
rect 111958 34246 112010 34298
rect 142486 34246 142538 34298
rect 142550 34246 142602 34298
rect 142614 34246 142666 34298
rect 142678 34246 142730 34298
rect 173206 34246 173258 34298
rect 173270 34246 173322 34298
rect 173334 34246 173386 34298
rect 173398 34246 173450 34298
rect 4246 33702 4298 33754
rect 4310 33702 4362 33754
rect 4374 33702 4426 33754
rect 4438 33702 4490 33754
rect 34966 33702 35018 33754
rect 35030 33702 35082 33754
rect 35094 33702 35146 33754
rect 35158 33702 35210 33754
rect 65686 33702 65738 33754
rect 65750 33702 65802 33754
rect 65814 33702 65866 33754
rect 65878 33702 65930 33754
rect 96406 33702 96458 33754
rect 96470 33702 96522 33754
rect 96534 33702 96586 33754
rect 96598 33702 96650 33754
rect 127126 33702 127178 33754
rect 127190 33702 127242 33754
rect 127254 33702 127306 33754
rect 127318 33702 127370 33754
rect 157846 33702 157898 33754
rect 157910 33702 157962 33754
rect 157974 33702 158026 33754
rect 158038 33702 158090 33754
rect 19606 33158 19658 33210
rect 19670 33158 19722 33210
rect 19734 33158 19786 33210
rect 19798 33158 19850 33210
rect 50326 33158 50378 33210
rect 50390 33158 50442 33210
rect 50454 33158 50506 33210
rect 50518 33158 50570 33210
rect 81046 33158 81098 33210
rect 81110 33158 81162 33210
rect 81174 33158 81226 33210
rect 81238 33158 81290 33210
rect 111766 33158 111818 33210
rect 111830 33158 111882 33210
rect 111894 33158 111946 33210
rect 111958 33158 112010 33210
rect 142486 33158 142538 33210
rect 142550 33158 142602 33210
rect 142614 33158 142666 33210
rect 142678 33158 142730 33210
rect 173206 33158 173258 33210
rect 173270 33158 173322 33210
rect 173334 33158 173386 33210
rect 173398 33158 173450 33210
rect 4246 32614 4298 32666
rect 4310 32614 4362 32666
rect 4374 32614 4426 32666
rect 4438 32614 4490 32666
rect 34966 32614 35018 32666
rect 35030 32614 35082 32666
rect 35094 32614 35146 32666
rect 35158 32614 35210 32666
rect 65686 32614 65738 32666
rect 65750 32614 65802 32666
rect 65814 32614 65866 32666
rect 65878 32614 65930 32666
rect 96406 32614 96458 32666
rect 96470 32614 96522 32666
rect 96534 32614 96586 32666
rect 96598 32614 96650 32666
rect 127126 32614 127178 32666
rect 127190 32614 127242 32666
rect 127254 32614 127306 32666
rect 127318 32614 127370 32666
rect 157846 32614 157898 32666
rect 157910 32614 157962 32666
rect 157974 32614 158026 32666
rect 158038 32614 158090 32666
rect 19606 32070 19658 32122
rect 19670 32070 19722 32122
rect 19734 32070 19786 32122
rect 19798 32070 19850 32122
rect 50326 32070 50378 32122
rect 50390 32070 50442 32122
rect 50454 32070 50506 32122
rect 50518 32070 50570 32122
rect 81046 32070 81098 32122
rect 81110 32070 81162 32122
rect 81174 32070 81226 32122
rect 81238 32070 81290 32122
rect 111766 32070 111818 32122
rect 111830 32070 111882 32122
rect 111894 32070 111946 32122
rect 111958 32070 112010 32122
rect 142486 32070 142538 32122
rect 142550 32070 142602 32122
rect 142614 32070 142666 32122
rect 142678 32070 142730 32122
rect 173206 32070 173258 32122
rect 173270 32070 173322 32122
rect 173334 32070 173386 32122
rect 173398 32070 173450 32122
rect 4246 31526 4298 31578
rect 4310 31526 4362 31578
rect 4374 31526 4426 31578
rect 4438 31526 4490 31578
rect 34966 31526 35018 31578
rect 35030 31526 35082 31578
rect 35094 31526 35146 31578
rect 35158 31526 35210 31578
rect 65686 31526 65738 31578
rect 65750 31526 65802 31578
rect 65814 31526 65866 31578
rect 65878 31526 65930 31578
rect 96406 31526 96458 31578
rect 96470 31526 96522 31578
rect 96534 31526 96586 31578
rect 96598 31526 96650 31578
rect 127126 31526 127178 31578
rect 127190 31526 127242 31578
rect 127254 31526 127306 31578
rect 127318 31526 127370 31578
rect 157846 31526 157898 31578
rect 157910 31526 157962 31578
rect 157974 31526 158026 31578
rect 158038 31526 158090 31578
rect 19606 30982 19658 31034
rect 19670 30982 19722 31034
rect 19734 30982 19786 31034
rect 19798 30982 19850 31034
rect 50326 30982 50378 31034
rect 50390 30982 50442 31034
rect 50454 30982 50506 31034
rect 50518 30982 50570 31034
rect 81046 30982 81098 31034
rect 81110 30982 81162 31034
rect 81174 30982 81226 31034
rect 81238 30982 81290 31034
rect 111766 30982 111818 31034
rect 111830 30982 111882 31034
rect 111894 30982 111946 31034
rect 111958 30982 112010 31034
rect 142486 30982 142538 31034
rect 142550 30982 142602 31034
rect 142614 30982 142666 31034
rect 142678 30982 142730 31034
rect 173206 30982 173258 31034
rect 173270 30982 173322 31034
rect 173334 30982 173386 31034
rect 173398 30982 173450 31034
rect 4246 30438 4298 30490
rect 4310 30438 4362 30490
rect 4374 30438 4426 30490
rect 4438 30438 4490 30490
rect 34966 30438 35018 30490
rect 35030 30438 35082 30490
rect 35094 30438 35146 30490
rect 35158 30438 35210 30490
rect 65686 30438 65738 30490
rect 65750 30438 65802 30490
rect 65814 30438 65866 30490
rect 65878 30438 65930 30490
rect 96406 30438 96458 30490
rect 96470 30438 96522 30490
rect 96534 30438 96586 30490
rect 96598 30438 96650 30490
rect 127126 30438 127178 30490
rect 127190 30438 127242 30490
rect 127254 30438 127306 30490
rect 127318 30438 127370 30490
rect 157846 30438 157898 30490
rect 157910 30438 157962 30490
rect 157974 30438 158026 30490
rect 158038 30438 158090 30490
rect 19606 29894 19658 29946
rect 19670 29894 19722 29946
rect 19734 29894 19786 29946
rect 19798 29894 19850 29946
rect 50326 29894 50378 29946
rect 50390 29894 50442 29946
rect 50454 29894 50506 29946
rect 50518 29894 50570 29946
rect 81046 29894 81098 29946
rect 81110 29894 81162 29946
rect 81174 29894 81226 29946
rect 81238 29894 81290 29946
rect 111766 29894 111818 29946
rect 111830 29894 111882 29946
rect 111894 29894 111946 29946
rect 111958 29894 112010 29946
rect 142486 29894 142538 29946
rect 142550 29894 142602 29946
rect 142614 29894 142666 29946
rect 142678 29894 142730 29946
rect 173206 29894 173258 29946
rect 173270 29894 173322 29946
rect 173334 29894 173386 29946
rect 173398 29894 173450 29946
rect 4246 29350 4298 29402
rect 4310 29350 4362 29402
rect 4374 29350 4426 29402
rect 4438 29350 4490 29402
rect 34966 29350 35018 29402
rect 35030 29350 35082 29402
rect 35094 29350 35146 29402
rect 35158 29350 35210 29402
rect 65686 29350 65738 29402
rect 65750 29350 65802 29402
rect 65814 29350 65866 29402
rect 65878 29350 65930 29402
rect 96406 29350 96458 29402
rect 96470 29350 96522 29402
rect 96534 29350 96586 29402
rect 96598 29350 96650 29402
rect 127126 29350 127178 29402
rect 127190 29350 127242 29402
rect 127254 29350 127306 29402
rect 127318 29350 127370 29402
rect 157846 29350 157898 29402
rect 157910 29350 157962 29402
rect 157974 29350 158026 29402
rect 158038 29350 158090 29402
rect 19606 28806 19658 28858
rect 19670 28806 19722 28858
rect 19734 28806 19786 28858
rect 19798 28806 19850 28858
rect 50326 28806 50378 28858
rect 50390 28806 50442 28858
rect 50454 28806 50506 28858
rect 50518 28806 50570 28858
rect 81046 28806 81098 28858
rect 81110 28806 81162 28858
rect 81174 28806 81226 28858
rect 81238 28806 81290 28858
rect 111766 28806 111818 28858
rect 111830 28806 111882 28858
rect 111894 28806 111946 28858
rect 111958 28806 112010 28858
rect 142486 28806 142538 28858
rect 142550 28806 142602 28858
rect 142614 28806 142666 28858
rect 142678 28806 142730 28858
rect 173206 28806 173258 28858
rect 173270 28806 173322 28858
rect 173334 28806 173386 28858
rect 173398 28806 173450 28858
rect 4246 28262 4298 28314
rect 4310 28262 4362 28314
rect 4374 28262 4426 28314
rect 4438 28262 4490 28314
rect 34966 28262 35018 28314
rect 35030 28262 35082 28314
rect 35094 28262 35146 28314
rect 35158 28262 35210 28314
rect 65686 28262 65738 28314
rect 65750 28262 65802 28314
rect 65814 28262 65866 28314
rect 65878 28262 65930 28314
rect 96406 28262 96458 28314
rect 96470 28262 96522 28314
rect 96534 28262 96586 28314
rect 96598 28262 96650 28314
rect 127126 28262 127178 28314
rect 127190 28262 127242 28314
rect 127254 28262 127306 28314
rect 127318 28262 127370 28314
rect 157846 28262 157898 28314
rect 157910 28262 157962 28314
rect 157974 28262 158026 28314
rect 158038 28262 158090 28314
rect 19606 27718 19658 27770
rect 19670 27718 19722 27770
rect 19734 27718 19786 27770
rect 19798 27718 19850 27770
rect 50326 27718 50378 27770
rect 50390 27718 50442 27770
rect 50454 27718 50506 27770
rect 50518 27718 50570 27770
rect 81046 27718 81098 27770
rect 81110 27718 81162 27770
rect 81174 27718 81226 27770
rect 81238 27718 81290 27770
rect 111766 27718 111818 27770
rect 111830 27718 111882 27770
rect 111894 27718 111946 27770
rect 111958 27718 112010 27770
rect 142486 27718 142538 27770
rect 142550 27718 142602 27770
rect 142614 27718 142666 27770
rect 142678 27718 142730 27770
rect 173206 27718 173258 27770
rect 173270 27718 173322 27770
rect 173334 27718 173386 27770
rect 173398 27718 173450 27770
rect 4246 27174 4298 27226
rect 4310 27174 4362 27226
rect 4374 27174 4426 27226
rect 4438 27174 4490 27226
rect 34966 27174 35018 27226
rect 35030 27174 35082 27226
rect 35094 27174 35146 27226
rect 35158 27174 35210 27226
rect 65686 27174 65738 27226
rect 65750 27174 65802 27226
rect 65814 27174 65866 27226
rect 65878 27174 65930 27226
rect 96406 27174 96458 27226
rect 96470 27174 96522 27226
rect 96534 27174 96586 27226
rect 96598 27174 96650 27226
rect 127126 27174 127178 27226
rect 127190 27174 127242 27226
rect 127254 27174 127306 27226
rect 127318 27174 127370 27226
rect 157846 27174 157898 27226
rect 157910 27174 157962 27226
rect 157974 27174 158026 27226
rect 158038 27174 158090 27226
rect 19606 26630 19658 26682
rect 19670 26630 19722 26682
rect 19734 26630 19786 26682
rect 19798 26630 19850 26682
rect 50326 26630 50378 26682
rect 50390 26630 50442 26682
rect 50454 26630 50506 26682
rect 50518 26630 50570 26682
rect 81046 26630 81098 26682
rect 81110 26630 81162 26682
rect 81174 26630 81226 26682
rect 81238 26630 81290 26682
rect 111766 26630 111818 26682
rect 111830 26630 111882 26682
rect 111894 26630 111946 26682
rect 111958 26630 112010 26682
rect 142486 26630 142538 26682
rect 142550 26630 142602 26682
rect 142614 26630 142666 26682
rect 142678 26630 142730 26682
rect 173206 26630 173258 26682
rect 173270 26630 173322 26682
rect 173334 26630 173386 26682
rect 173398 26630 173450 26682
rect 4246 26086 4298 26138
rect 4310 26086 4362 26138
rect 4374 26086 4426 26138
rect 4438 26086 4490 26138
rect 34966 26086 35018 26138
rect 35030 26086 35082 26138
rect 35094 26086 35146 26138
rect 35158 26086 35210 26138
rect 65686 26086 65738 26138
rect 65750 26086 65802 26138
rect 65814 26086 65866 26138
rect 65878 26086 65930 26138
rect 96406 26086 96458 26138
rect 96470 26086 96522 26138
rect 96534 26086 96586 26138
rect 96598 26086 96650 26138
rect 127126 26086 127178 26138
rect 127190 26086 127242 26138
rect 127254 26086 127306 26138
rect 127318 26086 127370 26138
rect 157846 26086 157898 26138
rect 157910 26086 157962 26138
rect 157974 26086 158026 26138
rect 158038 26086 158090 26138
rect 19606 25542 19658 25594
rect 19670 25542 19722 25594
rect 19734 25542 19786 25594
rect 19798 25542 19850 25594
rect 50326 25542 50378 25594
rect 50390 25542 50442 25594
rect 50454 25542 50506 25594
rect 50518 25542 50570 25594
rect 81046 25542 81098 25594
rect 81110 25542 81162 25594
rect 81174 25542 81226 25594
rect 81238 25542 81290 25594
rect 111766 25542 111818 25594
rect 111830 25542 111882 25594
rect 111894 25542 111946 25594
rect 111958 25542 112010 25594
rect 142486 25542 142538 25594
rect 142550 25542 142602 25594
rect 142614 25542 142666 25594
rect 142678 25542 142730 25594
rect 173206 25542 173258 25594
rect 173270 25542 173322 25594
rect 173334 25542 173386 25594
rect 173398 25542 173450 25594
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 34966 24998 35018 25050
rect 35030 24998 35082 25050
rect 35094 24998 35146 25050
rect 35158 24998 35210 25050
rect 65686 24998 65738 25050
rect 65750 24998 65802 25050
rect 65814 24998 65866 25050
rect 65878 24998 65930 25050
rect 96406 24998 96458 25050
rect 96470 24998 96522 25050
rect 96534 24998 96586 25050
rect 96598 24998 96650 25050
rect 127126 24998 127178 25050
rect 127190 24998 127242 25050
rect 127254 24998 127306 25050
rect 127318 24998 127370 25050
rect 157846 24998 157898 25050
rect 157910 24998 157962 25050
rect 157974 24998 158026 25050
rect 158038 24998 158090 25050
rect 19606 24454 19658 24506
rect 19670 24454 19722 24506
rect 19734 24454 19786 24506
rect 19798 24454 19850 24506
rect 50326 24454 50378 24506
rect 50390 24454 50442 24506
rect 50454 24454 50506 24506
rect 50518 24454 50570 24506
rect 81046 24454 81098 24506
rect 81110 24454 81162 24506
rect 81174 24454 81226 24506
rect 81238 24454 81290 24506
rect 111766 24454 111818 24506
rect 111830 24454 111882 24506
rect 111894 24454 111946 24506
rect 111958 24454 112010 24506
rect 142486 24454 142538 24506
rect 142550 24454 142602 24506
rect 142614 24454 142666 24506
rect 142678 24454 142730 24506
rect 173206 24454 173258 24506
rect 173270 24454 173322 24506
rect 173334 24454 173386 24506
rect 173398 24454 173450 24506
rect 31024 24216 31076 24268
rect 31392 24216 31444 24268
rect 35900 24216 35952 24268
rect 36820 24216 36872 24268
rect 33140 24012 33192 24064
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 34966 23910 35018 23962
rect 35030 23910 35082 23962
rect 35094 23910 35146 23962
rect 35158 23910 35210 23962
rect 65686 23910 65738 23962
rect 65750 23910 65802 23962
rect 65814 23910 65866 23962
rect 65878 23910 65930 23962
rect 96406 23910 96458 23962
rect 96470 23910 96522 23962
rect 96534 23910 96586 23962
rect 96598 23910 96650 23962
rect 127126 23910 127178 23962
rect 127190 23910 127242 23962
rect 127254 23910 127306 23962
rect 127318 23910 127370 23962
rect 157846 23910 157898 23962
rect 157910 23910 157962 23962
rect 157974 23910 158026 23962
rect 158038 23910 158090 23962
rect 19606 23366 19658 23418
rect 19670 23366 19722 23418
rect 19734 23366 19786 23418
rect 19798 23366 19850 23418
rect 50326 23366 50378 23418
rect 50390 23366 50442 23418
rect 50454 23366 50506 23418
rect 50518 23366 50570 23418
rect 81046 23366 81098 23418
rect 81110 23366 81162 23418
rect 81174 23366 81226 23418
rect 81238 23366 81290 23418
rect 111766 23366 111818 23418
rect 111830 23366 111882 23418
rect 111894 23366 111946 23418
rect 111958 23366 112010 23418
rect 142486 23366 142538 23418
rect 142550 23366 142602 23418
rect 142614 23366 142666 23418
rect 142678 23366 142730 23418
rect 173206 23366 173258 23418
rect 173270 23366 173322 23418
rect 173334 23366 173386 23418
rect 173398 23366 173450 23418
rect 26424 23171 26476 23180
rect 26424 23137 26433 23171
rect 26433 23137 26467 23171
rect 26467 23137 26476 23171
rect 26424 23128 26476 23137
rect 26608 23171 26660 23180
rect 26608 23137 26617 23171
rect 26617 23137 26651 23171
rect 26651 23137 26660 23171
rect 26608 23128 26660 23137
rect 28264 23128 28316 23180
rect 28172 23060 28224 23112
rect 27988 22924 28040 22976
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 34966 22822 35018 22874
rect 35030 22822 35082 22874
rect 35094 22822 35146 22874
rect 35158 22822 35210 22874
rect 65686 22822 65738 22874
rect 65750 22822 65802 22874
rect 65814 22822 65866 22874
rect 65878 22822 65930 22874
rect 96406 22822 96458 22874
rect 96470 22822 96522 22874
rect 96534 22822 96586 22874
rect 96598 22822 96650 22874
rect 127126 22822 127178 22874
rect 127190 22822 127242 22874
rect 127254 22822 127306 22874
rect 127318 22822 127370 22874
rect 157846 22822 157898 22874
rect 157910 22822 157962 22874
rect 157974 22822 158026 22874
rect 158038 22822 158090 22874
rect 33140 22627 33192 22636
rect 33140 22593 33149 22627
rect 33149 22593 33183 22627
rect 33183 22593 33192 22627
rect 33140 22584 33192 22593
rect 32128 22516 32180 22568
rect 30380 22448 30432 22500
rect 33416 22423 33468 22432
rect 33416 22389 33425 22423
rect 33425 22389 33459 22423
rect 33459 22389 33468 22423
rect 33416 22380 33468 22389
rect 35256 22380 35308 22432
rect 19606 22278 19658 22330
rect 19670 22278 19722 22330
rect 19734 22278 19786 22330
rect 19798 22278 19850 22330
rect 50326 22278 50378 22330
rect 50390 22278 50442 22330
rect 50454 22278 50506 22330
rect 50518 22278 50570 22330
rect 81046 22278 81098 22330
rect 81110 22278 81162 22330
rect 81174 22278 81226 22330
rect 81238 22278 81290 22330
rect 111766 22278 111818 22330
rect 111830 22278 111882 22330
rect 111894 22278 111946 22330
rect 111958 22278 112010 22330
rect 142486 22278 142538 22330
rect 142550 22278 142602 22330
rect 142614 22278 142666 22330
rect 142678 22278 142730 22330
rect 173206 22278 173258 22330
rect 173270 22278 173322 22330
rect 173334 22278 173386 22330
rect 173398 22278 173450 22330
rect 29092 22151 29144 22160
rect 29092 22117 29101 22151
rect 29101 22117 29135 22151
rect 29135 22117 29144 22151
rect 29092 22108 29144 22117
rect 29276 22151 29328 22160
rect 29276 22117 29306 22151
rect 29306 22117 29328 22151
rect 29276 22108 29328 22117
rect 30380 21904 30432 21956
rect 29184 21836 29236 21888
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 34966 21734 35018 21786
rect 35030 21734 35082 21786
rect 35094 21734 35146 21786
rect 35158 21734 35210 21786
rect 65686 21734 65738 21786
rect 65750 21734 65802 21786
rect 65814 21734 65866 21786
rect 65878 21734 65930 21786
rect 96406 21734 96458 21786
rect 96470 21734 96522 21786
rect 96534 21734 96586 21786
rect 96598 21734 96650 21786
rect 127126 21734 127178 21786
rect 127190 21734 127242 21786
rect 127254 21734 127306 21786
rect 127318 21734 127370 21786
rect 157846 21734 157898 21786
rect 157910 21734 157962 21786
rect 157974 21734 158026 21786
rect 158038 21734 158090 21786
rect 27988 21471 28040 21480
rect 27988 21437 27997 21471
rect 27997 21437 28031 21471
rect 28031 21437 28040 21471
rect 27988 21428 28040 21437
rect 29276 21292 29328 21344
rect 19606 21190 19658 21242
rect 19670 21190 19722 21242
rect 19734 21190 19786 21242
rect 19798 21190 19850 21242
rect 50326 21190 50378 21242
rect 50390 21190 50442 21242
rect 50454 21190 50506 21242
rect 50518 21190 50570 21242
rect 81046 21190 81098 21242
rect 81110 21190 81162 21242
rect 81174 21190 81226 21242
rect 81238 21190 81290 21242
rect 111766 21190 111818 21242
rect 111830 21190 111882 21242
rect 111894 21190 111946 21242
rect 111958 21190 112010 21242
rect 142486 21190 142538 21242
rect 142550 21190 142602 21242
rect 142614 21190 142666 21242
rect 142678 21190 142730 21242
rect 173206 21190 173258 21242
rect 173270 21190 173322 21242
rect 173334 21190 173386 21242
rect 173398 21190 173450 21242
rect 29092 21020 29144 21072
rect 32036 21020 32088 21072
rect 29184 20995 29236 21004
rect 29184 20961 29193 20995
rect 29193 20961 29227 20995
rect 29227 20961 29236 20995
rect 29184 20952 29236 20961
rect 29276 20995 29328 21004
rect 29276 20961 29285 20995
rect 29285 20961 29319 20995
rect 29319 20961 29328 20995
rect 29276 20952 29328 20961
rect 30656 20748 30708 20800
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 34966 20646 35018 20698
rect 35030 20646 35082 20698
rect 35094 20646 35146 20698
rect 35158 20646 35210 20698
rect 65686 20646 65738 20698
rect 65750 20646 65802 20698
rect 65814 20646 65866 20698
rect 65878 20646 65930 20698
rect 96406 20646 96458 20698
rect 96470 20646 96522 20698
rect 96534 20646 96586 20698
rect 96598 20646 96650 20698
rect 127126 20646 127178 20698
rect 127190 20646 127242 20698
rect 127254 20646 127306 20698
rect 127318 20646 127370 20698
rect 157846 20646 157898 20698
rect 157910 20646 157962 20698
rect 157974 20646 158026 20698
rect 158038 20646 158090 20698
rect 28172 20451 28224 20460
rect 28172 20417 28181 20451
rect 28181 20417 28215 20451
rect 28215 20417 28224 20451
rect 28172 20408 28224 20417
rect 33232 20408 33284 20460
rect 27988 20383 28040 20392
rect 27988 20349 27997 20383
rect 27997 20349 28031 20383
rect 28031 20349 28040 20383
rect 27988 20340 28040 20349
rect 28264 20383 28316 20392
rect 28264 20349 28273 20383
rect 28273 20349 28307 20383
rect 28307 20349 28316 20383
rect 28264 20340 28316 20349
rect 29092 20340 29144 20392
rect 29000 20204 29052 20256
rect 74540 20204 74592 20256
rect 149520 20340 149572 20392
rect 75828 20204 75880 20256
rect 19606 20102 19658 20154
rect 19670 20102 19722 20154
rect 19734 20102 19786 20154
rect 19798 20102 19850 20154
rect 50326 20102 50378 20154
rect 50390 20102 50442 20154
rect 50454 20102 50506 20154
rect 50518 20102 50570 20154
rect 81046 20102 81098 20154
rect 81110 20102 81162 20154
rect 81174 20102 81226 20154
rect 81238 20102 81290 20154
rect 111766 20102 111818 20154
rect 111830 20102 111882 20154
rect 111894 20102 111946 20154
rect 111958 20102 112010 20154
rect 142486 20102 142538 20154
rect 142550 20102 142602 20154
rect 142614 20102 142666 20154
rect 142678 20102 142730 20154
rect 173206 20102 173258 20154
rect 173270 20102 173322 20154
rect 173334 20102 173386 20154
rect 173398 20102 173450 20154
rect 29276 20000 29328 20052
rect 29184 19864 29236 19916
rect 72148 20000 72200 20052
rect 121736 20000 121788 20052
rect 73252 19932 73304 19984
rect 130752 19932 130804 19984
rect 30380 19864 30432 19916
rect 31208 19907 31260 19916
rect 31208 19873 31217 19907
rect 31217 19873 31251 19907
rect 31251 19873 31260 19907
rect 31208 19864 31260 19873
rect 31392 19907 31444 19916
rect 31392 19873 31401 19907
rect 31401 19873 31435 19907
rect 31435 19873 31444 19907
rect 31392 19864 31444 19873
rect 31944 19864 31996 19916
rect 31024 19796 31076 19848
rect 28908 19703 28960 19712
rect 28908 19669 28917 19703
rect 28917 19669 28951 19703
rect 28951 19669 28960 19703
rect 28908 19660 28960 19669
rect 31300 19703 31352 19712
rect 31300 19669 31309 19703
rect 31309 19669 31343 19703
rect 31343 19669 31352 19703
rect 31300 19660 31352 19669
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 34966 19558 35018 19610
rect 35030 19558 35082 19610
rect 35094 19558 35146 19610
rect 35158 19558 35210 19610
rect 65686 19558 65738 19610
rect 65750 19558 65802 19610
rect 65814 19558 65866 19610
rect 65878 19558 65930 19610
rect 96406 19558 96458 19610
rect 96470 19558 96522 19610
rect 96534 19558 96586 19610
rect 96598 19558 96650 19610
rect 127126 19558 127178 19610
rect 127190 19558 127242 19610
rect 127254 19558 127306 19610
rect 127318 19558 127370 19610
rect 157846 19558 157898 19610
rect 157910 19558 157962 19610
rect 157974 19558 158026 19610
rect 158038 19558 158090 19610
rect 135444 19456 135496 19508
rect 35256 19252 35308 19304
rect 35808 19252 35860 19304
rect 37740 19252 37792 19304
rect 41696 19252 41748 19304
rect 57152 19295 57204 19304
rect 57152 19261 57161 19295
rect 57161 19261 57195 19295
rect 57195 19261 57204 19295
rect 57152 19252 57204 19261
rect 58072 19252 58124 19304
rect 59268 19295 59320 19304
rect 59268 19261 59277 19295
rect 59277 19261 59311 19295
rect 59311 19261 59320 19295
rect 59268 19252 59320 19261
rect 60188 19295 60240 19304
rect 60188 19261 60197 19295
rect 60197 19261 60231 19295
rect 60231 19261 60240 19295
rect 60188 19252 60240 19261
rect 61016 19295 61068 19304
rect 61016 19261 61025 19295
rect 61025 19261 61059 19295
rect 61059 19261 61068 19295
rect 61016 19252 61068 19261
rect 65248 19295 65300 19304
rect 65248 19261 65257 19295
rect 65257 19261 65291 19295
rect 65291 19261 65300 19295
rect 65248 19252 65300 19261
rect 72884 19252 72936 19304
rect 73252 19252 73304 19304
rect 71320 19184 71372 19236
rect 37464 19116 37516 19168
rect 42800 19116 42852 19168
rect 43444 19116 43496 19168
rect 50896 19116 50948 19168
rect 57244 19159 57296 19168
rect 57244 19125 57253 19159
rect 57253 19125 57287 19159
rect 57287 19125 57296 19159
rect 57244 19116 57296 19125
rect 59360 19159 59412 19168
rect 59360 19125 59369 19159
rect 59369 19125 59403 19159
rect 59403 19125 59412 19159
rect 59360 19116 59412 19125
rect 60188 19116 60240 19168
rect 61108 19159 61160 19168
rect 61108 19125 61117 19159
rect 61117 19125 61151 19159
rect 61151 19125 61160 19159
rect 61108 19116 61160 19125
rect 65984 19116 66036 19168
rect 68652 19116 68704 19168
rect 72884 19116 72936 19168
rect 73160 19116 73212 19168
rect 75276 19184 75328 19236
rect 73528 19116 73580 19168
rect 75000 19159 75052 19168
rect 75000 19125 75009 19159
rect 75009 19125 75043 19159
rect 75043 19125 75052 19159
rect 75000 19116 75052 19125
rect 140412 19116 140464 19168
rect 19606 19014 19658 19066
rect 19670 19014 19722 19066
rect 19734 19014 19786 19066
rect 19798 19014 19850 19066
rect 50326 19014 50378 19066
rect 50390 19014 50442 19066
rect 50454 19014 50506 19066
rect 50518 19014 50570 19066
rect 81046 19014 81098 19066
rect 81110 19014 81162 19066
rect 81174 19014 81226 19066
rect 81238 19014 81290 19066
rect 111766 19014 111818 19066
rect 111830 19014 111882 19066
rect 111894 19014 111946 19066
rect 111958 19014 112010 19066
rect 142486 19014 142538 19066
rect 142550 19014 142602 19066
rect 142614 19014 142666 19066
rect 142678 19014 142730 19066
rect 173206 19014 173258 19066
rect 173270 19014 173322 19066
rect 173334 19014 173386 19066
rect 173398 19014 173450 19066
rect 33416 18776 33468 18828
rect 35348 18776 35400 18828
rect 42800 18776 42852 18828
rect 44640 18912 44692 18964
rect 32128 18640 32180 18692
rect 46940 18844 46992 18896
rect 73252 18844 73304 18896
rect 66076 18819 66128 18828
rect 66076 18785 66085 18819
rect 66085 18785 66119 18819
rect 66119 18785 66128 18819
rect 66076 18776 66128 18785
rect 67824 18819 67876 18828
rect 67824 18785 67833 18819
rect 67833 18785 67867 18819
rect 67867 18785 67876 18819
rect 67824 18776 67876 18785
rect 68468 18819 68520 18828
rect 68468 18785 68477 18819
rect 68477 18785 68511 18819
rect 68511 18785 68520 18819
rect 68468 18776 68520 18785
rect 72240 18776 72292 18828
rect 72424 18819 72476 18828
rect 72424 18785 72433 18819
rect 72433 18785 72467 18819
rect 72467 18785 72476 18819
rect 72424 18776 72476 18785
rect 72976 18776 73028 18828
rect 55588 18708 55640 18760
rect 47860 18640 47912 18692
rect 65524 18640 65576 18692
rect 67088 18640 67140 18692
rect 71136 18640 71188 18692
rect 42892 18572 42944 18624
rect 44088 18615 44140 18624
rect 44088 18581 44097 18615
rect 44097 18581 44131 18615
rect 44131 18581 44140 18615
rect 44088 18572 44140 18581
rect 47032 18615 47084 18624
rect 47032 18581 47041 18615
rect 47041 18581 47075 18615
rect 47075 18581 47084 18615
rect 47032 18572 47084 18581
rect 48320 18572 48372 18624
rect 66168 18615 66220 18624
rect 66168 18581 66177 18615
rect 66177 18581 66211 18615
rect 66211 18581 66220 18615
rect 66168 18572 66220 18581
rect 66904 18572 66956 18624
rect 70860 18572 70912 18624
rect 73896 18615 73948 18624
rect 73896 18581 73905 18615
rect 73905 18581 73939 18615
rect 73939 18581 73948 18615
rect 73896 18572 73948 18581
rect 74356 18887 74408 18896
rect 74356 18853 74391 18887
rect 74391 18853 74408 18887
rect 74356 18844 74408 18853
rect 74264 18819 74316 18828
rect 74264 18785 74273 18819
rect 74273 18785 74307 18819
rect 74307 18785 74316 18819
rect 75000 18819 75052 18828
rect 74264 18776 74316 18785
rect 75000 18785 75009 18819
rect 75009 18785 75043 18819
rect 75043 18785 75052 18819
rect 75000 18776 75052 18785
rect 75092 18751 75144 18760
rect 75092 18717 75101 18751
rect 75101 18717 75135 18751
rect 75135 18717 75144 18751
rect 75092 18708 75144 18717
rect 74264 18640 74316 18692
rect 144552 18776 144604 18828
rect 75828 18572 75880 18624
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 34966 18470 35018 18522
rect 35030 18470 35082 18522
rect 35094 18470 35146 18522
rect 35158 18470 35210 18522
rect 65686 18470 65738 18522
rect 65750 18470 65802 18522
rect 65814 18470 65866 18522
rect 65878 18470 65930 18522
rect 96406 18470 96458 18522
rect 96470 18470 96522 18522
rect 96534 18470 96586 18522
rect 96598 18470 96650 18522
rect 127126 18470 127178 18522
rect 127190 18470 127242 18522
rect 127254 18470 127306 18522
rect 127318 18470 127370 18522
rect 157846 18470 157898 18522
rect 157910 18470 157962 18522
rect 157974 18470 158026 18522
rect 158038 18470 158090 18522
rect 31208 18368 31260 18420
rect 47032 18368 47084 18420
rect 47584 18368 47636 18420
rect 60372 18368 60424 18420
rect 33048 18232 33100 18284
rect 47124 18232 47176 18284
rect 30656 18207 30708 18216
rect 30656 18173 30665 18207
rect 30665 18173 30699 18207
rect 30699 18173 30708 18207
rect 30656 18164 30708 18173
rect 31208 18164 31260 18216
rect 31300 18164 31352 18216
rect 31944 18207 31996 18216
rect 31944 18173 31953 18207
rect 31953 18173 31987 18207
rect 31987 18173 31996 18207
rect 31944 18164 31996 18173
rect 33140 18164 33192 18216
rect 37464 18164 37516 18216
rect 31852 18096 31904 18148
rect 41420 18164 41472 18216
rect 47032 18164 47084 18216
rect 48320 18164 48372 18216
rect 49516 18164 49568 18216
rect 69664 18232 69716 18284
rect 52460 18164 52512 18216
rect 53104 18164 53156 18216
rect 54208 18207 54260 18216
rect 54208 18173 54217 18207
rect 54217 18173 54251 18207
rect 54251 18173 54260 18207
rect 54208 18164 54260 18173
rect 72148 18207 72200 18216
rect 72148 18173 72157 18207
rect 72157 18173 72191 18207
rect 72191 18173 72200 18207
rect 72148 18164 72200 18173
rect 73528 18207 73580 18216
rect 73528 18173 73537 18207
rect 73537 18173 73571 18207
rect 73571 18173 73580 18207
rect 73528 18164 73580 18173
rect 41144 18139 41196 18148
rect 41144 18105 41153 18139
rect 41153 18105 41187 18139
rect 41187 18105 41196 18139
rect 41144 18096 41196 18105
rect 54392 18139 54444 18148
rect 54392 18105 54401 18139
rect 54401 18105 54435 18139
rect 54435 18105 54444 18139
rect 54392 18096 54444 18105
rect 41328 18028 41380 18080
rect 46388 18028 46440 18080
rect 49608 18071 49660 18080
rect 49608 18037 49617 18071
rect 49617 18037 49651 18071
rect 49651 18037 49660 18071
rect 49608 18028 49660 18037
rect 70768 18028 70820 18080
rect 73620 18071 73672 18080
rect 73620 18037 73629 18071
rect 73629 18037 73663 18071
rect 73663 18037 73672 18071
rect 73620 18028 73672 18037
rect 19606 17926 19658 17978
rect 19670 17926 19722 17978
rect 19734 17926 19786 17978
rect 19798 17926 19850 17978
rect 50326 17926 50378 17978
rect 50390 17926 50442 17978
rect 50454 17926 50506 17978
rect 50518 17926 50570 17978
rect 81046 17926 81098 17978
rect 81110 17926 81162 17978
rect 81174 17926 81226 17978
rect 81238 17926 81290 17978
rect 111766 17926 111818 17978
rect 111830 17926 111882 17978
rect 111894 17926 111946 17978
rect 111958 17926 112010 17978
rect 142486 17926 142538 17978
rect 142550 17926 142602 17978
rect 142614 17926 142666 17978
rect 142678 17926 142730 17978
rect 173206 17926 173258 17978
rect 173270 17926 173322 17978
rect 173334 17926 173386 17978
rect 173398 17926 173450 17978
rect 52460 17824 52512 17876
rect 31300 17688 31352 17740
rect 37464 17731 37516 17740
rect 37464 17697 37473 17731
rect 37473 17697 37507 17731
rect 37507 17697 37516 17731
rect 37464 17688 37516 17697
rect 37740 17731 37792 17740
rect 37740 17697 37749 17731
rect 37749 17697 37783 17731
rect 37783 17697 37792 17731
rect 37740 17688 37792 17697
rect 38752 17688 38804 17740
rect 49608 17688 49660 17740
rect 61108 17756 61160 17808
rect 59544 17688 59596 17740
rect 60188 17731 60240 17740
rect 60188 17697 60197 17731
rect 60197 17697 60231 17731
rect 60231 17697 60240 17731
rect 60188 17688 60240 17697
rect 35808 17620 35860 17672
rect 38844 17552 38896 17604
rect 58348 17552 58400 17604
rect 59176 17552 59228 17604
rect 32404 17484 32456 17536
rect 59544 17484 59596 17536
rect 60556 17527 60608 17536
rect 60556 17493 60565 17527
rect 60565 17493 60599 17527
rect 60599 17493 60608 17527
rect 60556 17484 60608 17493
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 34966 17382 35018 17434
rect 35030 17382 35082 17434
rect 35094 17382 35146 17434
rect 35158 17382 35210 17434
rect 65686 17382 65738 17434
rect 65750 17382 65802 17434
rect 65814 17382 65866 17434
rect 65878 17382 65930 17434
rect 96406 17382 96458 17434
rect 96470 17382 96522 17434
rect 96534 17382 96586 17434
rect 96598 17382 96650 17434
rect 127126 17382 127178 17434
rect 127190 17382 127242 17434
rect 127254 17382 127306 17434
rect 127318 17382 127370 17434
rect 157846 17382 157898 17434
rect 157910 17382 157962 17434
rect 157974 17382 158026 17434
rect 158038 17382 158090 17434
rect 46940 17280 46992 17332
rect 48320 17280 48372 17332
rect 60556 17280 60608 17332
rect 70400 17280 70452 17332
rect 70860 17280 70912 17332
rect 72332 17323 72384 17332
rect 72332 17289 72341 17323
rect 72341 17289 72375 17323
rect 72375 17289 72384 17323
rect 72332 17280 72384 17289
rect 73068 17280 73120 17332
rect 43628 17212 43680 17264
rect 57244 17212 57296 17264
rect 63592 17212 63644 17264
rect 65984 17255 66036 17264
rect 65984 17221 65993 17255
rect 65993 17221 66027 17255
rect 66027 17221 66036 17255
rect 65984 17212 66036 17221
rect 35808 17144 35860 17196
rect 35256 17119 35308 17128
rect 35256 17085 35265 17119
rect 35265 17085 35299 17119
rect 35299 17085 35308 17119
rect 35256 17076 35308 17085
rect 35900 17076 35952 17128
rect 43352 17076 43404 17128
rect 44088 17076 44140 17128
rect 46204 17076 46256 17128
rect 49608 17144 49660 17196
rect 49516 17119 49568 17128
rect 49516 17085 49525 17119
rect 49525 17085 49559 17119
rect 49559 17085 49568 17119
rect 49516 17076 49568 17085
rect 59360 17144 59412 17196
rect 58348 17119 58400 17128
rect 56692 17008 56744 17060
rect 56968 17008 57020 17060
rect 58348 17085 58357 17119
rect 58357 17085 58391 17119
rect 58391 17085 58400 17119
rect 58348 17076 58400 17085
rect 63500 17076 63552 17128
rect 66168 17144 66220 17196
rect 66904 17119 66956 17128
rect 66904 17085 66913 17119
rect 66913 17085 66947 17119
rect 66947 17085 66956 17119
rect 66904 17076 66956 17085
rect 67088 17119 67140 17128
rect 67088 17085 67097 17119
rect 67097 17085 67131 17119
rect 67131 17085 67140 17119
rect 67088 17076 67140 17085
rect 69848 17119 69900 17128
rect 69848 17085 69857 17119
rect 69857 17085 69891 17119
rect 69891 17085 69900 17119
rect 69848 17076 69900 17085
rect 70768 17076 70820 17128
rect 71136 17119 71188 17128
rect 71136 17085 71145 17119
rect 71145 17085 71179 17119
rect 71179 17085 71188 17119
rect 71136 17076 71188 17085
rect 71320 17119 71372 17128
rect 71320 17085 71329 17119
rect 71329 17085 71363 17119
rect 71363 17085 71372 17119
rect 71320 17076 71372 17085
rect 71688 17076 71740 17128
rect 75092 17144 75144 17196
rect 73252 17119 73304 17128
rect 73252 17085 73261 17119
rect 73261 17085 73295 17119
rect 73295 17085 73304 17119
rect 73252 17076 73304 17085
rect 36360 16940 36412 16992
rect 49056 16983 49108 16992
rect 49056 16949 49065 16983
rect 49065 16949 49099 16983
rect 49099 16949 49108 16983
rect 49056 16940 49108 16949
rect 59728 16940 59780 16992
rect 69940 17008 69992 17060
rect 74264 17076 74316 17128
rect 66168 16940 66220 16992
rect 66352 16983 66404 16992
rect 66352 16949 66361 16983
rect 66361 16949 66395 16983
rect 66395 16949 66404 16983
rect 66352 16940 66404 16949
rect 70216 16983 70268 16992
rect 70216 16949 70225 16983
rect 70225 16949 70259 16983
rect 70259 16949 70268 16983
rect 70216 16940 70268 16949
rect 71504 16983 71556 16992
rect 71504 16949 71513 16983
rect 71513 16949 71547 16983
rect 71547 16949 71556 16983
rect 71504 16940 71556 16949
rect 72516 16940 72568 16992
rect 19606 16838 19658 16890
rect 19670 16838 19722 16890
rect 19734 16838 19786 16890
rect 19798 16838 19850 16890
rect 50326 16838 50378 16890
rect 50390 16838 50442 16890
rect 50454 16838 50506 16890
rect 50518 16838 50570 16890
rect 81046 16838 81098 16890
rect 81110 16838 81162 16890
rect 81174 16838 81226 16890
rect 81238 16838 81290 16890
rect 111766 16838 111818 16890
rect 111830 16838 111882 16890
rect 111894 16838 111946 16890
rect 111958 16838 112010 16890
rect 142486 16838 142538 16890
rect 142550 16838 142602 16890
rect 142614 16838 142666 16890
rect 142678 16838 142730 16890
rect 173206 16838 173258 16890
rect 173270 16838 173322 16890
rect 173334 16838 173386 16890
rect 173398 16838 173450 16890
rect 32128 16736 32180 16788
rect 33692 16736 33744 16788
rect 42892 16779 42944 16788
rect 42892 16745 42901 16779
rect 42901 16745 42935 16779
rect 42935 16745 42944 16779
rect 42892 16736 42944 16745
rect 43628 16736 43680 16788
rect 43812 16711 43864 16720
rect 32220 16600 32272 16652
rect 32404 16643 32456 16652
rect 32404 16609 32413 16643
rect 32413 16609 32447 16643
rect 32447 16609 32456 16643
rect 32404 16600 32456 16609
rect 40960 16643 41012 16652
rect 40960 16609 40969 16643
rect 40969 16609 41003 16643
rect 41003 16609 41012 16643
rect 40960 16600 41012 16609
rect 41144 16643 41196 16652
rect 41144 16609 41153 16643
rect 41153 16609 41187 16643
rect 41187 16609 41196 16643
rect 43812 16677 43821 16711
rect 43821 16677 43855 16711
rect 43855 16677 43864 16711
rect 43812 16668 43864 16677
rect 41144 16600 41196 16609
rect 41328 16575 41380 16584
rect 41328 16541 41337 16575
rect 41337 16541 41371 16575
rect 41371 16541 41380 16575
rect 41328 16532 41380 16541
rect 41420 16575 41472 16584
rect 41420 16541 41429 16575
rect 41429 16541 41463 16575
rect 41463 16541 41472 16575
rect 43352 16600 43404 16652
rect 43628 16643 43680 16652
rect 43628 16609 43637 16643
rect 43637 16609 43671 16643
rect 43671 16609 43680 16643
rect 43628 16600 43680 16609
rect 46204 16643 46256 16652
rect 46204 16609 46213 16643
rect 46213 16609 46247 16643
rect 46247 16609 46256 16643
rect 46204 16600 46256 16609
rect 46388 16643 46440 16652
rect 46388 16609 46397 16643
rect 46397 16609 46431 16643
rect 46431 16609 46440 16643
rect 46388 16600 46440 16609
rect 47216 16643 47268 16652
rect 47216 16609 47225 16643
rect 47225 16609 47259 16643
rect 47259 16609 47268 16643
rect 47216 16600 47268 16609
rect 48320 16668 48372 16720
rect 47860 16643 47912 16652
rect 41420 16532 41472 16541
rect 46940 16532 46992 16584
rect 47860 16609 47869 16643
rect 47869 16609 47903 16643
rect 47903 16609 47912 16643
rect 47860 16600 47912 16609
rect 52736 16643 52788 16652
rect 52736 16609 52745 16643
rect 52745 16609 52779 16643
rect 52779 16609 52788 16643
rect 52736 16600 52788 16609
rect 54392 16668 54444 16720
rect 60096 16736 60148 16788
rect 53196 16643 53248 16652
rect 53196 16609 53205 16643
rect 53205 16609 53239 16643
rect 53239 16609 53248 16643
rect 53196 16600 53248 16609
rect 54208 16600 54260 16652
rect 56692 16643 56744 16652
rect 56692 16609 56701 16643
rect 56701 16609 56735 16643
rect 56735 16609 56744 16643
rect 56692 16600 56744 16609
rect 56876 16643 56928 16652
rect 56876 16609 56885 16643
rect 56885 16609 56919 16643
rect 56919 16609 56928 16643
rect 56876 16600 56928 16609
rect 57244 16600 57296 16652
rect 58256 16600 58308 16652
rect 58716 16643 58768 16652
rect 58716 16609 58725 16643
rect 58725 16609 58759 16643
rect 58759 16609 58768 16643
rect 58716 16600 58768 16609
rect 66352 16668 66404 16720
rect 59452 16600 59504 16652
rect 53104 16575 53156 16584
rect 53104 16541 53113 16575
rect 53113 16541 53147 16575
rect 53147 16541 53156 16575
rect 53104 16532 53156 16541
rect 59176 16532 59228 16584
rect 65524 16600 65576 16652
rect 67088 16600 67140 16652
rect 69848 16668 69900 16720
rect 66260 16575 66312 16584
rect 66260 16541 66269 16575
rect 66269 16541 66303 16575
rect 66303 16541 66312 16575
rect 66260 16532 66312 16541
rect 66904 16532 66956 16584
rect 71504 16600 71556 16652
rect 72424 16643 72476 16652
rect 72424 16609 72433 16643
rect 72433 16609 72467 16643
rect 72467 16609 72476 16643
rect 72424 16600 72476 16609
rect 73252 16668 73304 16720
rect 72884 16643 72936 16652
rect 72884 16609 72893 16643
rect 72893 16609 72927 16643
rect 72927 16609 72936 16643
rect 72884 16600 72936 16609
rect 73068 16643 73120 16652
rect 73068 16609 73077 16643
rect 73077 16609 73111 16643
rect 73111 16609 73120 16643
rect 73068 16600 73120 16609
rect 75276 16600 75328 16652
rect 70400 16532 70452 16584
rect 70768 16575 70820 16584
rect 70768 16541 70777 16575
rect 70777 16541 70811 16575
rect 70811 16541 70820 16575
rect 70768 16532 70820 16541
rect 71688 16532 71740 16584
rect 42800 16396 42852 16448
rect 56692 16439 56744 16448
rect 56692 16405 56701 16439
rect 56701 16405 56735 16439
rect 56735 16405 56744 16439
rect 56692 16396 56744 16405
rect 58992 16439 59044 16448
rect 58992 16405 59001 16439
rect 59001 16405 59035 16439
rect 59035 16405 59044 16439
rect 58992 16396 59044 16405
rect 66168 16439 66220 16448
rect 66168 16405 66177 16439
rect 66177 16405 66211 16439
rect 66211 16405 66220 16439
rect 66168 16396 66220 16405
rect 68928 16439 68980 16448
rect 68928 16405 68937 16439
rect 68937 16405 68971 16439
rect 68971 16405 68980 16439
rect 68928 16396 68980 16405
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 34966 16294 35018 16346
rect 35030 16294 35082 16346
rect 35094 16294 35146 16346
rect 35158 16294 35210 16346
rect 65686 16294 65738 16346
rect 65750 16294 65802 16346
rect 65814 16294 65866 16346
rect 65878 16294 65930 16346
rect 96406 16294 96458 16346
rect 96470 16294 96522 16346
rect 96534 16294 96586 16346
rect 96598 16294 96650 16346
rect 127126 16294 127178 16346
rect 127190 16294 127242 16346
rect 127254 16294 127306 16346
rect 127318 16294 127370 16346
rect 157846 16294 157898 16346
rect 157910 16294 157962 16346
rect 157974 16294 158026 16346
rect 158038 16294 158090 16346
rect 32404 16192 32456 16244
rect 31944 16124 31996 16176
rect 34520 16192 34572 16244
rect 35256 16192 35308 16244
rect 69020 16192 69072 16244
rect 71872 16235 71924 16244
rect 71872 16201 71881 16235
rect 71881 16201 71915 16235
rect 71915 16201 71924 16235
rect 71872 16192 71924 16201
rect 72884 16192 72936 16244
rect 44732 16124 44784 16176
rect 45836 16167 45888 16176
rect 45836 16133 45845 16167
rect 45845 16133 45879 16167
rect 45879 16133 45888 16167
rect 45836 16124 45888 16133
rect 32128 16031 32180 16040
rect 32128 15997 32137 16031
rect 32137 15997 32171 16031
rect 32171 15997 32180 16031
rect 32128 15988 32180 15997
rect 43812 15988 43864 16040
rect 46940 16056 46992 16108
rect 56692 16056 56744 16108
rect 67824 16124 67876 16176
rect 65708 16099 65760 16108
rect 46204 15988 46256 16040
rect 32220 15920 32272 15972
rect 36084 15920 36136 15972
rect 32404 15852 32456 15904
rect 44180 15920 44232 15972
rect 46388 15920 46440 15972
rect 58072 15988 58124 16040
rect 63500 15988 63552 16040
rect 63592 16031 63644 16040
rect 63592 15997 63601 16031
rect 63601 15997 63635 16031
rect 63635 15997 63644 16031
rect 63592 15988 63644 15997
rect 65340 15988 65392 16040
rect 65708 16065 65717 16099
rect 65717 16065 65751 16099
rect 65751 16065 65760 16099
rect 65708 16056 65760 16065
rect 66168 16056 66220 16108
rect 58992 15920 59044 15972
rect 66076 15988 66128 16040
rect 71136 16056 71188 16108
rect 70216 15988 70268 16040
rect 70492 16031 70544 16040
rect 70492 15997 70501 16031
rect 70501 15997 70535 16031
rect 70535 15997 70544 16031
rect 70492 15988 70544 15997
rect 47032 15852 47084 15904
rect 57060 15895 57112 15904
rect 57060 15861 57069 15895
rect 57069 15861 57103 15895
rect 57103 15861 57112 15895
rect 57060 15852 57112 15861
rect 64052 15852 64104 15904
rect 65248 15895 65300 15904
rect 65248 15861 65257 15895
rect 65257 15861 65291 15895
rect 65291 15861 65300 15895
rect 65248 15852 65300 15861
rect 69848 15852 69900 15904
rect 71688 15988 71740 16040
rect 72056 16031 72108 16040
rect 72056 15997 72065 16031
rect 72065 15997 72099 16031
rect 72099 15997 72108 16031
rect 72056 15988 72108 15997
rect 73620 15988 73672 16040
rect 71320 15963 71372 15972
rect 71320 15929 71329 15963
rect 71329 15929 71363 15963
rect 71363 15929 71372 15963
rect 71320 15920 71372 15929
rect 72332 15852 72384 15904
rect 19606 15750 19658 15802
rect 19670 15750 19722 15802
rect 19734 15750 19786 15802
rect 19798 15750 19850 15802
rect 50326 15750 50378 15802
rect 50390 15750 50442 15802
rect 50454 15750 50506 15802
rect 50518 15750 50570 15802
rect 81046 15750 81098 15802
rect 81110 15750 81162 15802
rect 81174 15750 81226 15802
rect 81238 15750 81290 15802
rect 111766 15750 111818 15802
rect 111830 15750 111882 15802
rect 111894 15750 111946 15802
rect 111958 15750 112010 15802
rect 142486 15750 142538 15802
rect 142550 15750 142602 15802
rect 142614 15750 142666 15802
rect 142678 15750 142730 15802
rect 173206 15750 173258 15802
rect 173270 15750 173322 15802
rect 173334 15750 173386 15802
rect 173398 15750 173450 15802
rect 29000 15648 29052 15700
rect 31852 15648 31904 15700
rect 56876 15691 56928 15700
rect 56876 15657 56885 15691
rect 56885 15657 56919 15691
rect 56919 15657 56928 15691
rect 56876 15648 56928 15657
rect 63592 15648 63644 15700
rect 70492 15648 70544 15700
rect 72056 15648 72108 15700
rect 29092 15512 29144 15564
rect 30012 15512 30064 15564
rect 32036 15580 32088 15632
rect 56692 15623 56744 15632
rect 56692 15589 56701 15623
rect 56701 15589 56735 15623
rect 56735 15589 56744 15623
rect 56692 15580 56744 15589
rect 33692 15555 33744 15564
rect 33692 15521 33701 15555
rect 33701 15521 33735 15555
rect 33735 15521 33744 15555
rect 33692 15512 33744 15521
rect 34520 15512 34572 15564
rect 56968 15555 57020 15564
rect 56968 15521 56977 15555
rect 56977 15521 57011 15555
rect 57011 15521 57020 15555
rect 56968 15512 57020 15521
rect 59728 15512 59780 15564
rect 31208 15444 31260 15496
rect 63500 15512 63552 15564
rect 64052 15555 64104 15564
rect 64052 15521 64061 15555
rect 64061 15521 64095 15555
rect 64095 15521 64104 15555
rect 64052 15512 64104 15521
rect 63960 15444 64012 15496
rect 65984 15512 66036 15564
rect 71872 15580 71924 15632
rect 69848 15555 69900 15564
rect 69848 15521 69857 15555
rect 69857 15521 69891 15555
rect 69891 15521 69900 15555
rect 69848 15512 69900 15521
rect 70216 15512 70268 15564
rect 71688 15512 71740 15564
rect 68928 15444 68980 15496
rect 69388 15487 69440 15496
rect 69388 15453 69397 15487
rect 69397 15453 69431 15487
rect 69431 15453 69440 15487
rect 69388 15444 69440 15453
rect 72148 15444 72200 15496
rect 65708 15376 65760 15428
rect 28816 15351 28868 15360
rect 28816 15317 28825 15351
rect 28825 15317 28859 15351
rect 28859 15317 28868 15351
rect 28816 15308 28868 15317
rect 31484 15351 31536 15360
rect 31484 15317 31493 15351
rect 31493 15317 31527 15351
rect 31527 15317 31536 15351
rect 31484 15308 31536 15317
rect 34796 15308 34848 15360
rect 55312 15308 55364 15360
rect 62488 15351 62540 15360
rect 62488 15317 62497 15351
rect 62497 15317 62531 15351
rect 62531 15317 62540 15351
rect 62488 15308 62540 15317
rect 63684 15351 63736 15360
rect 63684 15317 63693 15351
rect 63693 15317 63727 15351
rect 63727 15317 63736 15351
rect 63684 15308 63736 15317
rect 67640 15308 67692 15360
rect 70032 15351 70084 15360
rect 70032 15317 70041 15351
rect 70041 15317 70075 15351
rect 70075 15317 70084 15351
rect 70032 15308 70084 15317
rect 70124 15308 70176 15360
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 34966 15206 35018 15258
rect 35030 15206 35082 15258
rect 35094 15206 35146 15258
rect 35158 15206 35210 15258
rect 65686 15206 65738 15258
rect 65750 15206 65802 15258
rect 65814 15206 65866 15258
rect 65878 15206 65930 15258
rect 96406 15206 96458 15258
rect 96470 15206 96522 15258
rect 96534 15206 96586 15258
rect 96598 15206 96650 15258
rect 127126 15206 127178 15258
rect 127190 15206 127242 15258
rect 127254 15206 127306 15258
rect 127318 15206 127370 15258
rect 157846 15206 157898 15258
rect 157910 15206 157962 15258
rect 157974 15206 158026 15258
rect 158038 15206 158090 15258
rect 32496 15036 32548 15088
rect 28908 14968 28960 15020
rect 31208 15011 31260 15020
rect 31208 14977 31217 15011
rect 31217 14977 31251 15011
rect 31251 14977 31260 15011
rect 31208 14968 31260 14977
rect 63500 14968 63552 15020
rect 33508 14943 33560 14952
rect 33508 14909 33517 14943
rect 33517 14909 33551 14943
rect 33551 14909 33560 14943
rect 33508 14900 33560 14909
rect 33784 14943 33836 14952
rect 33784 14909 33793 14943
rect 33793 14909 33827 14943
rect 33827 14909 33836 14943
rect 33784 14900 33836 14909
rect 59544 14900 59596 14952
rect 65524 14900 65576 14952
rect 35348 14832 35400 14884
rect 59728 14875 59780 14884
rect 59728 14841 59737 14875
rect 59737 14841 59771 14875
rect 59771 14841 59780 14875
rect 59728 14832 59780 14841
rect 60096 14875 60148 14884
rect 60096 14841 60105 14875
rect 60105 14841 60139 14875
rect 60139 14841 60148 14875
rect 60096 14832 60148 14841
rect 66352 14832 66404 14884
rect 68560 14900 68612 14952
rect 68928 14832 68980 14884
rect 73528 14832 73580 14884
rect 31024 14807 31076 14816
rect 31024 14773 31033 14807
rect 31033 14773 31067 14807
rect 31067 14773 31076 14807
rect 31024 14764 31076 14773
rect 32220 14764 32272 14816
rect 65524 14764 65576 14816
rect 70400 14764 70452 14816
rect 19606 14662 19658 14714
rect 19670 14662 19722 14714
rect 19734 14662 19786 14714
rect 19798 14662 19850 14714
rect 50326 14662 50378 14714
rect 50390 14662 50442 14714
rect 50454 14662 50506 14714
rect 50518 14662 50570 14714
rect 81046 14662 81098 14714
rect 81110 14662 81162 14714
rect 81174 14662 81226 14714
rect 81238 14662 81290 14714
rect 111766 14662 111818 14714
rect 111830 14662 111882 14714
rect 111894 14662 111946 14714
rect 111958 14662 112010 14714
rect 142486 14662 142538 14714
rect 142550 14662 142602 14714
rect 142614 14662 142666 14714
rect 142678 14662 142730 14714
rect 173206 14662 173258 14714
rect 173270 14662 173322 14714
rect 173334 14662 173386 14714
rect 173398 14662 173450 14714
rect 33048 14560 33100 14612
rect 70124 14560 70176 14612
rect 31760 14492 31812 14544
rect 31116 14467 31168 14476
rect 31116 14433 31125 14467
rect 31125 14433 31159 14467
rect 31159 14433 31168 14467
rect 39672 14492 39724 14544
rect 31116 14424 31168 14433
rect 33140 14467 33192 14476
rect 33140 14433 33149 14467
rect 33149 14433 33183 14467
rect 33183 14433 33192 14467
rect 33140 14424 33192 14433
rect 34612 14424 34664 14476
rect 73896 14492 73948 14544
rect 68560 14467 68612 14476
rect 31208 14356 31260 14408
rect 33968 14356 34020 14408
rect 68560 14433 68569 14467
rect 68569 14433 68603 14467
rect 68603 14433 68612 14467
rect 68560 14424 68612 14433
rect 69756 14467 69808 14476
rect 69756 14433 69765 14467
rect 69765 14433 69799 14467
rect 69799 14433 69808 14467
rect 69756 14424 69808 14433
rect 74356 14424 74408 14476
rect 69112 14356 69164 14408
rect 70308 14356 70360 14408
rect 34244 14331 34296 14340
rect 34244 14297 34253 14331
rect 34253 14297 34287 14331
rect 34287 14297 34296 14331
rect 34244 14288 34296 14297
rect 55220 14288 55272 14340
rect 101312 14288 101364 14340
rect 33140 14220 33192 14272
rect 46940 14263 46992 14272
rect 46940 14229 46949 14263
rect 46949 14229 46983 14263
rect 46983 14229 46992 14263
rect 46940 14220 46992 14229
rect 68192 14263 68244 14272
rect 68192 14229 68201 14263
rect 68201 14229 68235 14263
rect 68235 14229 68244 14263
rect 68192 14220 68244 14229
rect 68284 14220 68336 14272
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 34966 14118 35018 14170
rect 35030 14118 35082 14170
rect 35094 14118 35146 14170
rect 35158 14118 35210 14170
rect 65686 14118 65738 14170
rect 65750 14118 65802 14170
rect 65814 14118 65866 14170
rect 65878 14118 65930 14170
rect 96406 14118 96458 14170
rect 96470 14118 96522 14170
rect 96534 14118 96586 14170
rect 96598 14118 96650 14170
rect 127126 14118 127178 14170
rect 127190 14118 127242 14170
rect 127254 14118 127306 14170
rect 127318 14118 127370 14170
rect 157846 14118 157898 14170
rect 157910 14118 157962 14170
rect 157974 14118 158026 14170
rect 158038 14118 158090 14170
rect 30012 14016 30064 14068
rect 41144 14016 41196 14068
rect 48044 14016 48096 14068
rect 57244 14016 57296 14068
rect 62396 14016 62448 14068
rect 35256 13948 35308 14000
rect 36636 13948 36688 14000
rect 39580 13948 39632 14000
rect 30840 13880 30892 13932
rect 31944 13880 31996 13932
rect 36360 13923 36412 13932
rect 31668 13812 31720 13864
rect 33968 13812 34020 13864
rect 36360 13889 36369 13923
rect 36369 13889 36403 13923
rect 36403 13889 36412 13923
rect 36360 13880 36412 13889
rect 38844 13923 38896 13932
rect 38844 13889 38853 13923
rect 38853 13889 38887 13923
rect 38887 13889 38896 13923
rect 38844 13880 38896 13889
rect 40960 13880 41012 13932
rect 47860 13948 47912 14000
rect 56600 13948 56652 14000
rect 43628 13880 43680 13932
rect 47216 13880 47268 13932
rect 39672 13855 39724 13864
rect 35900 13744 35952 13796
rect 36544 13744 36596 13796
rect 39672 13821 39681 13855
rect 39681 13821 39715 13855
rect 39715 13821 39724 13855
rect 39672 13812 39724 13821
rect 39856 13855 39908 13864
rect 39856 13821 39865 13855
rect 39865 13821 39899 13855
rect 39899 13821 39908 13855
rect 39856 13812 39908 13821
rect 44824 13812 44876 13864
rect 47032 13812 47084 13864
rect 49056 13880 49108 13932
rect 49424 13923 49476 13932
rect 49424 13889 49433 13923
rect 49433 13889 49467 13923
rect 49467 13889 49476 13923
rect 49424 13880 49476 13889
rect 60096 13948 60148 14000
rect 64972 13948 65024 14000
rect 66904 13948 66956 14000
rect 69572 13948 69624 14000
rect 59912 13923 59964 13932
rect 59912 13889 59921 13923
rect 59921 13889 59955 13923
rect 59955 13889 59964 13923
rect 59912 13880 59964 13889
rect 65524 13923 65576 13932
rect 65524 13889 65533 13923
rect 65533 13889 65567 13923
rect 65567 13889 65576 13923
rect 65524 13880 65576 13889
rect 55220 13855 55272 13864
rect 55220 13821 55229 13855
rect 55229 13821 55263 13855
rect 55263 13821 55272 13855
rect 55404 13855 55456 13864
rect 55220 13812 55272 13821
rect 55404 13821 55413 13855
rect 55413 13821 55447 13855
rect 55447 13821 55456 13855
rect 55404 13812 55456 13821
rect 60372 13812 60424 13864
rect 62488 13812 62540 13864
rect 63408 13812 63460 13864
rect 69112 13880 69164 13932
rect 70216 13948 70268 14000
rect 70308 13923 70360 13932
rect 70308 13889 70317 13923
rect 70317 13889 70351 13923
rect 70351 13889 70360 13923
rect 70308 13880 70360 13889
rect 67640 13812 67692 13864
rect 69020 13812 69072 13864
rect 69848 13812 69900 13864
rect 72516 13812 72568 13864
rect 38752 13787 38804 13796
rect 38752 13753 38761 13787
rect 38761 13753 38795 13787
rect 38795 13753 38804 13787
rect 38752 13744 38804 13753
rect 41420 13744 41472 13796
rect 47768 13744 47820 13796
rect 48412 13744 48464 13796
rect 35348 13676 35400 13728
rect 40132 13676 40184 13728
rect 49516 13676 49568 13728
rect 50620 13676 50672 13728
rect 56692 13676 56744 13728
rect 60832 13676 60884 13728
rect 62488 13676 62540 13728
rect 65156 13676 65208 13728
rect 66260 13676 66312 13728
rect 68008 13676 68060 13728
rect 68652 13676 68704 13728
rect 19606 13574 19658 13626
rect 19670 13574 19722 13626
rect 19734 13574 19786 13626
rect 19798 13574 19850 13626
rect 50326 13574 50378 13626
rect 50390 13574 50442 13626
rect 50454 13574 50506 13626
rect 50518 13574 50570 13626
rect 81046 13574 81098 13626
rect 81110 13574 81162 13626
rect 81174 13574 81226 13626
rect 81238 13574 81290 13626
rect 111766 13574 111818 13626
rect 111830 13574 111882 13626
rect 111894 13574 111946 13626
rect 111958 13574 112010 13626
rect 142486 13574 142538 13626
rect 142550 13574 142602 13626
rect 142614 13574 142666 13626
rect 142678 13574 142730 13626
rect 173206 13574 173258 13626
rect 173270 13574 173322 13626
rect 173334 13574 173386 13626
rect 173398 13574 173450 13626
rect 32220 13515 32272 13524
rect 32220 13481 32229 13515
rect 32229 13481 32263 13515
rect 32263 13481 32272 13515
rect 32220 13472 32272 13481
rect 38200 13472 38252 13524
rect 42800 13472 42852 13524
rect 44732 13515 44784 13524
rect 44732 13481 44741 13515
rect 44741 13481 44775 13515
rect 44775 13481 44784 13515
rect 44732 13472 44784 13481
rect 47584 13515 47636 13524
rect 47584 13481 47593 13515
rect 47593 13481 47627 13515
rect 47627 13481 47636 13515
rect 47584 13472 47636 13481
rect 52736 13472 52788 13524
rect 55312 13515 55364 13524
rect 55312 13481 55321 13515
rect 55321 13481 55355 13515
rect 55355 13481 55364 13515
rect 55312 13472 55364 13481
rect 58256 13472 58308 13524
rect 30840 13379 30892 13388
rect 30840 13345 30849 13379
rect 30849 13345 30883 13379
rect 30883 13345 30892 13379
rect 30840 13336 30892 13345
rect 43444 13447 43496 13456
rect 43444 13413 43453 13447
rect 43453 13413 43487 13447
rect 43487 13413 43496 13447
rect 43444 13404 43496 13413
rect 44640 13447 44692 13456
rect 44640 13413 44649 13447
rect 44649 13413 44683 13447
rect 44683 13413 44692 13447
rect 44640 13404 44692 13413
rect 59912 13472 59964 13524
rect 65248 13472 65300 13524
rect 66260 13472 66312 13524
rect 72424 13472 72476 13524
rect 33232 13336 33284 13388
rect 33968 13379 34020 13388
rect 33968 13345 33977 13379
rect 33977 13345 34011 13379
rect 34011 13345 34020 13379
rect 33968 13336 34020 13345
rect 42800 13336 42852 13388
rect 45468 13336 45520 13388
rect 34520 13268 34572 13320
rect 36176 13268 36228 13320
rect 38568 13268 38620 13320
rect 40960 13311 41012 13320
rect 40960 13277 40969 13311
rect 40969 13277 41003 13311
rect 41003 13277 41012 13311
rect 40960 13268 41012 13277
rect 41604 13268 41656 13320
rect 43628 13311 43680 13320
rect 43628 13277 43637 13311
rect 43637 13277 43671 13311
rect 43671 13277 43680 13311
rect 43628 13268 43680 13277
rect 44824 13311 44876 13320
rect 44824 13277 44833 13311
rect 44833 13277 44867 13311
rect 44867 13277 44876 13311
rect 44824 13268 44876 13277
rect 46480 13311 46532 13320
rect 46480 13277 46489 13311
rect 46489 13277 46523 13311
rect 46523 13277 46532 13311
rect 46480 13268 46532 13277
rect 48780 13336 48832 13388
rect 52276 13336 52328 13388
rect 53196 13336 53248 13388
rect 55220 13379 55272 13388
rect 55220 13345 55229 13379
rect 55229 13345 55263 13379
rect 55263 13345 55272 13379
rect 55220 13336 55272 13345
rect 57152 13336 57204 13388
rect 57520 13379 57572 13388
rect 57520 13345 57529 13379
rect 57529 13345 57563 13379
rect 57563 13345 57572 13379
rect 57520 13336 57572 13345
rect 49424 13268 49476 13320
rect 57612 13268 57664 13320
rect 72240 13404 72292 13456
rect 57980 13336 58032 13388
rect 65340 13336 65392 13388
rect 70308 13336 70360 13388
rect 71136 13379 71188 13388
rect 71136 13345 71145 13379
rect 71145 13345 71179 13379
rect 71179 13345 71188 13379
rect 71136 13336 71188 13345
rect 73068 13336 73120 13388
rect 33232 13200 33284 13252
rect 41972 13200 42024 13252
rect 56692 13200 56744 13252
rect 57888 13200 57940 13252
rect 60832 13268 60884 13320
rect 61844 13268 61896 13320
rect 63408 13311 63460 13320
rect 63408 13277 63417 13311
rect 63417 13277 63451 13311
rect 63451 13277 63460 13311
rect 63408 13268 63460 13277
rect 64604 13311 64656 13320
rect 64604 13277 64613 13311
rect 64613 13277 64647 13311
rect 64647 13277 64656 13311
rect 64604 13268 64656 13277
rect 64880 13311 64932 13320
rect 64880 13277 64889 13311
rect 64889 13277 64923 13311
rect 64923 13277 64932 13311
rect 64880 13268 64932 13277
rect 66628 13268 66680 13320
rect 67456 13311 67508 13320
rect 67456 13277 67465 13311
rect 67465 13277 67499 13311
rect 67499 13277 67508 13311
rect 67456 13268 67508 13277
rect 70216 13268 70268 13320
rect 35900 13132 35952 13184
rect 44456 13132 44508 13184
rect 48596 13132 48648 13184
rect 54668 13132 54720 13184
rect 54944 13132 54996 13184
rect 57520 13132 57572 13184
rect 58716 13132 58768 13184
rect 60280 13200 60332 13252
rect 60096 13132 60148 13184
rect 67088 13132 67140 13184
rect 69756 13200 69808 13252
rect 73896 13268 73948 13320
rect 70124 13132 70176 13184
rect 70676 13132 70728 13184
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 34966 13030 35018 13082
rect 35030 13030 35082 13082
rect 35094 13030 35146 13082
rect 35158 13030 35210 13082
rect 65686 13030 65738 13082
rect 65750 13030 65802 13082
rect 65814 13030 65866 13082
rect 65878 13030 65930 13082
rect 96406 13030 96458 13082
rect 96470 13030 96522 13082
rect 96534 13030 96586 13082
rect 96598 13030 96650 13082
rect 127126 13030 127178 13082
rect 127190 13030 127242 13082
rect 127254 13030 127306 13082
rect 127318 13030 127370 13082
rect 157846 13030 157898 13082
rect 157910 13030 157962 13082
rect 157974 13030 158026 13082
rect 158038 13030 158090 13082
rect 32036 12971 32088 12980
rect 32036 12937 32045 12971
rect 32045 12937 32079 12971
rect 32079 12937 32088 12971
rect 32036 12928 32088 12937
rect 34612 12971 34664 12980
rect 34612 12937 34621 12971
rect 34621 12937 34655 12971
rect 34655 12937 34664 12971
rect 34612 12928 34664 12937
rect 36084 12928 36136 12980
rect 38752 12928 38804 12980
rect 39212 12928 39264 12980
rect 41512 12928 41564 12980
rect 42616 12928 42668 12980
rect 44640 12928 44692 12980
rect 45652 12971 45704 12980
rect 45652 12937 45661 12971
rect 45661 12937 45695 12971
rect 45695 12937 45704 12971
rect 45652 12928 45704 12937
rect 57152 12928 57204 12980
rect 58532 12928 58584 12980
rect 30840 12792 30892 12844
rect 33508 12792 33560 12844
rect 36176 12792 36228 12844
rect 37004 12792 37056 12844
rect 40960 12792 41012 12844
rect 45468 12792 45520 12844
rect 45836 12792 45888 12844
rect 47032 12835 47084 12844
rect 47032 12801 47041 12835
rect 47041 12801 47075 12835
rect 47075 12801 47084 12835
rect 47032 12792 47084 12801
rect 47952 12792 48004 12844
rect 32956 12724 33008 12776
rect 33324 12767 33376 12776
rect 33324 12733 33333 12767
rect 33333 12733 33367 12767
rect 33367 12733 33376 12767
rect 33324 12724 33376 12733
rect 37188 12724 37240 12776
rect 38752 12767 38804 12776
rect 38752 12733 38761 12767
rect 38761 12733 38795 12767
rect 38795 12733 38804 12767
rect 38752 12724 38804 12733
rect 40868 12767 40920 12776
rect 40868 12733 40877 12767
rect 40877 12733 40911 12767
rect 40911 12733 40920 12767
rect 40868 12724 40920 12733
rect 44548 12767 44600 12776
rect 44548 12733 44557 12767
rect 44557 12733 44591 12767
rect 44591 12733 44600 12767
rect 44548 12724 44600 12733
rect 47124 12724 47176 12776
rect 47584 12724 47636 12776
rect 48780 12767 48832 12776
rect 48780 12733 48789 12767
rect 48789 12733 48823 12767
rect 48823 12733 48832 12767
rect 56692 12792 56744 12844
rect 57060 12792 57112 12844
rect 57612 12835 57664 12844
rect 57612 12801 57621 12835
rect 57621 12801 57655 12835
rect 57655 12801 57664 12835
rect 57612 12792 57664 12801
rect 57888 12792 57940 12844
rect 48780 12724 48832 12733
rect 50988 12724 51040 12776
rect 55128 12767 55180 12776
rect 55128 12733 55137 12767
rect 55137 12733 55171 12767
rect 55171 12733 55180 12767
rect 55128 12724 55180 12733
rect 59820 12767 59872 12776
rect 59820 12733 59829 12767
rect 59829 12733 59863 12767
rect 59863 12733 59872 12767
rect 59820 12724 59872 12733
rect 63960 12928 64012 12980
rect 67272 12928 67324 12980
rect 63408 12835 63460 12844
rect 63408 12801 63417 12835
rect 63417 12801 63451 12835
rect 63451 12801 63460 12835
rect 63408 12792 63460 12801
rect 66628 12835 66680 12844
rect 66628 12801 66637 12835
rect 66637 12801 66671 12835
rect 66671 12801 66680 12835
rect 66628 12792 66680 12801
rect 68008 12792 68060 12844
rect 69388 12792 69440 12844
rect 70216 12792 70268 12844
rect 63684 12724 63736 12776
rect 64052 12724 64104 12776
rect 64604 12724 64656 12776
rect 64788 12767 64840 12776
rect 64788 12733 64797 12767
rect 64797 12733 64831 12767
rect 64831 12733 64840 12767
rect 64788 12724 64840 12733
rect 65524 12724 65576 12776
rect 70124 12767 70176 12776
rect 70124 12733 70133 12767
rect 70133 12733 70167 12767
rect 70167 12733 70176 12767
rect 70124 12724 70176 12733
rect 72976 12724 73028 12776
rect 50620 12656 50672 12708
rect 62488 12656 62540 12708
rect 63500 12656 63552 12708
rect 70032 12656 70084 12708
rect 46112 12588 46164 12640
rect 52276 12631 52328 12640
rect 52276 12597 52285 12631
rect 52285 12597 52319 12631
rect 52319 12597 52328 12631
rect 52276 12588 52328 12597
rect 56968 12631 57020 12640
rect 56968 12597 56977 12631
rect 56977 12597 57011 12631
rect 57011 12597 57020 12631
rect 56968 12588 57020 12597
rect 58072 12588 58124 12640
rect 61292 12588 61344 12640
rect 65064 12588 65116 12640
rect 68468 12588 68520 12640
rect 19606 12486 19658 12538
rect 19670 12486 19722 12538
rect 19734 12486 19786 12538
rect 19798 12486 19850 12538
rect 50326 12486 50378 12538
rect 50390 12486 50442 12538
rect 50454 12486 50506 12538
rect 50518 12486 50570 12538
rect 81046 12486 81098 12538
rect 81110 12486 81162 12538
rect 81174 12486 81226 12538
rect 81238 12486 81290 12538
rect 111766 12486 111818 12538
rect 111830 12486 111882 12538
rect 111894 12486 111946 12538
rect 111958 12486 112010 12538
rect 142486 12486 142538 12538
rect 142550 12486 142602 12538
rect 142614 12486 142666 12538
rect 142678 12486 142730 12538
rect 173206 12486 173258 12538
rect 173270 12486 173322 12538
rect 173334 12486 173386 12538
rect 173398 12486 173450 12538
rect 34796 12384 34848 12436
rect 34520 12316 34572 12368
rect 35440 12316 35492 12368
rect 60372 12427 60424 12436
rect 60372 12393 60381 12427
rect 60381 12393 60415 12427
rect 60415 12393 60424 12427
rect 60372 12384 60424 12393
rect 36084 12291 36136 12300
rect 36084 12257 36093 12291
rect 36093 12257 36127 12291
rect 36127 12257 36136 12291
rect 36084 12248 36136 12257
rect 37004 12291 37056 12300
rect 37004 12257 37013 12291
rect 37013 12257 37047 12291
rect 37047 12257 37056 12291
rect 37004 12248 37056 12257
rect 44916 12248 44968 12300
rect 45468 12248 45520 12300
rect 56692 12291 56744 12300
rect 56692 12257 56701 12291
rect 56701 12257 56735 12291
rect 56735 12257 56744 12291
rect 56692 12248 56744 12257
rect 62948 12316 63000 12368
rect 36544 12180 36596 12232
rect 42432 12180 42484 12232
rect 47216 12180 47268 12232
rect 55772 12180 55824 12232
rect 37004 12112 37056 12164
rect 35532 12044 35584 12096
rect 48412 12087 48464 12096
rect 48412 12053 48421 12087
rect 48421 12053 48455 12087
rect 48455 12053 48464 12087
rect 48412 12044 48464 12053
rect 58072 12087 58124 12096
rect 58072 12053 58081 12087
rect 58081 12053 58115 12087
rect 58115 12053 58124 12087
rect 58072 12044 58124 12053
rect 61660 12044 61712 12096
rect 62120 12180 62172 12232
rect 64052 12223 64104 12232
rect 64052 12189 64061 12223
rect 64061 12189 64095 12223
rect 64095 12189 64104 12223
rect 64052 12180 64104 12189
rect 66076 12316 66128 12368
rect 66628 12180 66680 12232
rect 93952 12248 94004 12300
rect 63868 12044 63920 12096
rect 65156 12044 65208 12096
rect 65340 12044 65392 12096
rect 67180 12044 67232 12096
rect 69664 12223 69716 12232
rect 69664 12189 69673 12223
rect 69673 12189 69707 12223
rect 69707 12189 69716 12223
rect 69664 12180 69716 12189
rect 68652 12087 68704 12096
rect 68652 12053 68661 12087
rect 68661 12053 68695 12087
rect 68695 12053 68704 12087
rect 68652 12044 68704 12053
rect 69848 12044 69900 12096
rect 70952 12087 71004 12096
rect 70952 12053 70961 12087
rect 70961 12053 70995 12087
rect 70995 12053 71004 12087
rect 70952 12044 71004 12053
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 34966 11942 35018 11994
rect 35030 11942 35082 11994
rect 35094 11942 35146 11994
rect 35158 11942 35210 11994
rect 65686 11942 65738 11994
rect 65750 11942 65802 11994
rect 65814 11942 65866 11994
rect 65878 11942 65930 11994
rect 96406 11942 96458 11994
rect 96470 11942 96522 11994
rect 96534 11942 96586 11994
rect 96598 11942 96650 11994
rect 127126 11942 127178 11994
rect 127190 11942 127242 11994
rect 127254 11942 127306 11994
rect 127318 11942 127370 11994
rect 157846 11942 157898 11994
rect 157910 11942 157962 11994
rect 157974 11942 158026 11994
rect 158038 11942 158090 11994
rect 61660 11883 61712 11892
rect 61660 11849 61669 11883
rect 61669 11849 61703 11883
rect 61703 11849 61712 11883
rect 61660 11840 61712 11849
rect 57888 11704 57940 11756
rect 63592 11704 63644 11756
rect 65984 11704 66036 11756
rect 59544 11679 59596 11688
rect 59544 11645 59553 11679
rect 59553 11645 59587 11679
rect 59587 11645 59596 11679
rect 59544 11636 59596 11645
rect 60372 11636 60424 11688
rect 64052 11636 64104 11688
rect 67180 11679 67232 11688
rect 67180 11645 67189 11679
rect 67189 11645 67223 11679
rect 67223 11645 67232 11679
rect 67180 11636 67232 11645
rect 60280 11500 60332 11552
rect 60556 11500 60608 11552
rect 66260 11500 66312 11552
rect 68560 11543 68612 11552
rect 68560 11509 68569 11543
rect 68569 11509 68603 11543
rect 68603 11509 68612 11543
rect 68560 11500 68612 11509
rect 19606 11398 19658 11450
rect 19670 11398 19722 11450
rect 19734 11398 19786 11450
rect 19798 11398 19850 11450
rect 50326 11398 50378 11450
rect 50390 11398 50442 11450
rect 50454 11398 50506 11450
rect 50518 11398 50570 11450
rect 81046 11398 81098 11450
rect 81110 11398 81162 11450
rect 81174 11398 81226 11450
rect 81238 11398 81290 11450
rect 111766 11398 111818 11450
rect 111830 11398 111882 11450
rect 111894 11398 111946 11450
rect 111958 11398 112010 11450
rect 142486 11398 142538 11450
rect 142550 11398 142602 11450
rect 142614 11398 142666 11450
rect 142678 11398 142730 11450
rect 173206 11398 173258 11450
rect 173270 11398 173322 11450
rect 173334 11398 173386 11450
rect 173398 11398 173450 11450
rect 70400 11296 70452 11348
rect 71136 11296 71188 11348
rect 67180 11160 67232 11212
rect 67548 11092 67600 11144
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 34966 10854 35018 10906
rect 35030 10854 35082 10906
rect 35094 10854 35146 10906
rect 35158 10854 35210 10906
rect 65686 10854 65738 10906
rect 65750 10854 65802 10906
rect 65814 10854 65866 10906
rect 65878 10854 65930 10906
rect 96406 10854 96458 10906
rect 96470 10854 96522 10906
rect 96534 10854 96586 10906
rect 96598 10854 96650 10906
rect 127126 10854 127178 10906
rect 127190 10854 127242 10906
rect 127254 10854 127306 10906
rect 127318 10854 127370 10906
rect 157846 10854 157898 10906
rect 157910 10854 157962 10906
rect 157974 10854 158026 10906
rect 158038 10854 158090 10906
rect 33232 10752 33284 10804
rect 33784 10752 33836 10804
rect 33600 10548 33652 10600
rect 34244 10548 34296 10600
rect 60372 10591 60424 10600
rect 60372 10557 60381 10591
rect 60381 10557 60415 10591
rect 60415 10557 60424 10591
rect 60372 10548 60424 10557
rect 65432 10548 65484 10600
rect 33784 10480 33836 10532
rect 35808 10480 35860 10532
rect 19606 10310 19658 10362
rect 19670 10310 19722 10362
rect 19734 10310 19786 10362
rect 19798 10310 19850 10362
rect 50326 10310 50378 10362
rect 50390 10310 50442 10362
rect 50454 10310 50506 10362
rect 50518 10310 50570 10362
rect 81046 10310 81098 10362
rect 81110 10310 81162 10362
rect 81174 10310 81226 10362
rect 81238 10310 81290 10362
rect 111766 10310 111818 10362
rect 111830 10310 111882 10362
rect 111894 10310 111946 10362
rect 111958 10310 112010 10362
rect 142486 10310 142538 10362
rect 142550 10310 142602 10362
rect 142614 10310 142666 10362
rect 142678 10310 142730 10362
rect 173206 10310 173258 10362
rect 173270 10310 173322 10362
rect 173334 10310 173386 10362
rect 173398 10310 173450 10362
rect 32680 10208 32732 10260
rect 31668 10140 31720 10192
rect 33600 10208 33652 10260
rect 32956 10183 33008 10192
rect 32956 10149 32965 10183
rect 32965 10149 32999 10183
rect 32999 10149 33008 10183
rect 32956 10140 33008 10149
rect 33324 10140 33376 10192
rect 38752 10140 38804 10192
rect 41604 10183 41656 10192
rect 33600 10115 33652 10124
rect 33600 10081 33609 10115
rect 33609 10081 33643 10115
rect 33643 10081 33652 10115
rect 33600 10072 33652 10081
rect 39764 10115 39816 10124
rect 34704 10004 34756 10056
rect 39764 10081 39773 10115
rect 39773 10081 39807 10115
rect 39807 10081 39816 10115
rect 41604 10149 41613 10183
rect 41613 10149 41647 10183
rect 41647 10149 41656 10183
rect 41604 10140 41656 10149
rect 44548 10140 44600 10192
rect 46480 10140 46532 10192
rect 47952 10183 48004 10192
rect 47952 10149 47961 10183
rect 47961 10149 47995 10183
rect 47995 10149 48004 10183
rect 47952 10140 48004 10149
rect 39764 10072 39816 10081
rect 46204 10115 46256 10124
rect 40776 10004 40828 10056
rect 42524 10004 42576 10056
rect 34428 9936 34480 9988
rect 46204 10081 46213 10115
rect 46213 10081 46247 10115
rect 46247 10081 46256 10115
rect 46204 10072 46256 10081
rect 47032 10072 47084 10124
rect 47768 10115 47820 10124
rect 47768 10081 47777 10115
rect 47777 10081 47811 10115
rect 47811 10081 47820 10115
rect 47768 10072 47820 10081
rect 56508 10072 56560 10124
rect 60372 10140 60424 10192
rect 64880 10140 64932 10192
rect 67548 10140 67600 10192
rect 46940 10004 46992 10056
rect 63684 10072 63736 10124
rect 64604 10004 64656 10056
rect 65432 10004 65484 10056
rect 45284 9936 45336 9988
rect 60096 9936 60148 9988
rect 56876 9911 56928 9920
rect 56876 9877 56885 9911
rect 56885 9877 56919 9911
rect 56919 9877 56928 9911
rect 56876 9868 56928 9877
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 34966 9766 35018 9818
rect 35030 9766 35082 9818
rect 35094 9766 35146 9818
rect 35158 9766 35210 9818
rect 65686 9766 65738 9818
rect 65750 9766 65802 9818
rect 65814 9766 65866 9818
rect 65878 9766 65930 9818
rect 96406 9766 96458 9818
rect 96470 9766 96522 9818
rect 96534 9766 96586 9818
rect 96598 9766 96650 9818
rect 127126 9766 127178 9818
rect 127190 9766 127242 9818
rect 127254 9766 127306 9818
rect 127318 9766 127370 9818
rect 157846 9766 157898 9818
rect 157910 9766 157962 9818
rect 157974 9766 158026 9818
rect 158038 9766 158090 9818
rect 37188 9596 37240 9648
rect 38568 9596 38620 9648
rect 40868 9639 40920 9648
rect 40868 9605 40877 9639
rect 40877 9605 40911 9639
rect 40911 9605 40920 9639
rect 40868 9596 40920 9605
rect 42432 9639 42484 9648
rect 42432 9605 42441 9639
rect 42441 9605 42475 9639
rect 42475 9605 42484 9639
rect 42432 9596 42484 9605
rect 47216 9639 47268 9648
rect 47216 9605 47225 9639
rect 47225 9605 47259 9639
rect 47259 9605 47268 9639
rect 47216 9596 47268 9605
rect 50988 9596 51040 9648
rect 55128 9596 55180 9648
rect 57980 9596 58032 9648
rect 59820 9596 59872 9648
rect 29092 9460 29144 9512
rect 32036 9460 32088 9512
rect 36268 9460 36320 9512
rect 39764 9460 39816 9512
rect 47768 9460 47820 9512
rect 49700 9528 49752 9580
rect 50620 9528 50672 9580
rect 54484 9528 54536 9580
rect 55404 9528 55456 9580
rect 56508 9528 56560 9580
rect 59544 9528 59596 9580
rect 72516 9596 72568 9648
rect 63592 9571 63644 9580
rect 56876 9460 56928 9512
rect 30196 9392 30248 9444
rect 36084 9392 36136 9444
rect 37372 9392 37424 9444
rect 38384 9392 38436 9444
rect 37740 9324 37792 9376
rect 40592 9392 40644 9444
rect 46664 9392 46716 9444
rect 49424 9392 49476 9444
rect 53472 9392 53524 9444
rect 56232 9435 56284 9444
rect 56232 9401 56241 9435
rect 56241 9401 56275 9435
rect 56275 9401 56284 9435
rect 56232 9392 56284 9401
rect 57060 9435 57112 9444
rect 57060 9401 57069 9435
rect 57069 9401 57103 9435
rect 57103 9401 57112 9435
rect 57060 9392 57112 9401
rect 57980 9435 58032 9444
rect 57980 9401 57989 9435
rect 57989 9401 58023 9435
rect 58023 9401 58032 9435
rect 57980 9392 58032 9401
rect 42432 9324 42484 9376
rect 54760 9324 54812 9376
rect 63592 9537 63601 9571
rect 63601 9537 63635 9571
rect 63635 9537 63644 9571
rect 63592 9528 63644 9537
rect 65984 9528 66036 9580
rect 60096 9460 60148 9512
rect 60648 9460 60700 9512
rect 64512 9460 64564 9512
rect 61844 9435 61896 9444
rect 61844 9401 61853 9435
rect 61853 9401 61887 9435
rect 61887 9401 61896 9435
rect 61844 9392 61896 9401
rect 63224 9435 63276 9444
rect 63224 9401 63233 9435
rect 63233 9401 63267 9435
rect 63267 9401 63276 9435
rect 63224 9392 63276 9401
rect 65248 9435 65300 9444
rect 65248 9401 65257 9435
rect 65257 9401 65291 9435
rect 65291 9401 65300 9435
rect 65248 9392 65300 9401
rect 65432 9503 65484 9512
rect 65432 9469 65441 9503
rect 65441 9469 65475 9503
rect 65475 9469 65484 9503
rect 65432 9460 65484 9469
rect 65800 9460 65852 9512
rect 67456 9528 67508 9580
rect 69664 9460 69716 9512
rect 64788 9324 64840 9376
rect 65340 9324 65392 9376
rect 19606 9222 19658 9274
rect 19670 9222 19722 9274
rect 19734 9222 19786 9274
rect 19798 9222 19850 9274
rect 50326 9222 50378 9274
rect 50390 9222 50442 9274
rect 50454 9222 50506 9274
rect 50518 9222 50570 9274
rect 81046 9222 81098 9274
rect 81110 9222 81162 9274
rect 81174 9222 81226 9274
rect 81238 9222 81290 9274
rect 111766 9222 111818 9274
rect 111830 9222 111882 9274
rect 111894 9222 111946 9274
rect 111958 9222 112010 9274
rect 142486 9222 142538 9274
rect 142550 9222 142602 9274
rect 142614 9222 142666 9274
rect 142678 9222 142730 9274
rect 173206 9222 173258 9274
rect 173270 9222 173322 9274
rect 173334 9222 173386 9274
rect 173398 9222 173450 9274
rect 48412 9120 48464 9172
rect 52092 9120 52144 9172
rect 41052 9052 41104 9104
rect 61660 9120 61712 9172
rect 32588 9027 32640 9036
rect 32588 8993 32597 9027
rect 32597 8993 32631 9027
rect 32631 8993 32640 9027
rect 32588 8984 32640 8993
rect 30932 8916 30984 8968
rect 31392 8848 31444 8900
rect 33876 8984 33928 9036
rect 40684 8984 40736 9036
rect 54760 8984 54812 9036
rect 55036 8984 55088 9036
rect 56876 8984 56928 9036
rect 59544 8984 59596 9036
rect 60648 8984 60700 9036
rect 61476 8984 61528 9036
rect 63316 9027 63368 9036
rect 63316 8993 63325 9027
rect 63325 8993 63359 9027
rect 63359 8993 63368 9027
rect 63316 8984 63368 8993
rect 65524 9052 65576 9104
rect 66076 9052 66128 9104
rect 63592 8984 63644 9036
rect 65800 9027 65852 9036
rect 65800 8993 65809 9027
rect 65809 8993 65843 9027
rect 65843 8993 65852 9027
rect 65800 8984 65852 8993
rect 55772 8959 55824 8968
rect 55772 8925 55781 8959
rect 55781 8925 55815 8959
rect 55815 8925 55824 8959
rect 55772 8916 55824 8925
rect 62028 8916 62080 8968
rect 62948 8916 63000 8968
rect 65064 8916 65116 8968
rect 66996 8916 67048 8968
rect 38476 8848 38528 8900
rect 41420 8848 41472 8900
rect 33232 8780 33284 8832
rect 33416 8780 33468 8832
rect 49700 8780 49752 8832
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 34966 8678 35018 8730
rect 35030 8678 35082 8730
rect 35094 8678 35146 8730
rect 35158 8678 35210 8730
rect 65686 8678 65738 8730
rect 65750 8678 65802 8730
rect 65814 8678 65866 8730
rect 65878 8678 65930 8730
rect 96406 8678 96458 8730
rect 96470 8678 96522 8730
rect 96534 8678 96586 8730
rect 96598 8678 96650 8730
rect 127126 8678 127178 8730
rect 127190 8678 127242 8730
rect 127254 8678 127306 8730
rect 127318 8678 127370 8730
rect 157846 8678 157898 8730
rect 157910 8678 157962 8730
rect 157974 8678 158026 8730
rect 158038 8678 158090 8730
rect 33600 8576 33652 8628
rect 41328 8576 41380 8628
rect 41420 8619 41472 8628
rect 41420 8585 41429 8619
rect 41429 8585 41463 8619
rect 41463 8585 41472 8619
rect 41420 8576 41472 8585
rect 41604 8576 41656 8628
rect 67640 8576 67692 8628
rect 33692 8508 33744 8560
rect 35624 8508 35676 8560
rect 70032 8508 70084 8560
rect 31668 8440 31720 8492
rect 31852 8372 31904 8424
rect 32588 8372 32640 8424
rect 33048 8372 33100 8424
rect 33416 8415 33468 8424
rect 33416 8381 33425 8415
rect 33425 8381 33459 8415
rect 33459 8381 33468 8415
rect 33416 8372 33468 8381
rect 33876 8372 33928 8424
rect 35900 8440 35952 8492
rect 38292 8440 38344 8492
rect 39856 8440 39908 8492
rect 39304 8372 39356 8424
rect 40868 8415 40920 8424
rect 40868 8381 40877 8415
rect 40877 8381 40911 8415
rect 40911 8381 40920 8415
rect 40868 8372 40920 8381
rect 41052 8415 41104 8424
rect 41052 8381 41061 8415
rect 41061 8381 41095 8415
rect 41095 8381 41104 8415
rect 41052 8372 41104 8381
rect 41236 8415 41288 8424
rect 41236 8381 41245 8415
rect 41245 8381 41279 8415
rect 41279 8381 41288 8415
rect 41236 8372 41288 8381
rect 31944 8304 31996 8356
rect 35900 8347 35952 8356
rect 35900 8313 35909 8347
rect 35909 8313 35943 8347
rect 35943 8313 35952 8347
rect 35900 8304 35952 8313
rect 38660 8304 38712 8356
rect 39488 8304 39540 8356
rect 27804 8236 27856 8288
rect 41052 8236 41104 8288
rect 45560 8372 45612 8424
rect 46020 8372 46072 8424
rect 65064 8440 65116 8492
rect 46296 8415 46348 8424
rect 46296 8381 46305 8415
rect 46305 8381 46339 8415
rect 46339 8381 46348 8415
rect 46296 8372 46348 8381
rect 63132 8372 63184 8424
rect 67272 8372 67324 8424
rect 43260 8304 43312 8356
rect 54300 8304 54352 8356
rect 56968 8304 57020 8356
rect 45928 8236 45980 8288
rect 46572 8236 46624 8288
rect 55680 8236 55732 8288
rect 55772 8236 55824 8288
rect 64420 8304 64472 8356
rect 62304 8236 62356 8288
rect 68652 8236 68704 8288
rect 71320 8236 71372 8288
rect 19606 8134 19658 8186
rect 19670 8134 19722 8186
rect 19734 8134 19786 8186
rect 19798 8134 19850 8186
rect 50326 8134 50378 8186
rect 50390 8134 50442 8186
rect 50454 8134 50506 8186
rect 50518 8134 50570 8186
rect 81046 8134 81098 8186
rect 81110 8134 81162 8186
rect 81174 8134 81226 8186
rect 81238 8134 81290 8186
rect 111766 8134 111818 8186
rect 111830 8134 111882 8186
rect 111894 8134 111946 8186
rect 111958 8134 112010 8186
rect 142486 8134 142538 8186
rect 142550 8134 142602 8186
rect 142614 8134 142666 8186
rect 142678 8134 142730 8186
rect 173206 8134 173258 8186
rect 173270 8134 173322 8186
rect 173334 8134 173386 8186
rect 173398 8134 173450 8186
rect 20996 8007 21048 8016
rect 20996 7973 21005 8007
rect 21005 7973 21039 8007
rect 21039 7973 21048 8007
rect 20996 7964 21048 7973
rect 21272 7964 21324 8016
rect 24216 7964 24268 8016
rect 31576 8032 31628 8084
rect 33600 8075 33652 8084
rect 21180 7939 21232 7948
rect 21180 7905 21189 7939
rect 21189 7905 21223 7939
rect 21223 7905 21232 7939
rect 25596 7939 25648 7948
rect 21180 7896 21232 7905
rect 25596 7905 25605 7939
rect 25605 7905 25639 7939
rect 25639 7905 25648 7939
rect 25596 7896 25648 7905
rect 27804 8007 27856 8016
rect 27804 7973 27813 8007
rect 27813 7973 27847 8007
rect 27847 7973 27856 8007
rect 27804 7964 27856 7973
rect 28172 7964 28224 8016
rect 29920 7964 29972 8016
rect 30380 7964 30432 8016
rect 25964 7939 26016 7948
rect 25964 7905 25973 7939
rect 25973 7905 26007 7939
rect 26007 7905 26016 7939
rect 25964 7896 26016 7905
rect 26424 7896 26476 7948
rect 27620 7939 27672 7948
rect 27620 7905 27629 7939
rect 27629 7905 27663 7939
rect 27663 7905 27672 7939
rect 27896 7939 27948 7948
rect 27620 7896 27672 7905
rect 27896 7905 27905 7939
rect 27905 7905 27939 7939
rect 27939 7905 27948 7939
rect 27896 7896 27948 7905
rect 20996 7828 21048 7880
rect 28264 7896 28316 7948
rect 29368 7896 29420 7948
rect 30472 7939 30524 7948
rect 30472 7905 30481 7939
rect 30481 7905 30515 7939
rect 30515 7905 30524 7939
rect 30472 7896 30524 7905
rect 31852 8007 31904 8016
rect 31852 7973 31861 8007
rect 31861 7973 31895 8007
rect 31895 7973 31904 8007
rect 31852 7964 31904 7973
rect 32496 8007 32548 8016
rect 32496 7973 32505 8007
rect 32505 7973 32539 8007
rect 32539 7973 32548 8007
rect 32496 7964 32548 7973
rect 32588 7964 32640 8016
rect 32956 7964 33008 8016
rect 33600 8041 33609 8075
rect 33609 8041 33643 8075
rect 33643 8041 33652 8075
rect 33600 8032 33652 8041
rect 33784 8075 33836 8084
rect 33784 8041 33793 8075
rect 33793 8041 33827 8075
rect 33827 8041 33836 8075
rect 33784 8032 33836 8041
rect 33968 8032 34020 8084
rect 39488 8032 39540 8084
rect 31024 7896 31076 7948
rect 31392 7896 31444 7948
rect 31668 7939 31720 7948
rect 31668 7905 31677 7939
rect 31677 7905 31711 7939
rect 31711 7905 31720 7939
rect 31668 7896 31720 7905
rect 32864 7939 32916 7948
rect 32864 7905 32873 7939
rect 32873 7905 32907 7939
rect 32907 7905 32916 7939
rect 32864 7896 32916 7905
rect 28816 7828 28868 7880
rect 29184 7828 29236 7880
rect 33324 7828 33376 7880
rect 26240 7760 26292 7812
rect 28264 7760 28316 7812
rect 20812 7692 20864 7744
rect 23480 7692 23532 7744
rect 26332 7692 26384 7744
rect 29276 7692 29328 7744
rect 34336 7964 34388 8016
rect 36360 7964 36412 8016
rect 38292 8007 38344 8016
rect 38292 7973 38301 8007
rect 38301 7973 38335 8007
rect 38335 7973 38344 8007
rect 38292 7964 38344 7973
rect 38568 7964 38620 8016
rect 39304 7964 39356 8016
rect 46020 8032 46072 8084
rect 46848 8032 46900 8084
rect 35992 7896 36044 7948
rect 37464 7896 37516 7948
rect 40868 7964 40920 8016
rect 41880 8007 41932 8016
rect 41880 7973 41889 8007
rect 41889 7973 41923 8007
rect 41923 7973 41932 8007
rect 41880 7964 41932 7973
rect 41972 8007 42024 8016
rect 41972 7973 41981 8007
rect 41981 7973 42015 8007
rect 42015 7973 42024 8007
rect 41972 7964 42024 7973
rect 43996 7964 44048 8016
rect 46296 7964 46348 8016
rect 33876 7828 33928 7880
rect 33784 7760 33836 7812
rect 36360 7760 36412 7812
rect 39120 7828 39172 7880
rect 39948 7896 40000 7948
rect 40132 7896 40184 7948
rect 40040 7828 40092 7880
rect 41604 7896 41656 7948
rect 41696 7939 41748 7948
rect 41696 7905 41705 7939
rect 41705 7905 41739 7939
rect 41739 7905 41748 7939
rect 41696 7896 41748 7905
rect 41236 7828 41288 7880
rect 44180 7896 44232 7948
rect 46388 7939 46440 7948
rect 46388 7905 46397 7939
rect 46397 7905 46431 7939
rect 46431 7905 46440 7939
rect 46388 7896 46440 7905
rect 46572 7939 46624 7948
rect 46572 7905 46581 7939
rect 46581 7905 46615 7939
rect 46615 7905 46624 7939
rect 46572 7896 46624 7905
rect 45100 7828 45152 7880
rect 47308 7896 47360 7948
rect 47492 7896 47544 7948
rect 47676 7939 47728 7948
rect 47676 7905 47685 7939
rect 47685 7905 47719 7939
rect 47719 7905 47728 7939
rect 47676 7896 47728 7905
rect 47952 7964 48004 8016
rect 48504 7964 48556 8016
rect 55772 8032 55824 8084
rect 55864 8032 55916 8084
rect 60556 8032 60608 8084
rect 48688 8007 48740 8016
rect 48688 7973 48697 8007
rect 48697 7973 48731 8007
rect 48731 7973 48740 8007
rect 48688 7964 48740 7973
rect 54760 7964 54812 8016
rect 58072 7964 58124 8016
rect 59452 7964 59504 8016
rect 48412 7939 48464 7948
rect 48412 7905 48421 7939
rect 48421 7905 48455 7939
rect 48455 7905 48464 7939
rect 48412 7896 48464 7905
rect 49148 7896 49200 7948
rect 49976 7896 50028 7948
rect 62304 7896 62356 7948
rect 63132 8032 63184 8084
rect 65340 8032 65392 8084
rect 63500 7939 63552 7948
rect 63500 7905 63527 7939
rect 63527 7905 63552 7939
rect 63500 7896 63552 7905
rect 46940 7828 46992 7880
rect 56692 7828 56744 7880
rect 62396 7828 62448 7880
rect 62672 7828 62724 7880
rect 62948 7828 63000 7880
rect 63132 7828 63184 7880
rect 64420 7896 64472 7948
rect 68560 7896 68612 7948
rect 72608 7896 72660 7948
rect 64144 7828 64196 7880
rect 65524 7828 65576 7880
rect 36728 7760 36780 7812
rect 40868 7760 40920 7812
rect 40960 7760 41012 7812
rect 41512 7760 41564 7812
rect 46572 7760 46624 7812
rect 47492 7760 47544 7812
rect 50988 7760 51040 7812
rect 55220 7760 55272 7812
rect 56876 7760 56928 7812
rect 61108 7760 61160 7812
rect 62580 7760 62632 7812
rect 62856 7760 62908 7812
rect 64236 7760 64288 7812
rect 70124 7760 70176 7812
rect 70308 7760 70360 7812
rect 39948 7692 40000 7744
rect 40132 7692 40184 7744
rect 40224 7692 40276 7744
rect 44732 7692 44784 7744
rect 47308 7692 47360 7744
rect 48136 7692 48188 7744
rect 48780 7692 48832 7744
rect 49056 7692 49108 7744
rect 65432 7692 65484 7744
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 34966 7590 35018 7642
rect 35030 7590 35082 7642
rect 35094 7590 35146 7642
rect 35158 7590 35210 7642
rect 65686 7590 65738 7642
rect 65750 7590 65802 7642
rect 65814 7590 65866 7642
rect 65878 7590 65930 7642
rect 96406 7590 96458 7642
rect 96470 7590 96522 7642
rect 96534 7590 96586 7642
rect 96598 7590 96650 7642
rect 127126 7590 127178 7642
rect 127190 7590 127242 7642
rect 127254 7590 127306 7642
rect 127318 7590 127370 7642
rect 157846 7590 157898 7642
rect 157910 7590 157962 7642
rect 157974 7590 158026 7642
rect 158038 7590 158090 7642
rect 18604 7327 18656 7336
rect 18604 7293 18613 7327
rect 18613 7293 18647 7327
rect 18647 7293 18656 7327
rect 18604 7284 18656 7293
rect 22192 7488 22244 7540
rect 29644 7531 29696 7540
rect 29644 7497 29653 7531
rect 29653 7497 29687 7531
rect 29687 7497 29696 7531
rect 29644 7488 29696 7497
rect 30472 7488 30524 7540
rect 32128 7488 32180 7540
rect 35808 7531 35860 7540
rect 35808 7497 35817 7531
rect 35817 7497 35851 7531
rect 35851 7497 35860 7531
rect 35808 7488 35860 7497
rect 36176 7488 36228 7540
rect 39396 7488 39448 7540
rect 40776 7488 40828 7540
rect 40960 7488 41012 7540
rect 50896 7488 50948 7540
rect 50988 7488 51040 7540
rect 18972 7327 19024 7336
rect 18972 7293 18981 7327
rect 18981 7293 19015 7327
rect 19015 7293 19024 7327
rect 20168 7327 20220 7336
rect 18972 7284 19024 7293
rect 18052 7216 18104 7268
rect 17960 7148 18012 7200
rect 20168 7293 20177 7327
rect 20177 7293 20211 7327
rect 20211 7293 20220 7327
rect 20168 7284 20220 7293
rect 20444 7259 20496 7268
rect 20444 7225 20453 7259
rect 20453 7225 20487 7259
rect 20487 7225 20496 7259
rect 20444 7216 20496 7225
rect 20904 7284 20956 7336
rect 23020 7327 23072 7336
rect 23020 7293 23029 7327
rect 23029 7293 23063 7327
rect 23063 7293 23072 7327
rect 23020 7284 23072 7293
rect 25964 7352 26016 7404
rect 22008 7216 22060 7268
rect 25596 7284 25648 7336
rect 26424 7284 26476 7336
rect 26516 7327 26568 7336
rect 26516 7293 26525 7327
rect 26525 7293 26559 7327
rect 26559 7293 26568 7327
rect 27436 7352 27488 7404
rect 30748 7420 30800 7472
rect 31576 7420 31628 7472
rect 26516 7284 26568 7293
rect 27620 7284 27672 7336
rect 28448 7327 28500 7336
rect 28448 7293 28457 7327
rect 28457 7293 28491 7327
rect 28491 7293 28500 7327
rect 28448 7284 28500 7293
rect 28540 7284 28592 7336
rect 28908 7284 28960 7336
rect 23204 7259 23256 7268
rect 23204 7225 23213 7259
rect 23213 7225 23247 7259
rect 23247 7225 23256 7259
rect 23204 7216 23256 7225
rect 26240 7216 26292 7268
rect 26608 7259 26660 7268
rect 26608 7225 26617 7259
rect 26617 7225 26651 7259
rect 26651 7225 26660 7259
rect 28724 7259 28776 7268
rect 26608 7216 26660 7225
rect 28724 7225 28733 7259
rect 28733 7225 28767 7259
rect 28767 7225 28776 7259
rect 28724 7216 28776 7225
rect 20720 7191 20772 7200
rect 20720 7157 20729 7191
rect 20729 7157 20763 7191
rect 20763 7157 20772 7191
rect 20720 7148 20772 7157
rect 22284 7148 22336 7200
rect 24952 7191 25004 7200
rect 24952 7157 24961 7191
rect 24961 7157 24995 7191
rect 24995 7157 25004 7191
rect 24952 7148 25004 7157
rect 25044 7148 25096 7200
rect 32772 7352 32824 7404
rect 33048 7352 33100 7404
rect 29920 7284 29972 7336
rect 30656 7284 30708 7336
rect 29184 7216 29236 7268
rect 31300 7284 31352 7336
rect 33784 7352 33836 7404
rect 33508 7327 33560 7336
rect 33508 7293 33517 7327
rect 33517 7293 33551 7327
rect 33551 7293 33560 7327
rect 33508 7284 33560 7293
rect 33876 7284 33928 7336
rect 31116 7216 31168 7268
rect 33600 7259 33652 7268
rect 33600 7225 33609 7259
rect 33609 7225 33643 7259
rect 33643 7225 33652 7259
rect 33600 7216 33652 7225
rect 34060 7284 34112 7336
rect 35256 7327 35308 7336
rect 35256 7293 35265 7327
rect 35265 7293 35299 7327
rect 35299 7293 35308 7327
rect 35256 7284 35308 7293
rect 36360 7327 36412 7336
rect 36360 7293 36369 7327
rect 36369 7293 36403 7327
rect 36403 7293 36412 7327
rect 36360 7284 36412 7293
rect 39488 7420 39540 7472
rect 43996 7420 44048 7472
rect 44180 7463 44232 7472
rect 44180 7429 44189 7463
rect 44189 7429 44223 7463
rect 44223 7429 44232 7463
rect 44180 7420 44232 7429
rect 46296 7420 46348 7472
rect 46572 7420 46624 7472
rect 37096 7352 37148 7404
rect 36728 7327 36780 7336
rect 36728 7293 36737 7327
rect 36737 7293 36771 7327
rect 36771 7293 36780 7327
rect 36728 7284 36780 7293
rect 29092 7148 29144 7200
rect 29276 7148 29328 7200
rect 29368 7148 29420 7200
rect 30564 7148 30616 7200
rect 33048 7148 33100 7200
rect 33324 7148 33376 7200
rect 34796 7259 34848 7268
rect 34796 7225 34805 7259
rect 34805 7225 34839 7259
rect 34839 7225 34848 7259
rect 34796 7216 34848 7225
rect 33876 7191 33928 7200
rect 33876 7157 33885 7191
rect 33885 7157 33919 7191
rect 33919 7157 33928 7191
rect 33876 7148 33928 7157
rect 34152 7191 34204 7200
rect 34152 7157 34161 7191
rect 34161 7157 34195 7191
rect 34195 7157 34204 7191
rect 34152 7148 34204 7157
rect 34244 7148 34296 7200
rect 35624 7191 35676 7200
rect 35624 7157 35633 7191
rect 35633 7157 35667 7191
rect 35667 7157 35676 7191
rect 35624 7148 35676 7157
rect 36452 7216 36504 7268
rect 38660 7327 38712 7336
rect 38660 7293 38669 7327
rect 38669 7293 38703 7327
rect 38703 7293 38712 7327
rect 38660 7284 38712 7293
rect 38844 7284 38896 7336
rect 39764 7352 39816 7404
rect 40868 7352 40920 7404
rect 41236 7352 41288 7404
rect 41696 7327 41748 7336
rect 36820 7148 36872 7200
rect 37280 7148 37332 7200
rect 39580 7259 39632 7268
rect 39580 7225 39589 7259
rect 39589 7225 39623 7259
rect 39623 7225 39632 7259
rect 39580 7216 39632 7225
rect 39672 7216 39724 7268
rect 39948 7259 40000 7268
rect 39948 7225 39957 7259
rect 39957 7225 39991 7259
rect 39991 7225 40000 7259
rect 39948 7216 40000 7225
rect 39488 7148 39540 7200
rect 41696 7293 41705 7327
rect 41705 7293 41739 7327
rect 41739 7293 41748 7327
rect 41696 7284 41748 7293
rect 41880 7327 41932 7336
rect 41880 7293 41889 7327
rect 41889 7293 41923 7327
rect 41923 7293 41932 7327
rect 41880 7284 41932 7293
rect 42156 7284 42208 7336
rect 43628 7327 43680 7336
rect 40684 7259 40736 7268
rect 40684 7225 40693 7259
rect 40693 7225 40727 7259
rect 40727 7225 40736 7259
rect 40684 7216 40736 7225
rect 40776 7216 40828 7268
rect 43628 7293 43637 7327
rect 43637 7293 43671 7327
rect 43671 7293 43680 7327
rect 43628 7284 43680 7293
rect 44916 7352 44968 7404
rect 48688 7352 48740 7404
rect 47584 7284 47636 7336
rect 48412 7284 48464 7336
rect 48872 7284 48924 7336
rect 49056 7352 49108 7404
rect 49240 7420 49292 7472
rect 54760 7420 54812 7472
rect 57060 7488 57112 7540
rect 59268 7488 59320 7540
rect 60188 7488 60240 7540
rect 61292 7488 61344 7540
rect 63316 7488 63368 7540
rect 64604 7531 64656 7540
rect 64604 7497 64613 7531
rect 64613 7497 64647 7531
rect 64647 7497 64656 7531
rect 64604 7488 64656 7497
rect 49148 7327 49200 7336
rect 49148 7293 49157 7327
rect 49157 7293 49191 7327
rect 49191 7293 49200 7327
rect 49148 7284 49200 7293
rect 49332 7284 49384 7336
rect 49976 7327 50028 7336
rect 49976 7293 49985 7327
rect 49985 7293 50019 7327
rect 50019 7293 50028 7327
rect 49976 7284 50028 7293
rect 50160 7327 50212 7336
rect 50160 7293 50169 7327
rect 50169 7293 50203 7327
rect 50203 7293 50212 7327
rect 50160 7284 50212 7293
rect 55128 7352 55180 7404
rect 55496 7395 55548 7404
rect 55496 7361 55505 7395
rect 55505 7361 55539 7395
rect 55539 7361 55548 7395
rect 55496 7352 55548 7361
rect 59912 7420 59964 7472
rect 56600 7352 56652 7404
rect 62279 7395 62331 7404
rect 62279 7361 62301 7395
rect 62301 7361 62331 7395
rect 62279 7352 62331 7361
rect 62764 7352 62816 7404
rect 63316 7395 63368 7404
rect 63316 7361 63325 7395
rect 63325 7361 63359 7395
rect 63359 7361 63368 7395
rect 63316 7352 63368 7361
rect 64788 7352 64840 7404
rect 65064 7352 65116 7404
rect 55220 7284 55272 7336
rect 55772 7327 55824 7336
rect 55772 7293 55799 7327
rect 55799 7293 55824 7327
rect 56048 7327 56100 7336
rect 55772 7284 55824 7293
rect 56048 7293 56057 7327
rect 56057 7293 56091 7327
rect 56091 7293 56100 7327
rect 56048 7284 56100 7293
rect 56692 7284 56744 7336
rect 61384 7284 61436 7336
rect 62120 7327 62172 7336
rect 62120 7293 62129 7327
rect 62129 7293 62163 7327
rect 62163 7293 62172 7327
rect 62377 7327 62429 7336
rect 62120 7284 62172 7293
rect 62377 7293 62386 7327
rect 62386 7293 62420 7327
rect 62420 7293 62429 7327
rect 62377 7284 62429 7293
rect 42248 7191 42300 7200
rect 42248 7157 42257 7191
rect 42257 7157 42291 7191
rect 42291 7157 42300 7191
rect 47676 7259 47728 7268
rect 42248 7148 42300 7157
rect 46940 7148 46992 7200
rect 47676 7225 47685 7259
rect 47685 7225 47719 7259
rect 47719 7225 47728 7259
rect 47676 7216 47728 7225
rect 48228 7216 48280 7268
rect 49332 7191 49384 7200
rect 49332 7157 49341 7191
rect 49341 7157 49375 7191
rect 49375 7157 49384 7191
rect 49332 7148 49384 7157
rect 49608 7216 49660 7268
rect 50620 7148 50672 7200
rect 56600 7216 56652 7268
rect 61568 7216 61620 7268
rect 86592 7284 86644 7336
rect 61200 7148 61252 7200
rect 65524 7259 65576 7268
rect 64788 7191 64840 7200
rect 64788 7157 64797 7191
rect 64797 7157 64831 7191
rect 64831 7157 64840 7191
rect 64788 7148 64840 7157
rect 65524 7225 65533 7259
rect 65533 7225 65567 7259
rect 65567 7225 65576 7259
rect 65524 7216 65576 7225
rect 66076 7216 66128 7268
rect 66260 7216 66312 7268
rect 68100 7216 68152 7268
rect 68284 7148 68336 7200
rect 19606 7046 19658 7098
rect 19670 7046 19722 7098
rect 19734 7046 19786 7098
rect 19798 7046 19850 7098
rect 50326 7046 50378 7098
rect 50390 7046 50442 7098
rect 50454 7046 50506 7098
rect 50518 7046 50570 7098
rect 81046 7046 81098 7098
rect 81110 7046 81162 7098
rect 81174 7046 81226 7098
rect 81238 7046 81290 7098
rect 111766 7046 111818 7098
rect 111830 7046 111882 7098
rect 111894 7046 111946 7098
rect 111958 7046 112010 7098
rect 142486 7046 142538 7098
rect 142550 7046 142602 7098
rect 142614 7046 142666 7098
rect 142678 7046 142730 7098
rect 173206 7046 173258 7098
rect 173270 7046 173322 7098
rect 173334 7046 173386 7098
rect 173398 7046 173450 7098
rect 21088 6987 21140 6996
rect 21088 6953 21097 6987
rect 21097 6953 21131 6987
rect 21131 6953 21140 6987
rect 21088 6944 21140 6953
rect 17960 6808 18012 6860
rect 18604 6876 18656 6928
rect 18696 6851 18748 6860
rect 18696 6817 18705 6851
rect 18705 6817 18739 6851
rect 18739 6817 18748 6851
rect 18696 6808 18748 6817
rect 18604 6740 18656 6792
rect 18972 6808 19024 6860
rect 20168 6808 20220 6860
rect 20536 6851 20588 6860
rect 20536 6817 20545 6851
rect 20545 6817 20579 6851
rect 20579 6817 20588 6851
rect 20536 6808 20588 6817
rect 20628 6808 20680 6860
rect 17408 6672 17460 6724
rect 17316 6604 17368 6656
rect 17960 6604 18012 6656
rect 18052 6604 18104 6656
rect 20536 6672 20588 6724
rect 20904 6851 20956 6860
rect 20904 6817 20913 6851
rect 20913 6817 20947 6851
rect 20947 6817 20956 6851
rect 21732 6919 21784 6928
rect 21732 6885 21741 6919
rect 21741 6885 21775 6919
rect 21775 6885 21784 6919
rect 21732 6876 21784 6885
rect 23204 6944 23256 6996
rect 33324 6944 33376 6996
rect 33508 6944 33560 6996
rect 40960 6944 41012 6996
rect 41144 6987 41196 6996
rect 41144 6953 41153 6987
rect 41153 6953 41187 6987
rect 41187 6953 41196 6987
rect 41144 6944 41196 6953
rect 41236 6944 41288 6996
rect 21548 6851 21600 6860
rect 20904 6808 20956 6817
rect 21548 6817 21557 6851
rect 21557 6817 21591 6851
rect 21591 6817 21600 6851
rect 21548 6808 21600 6817
rect 24952 6876 25004 6928
rect 29184 6876 29236 6928
rect 28908 6808 28960 6860
rect 29368 6851 29420 6860
rect 29368 6817 29377 6851
rect 29377 6817 29411 6851
rect 29411 6817 29420 6851
rect 30564 6851 30616 6860
rect 29368 6808 29420 6817
rect 30564 6817 30573 6851
rect 30573 6817 30607 6851
rect 30607 6817 30616 6851
rect 30564 6808 30616 6817
rect 31024 6876 31076 6928
rect 31208 6876 31260 6928
rect 31484 6876 31536 6928
rect 31760 6919 31812 6928
rect 31760 6885 31769 6919
rect 31769 6885 31803 6919
rect 31803 6885 31812 6919
rect 31760 6876 31812 6885
rect 32956 6808 33008 6860
rect 33140 6808 33192 6860
rect 33508 6808 33560 6860
rect 33784 6851 33836 6860
rect 33784 6817 33793 6851
rect 33793 6817 33827 6851
rect 33827 6817 33836 6851
rect 33784 6808 33836 6817
rect 34060 6808 34112 6860
rect 34796 6876 34848 6928
rect 36820 6876 36872 6928
rect 40040 6876 40092 6928
rect 35992 6851 36044 6860
rect 21732 6672 21784 6724
rect 30288 6740 30340 6792
rect 31024 6740 31076 6792
rect 35992 6817 36001 6851
rect 36001 6817 36035 6851
rect 36035 6817 36044 6851
rect 35992 6808 36044 6817
rect 36636 6851 36688 6860
rect 36636 6817 36645 6851
rect 36645 6817 36679 6851
rect 36679 6817 36688 6851
rect 36636 6808 36688 6817
rect 37648 6851 37700 6860
rect 37648 6817 37682 6851
rect 37682 6817 37700 6851
rect 37648 6808 37700 6817
rect 38568 6808 38620 6860
rect 41880 6944 41932 6996
rect 56600 6944 56652 6996
rect 41696 6808 41748 6860
rect 41880 6851 41932 6860
rect 41880 6817 41889 6851
rect 41889 6817 41923 6851
rect 41923 6817 41932 6851
rect 41880 6808 41932 6817
rect 43536 6808 43588 6860
rect 44456 6851 44508 6860
rect 44456 6817 44490 6851
rect 44490 6817 44508 6851
rect 44640 6851 44692 6860
rect 44456 6808 44508 6817
rect 44640 6817 44649 6851
rect 44649 6817 44683 6851
rect 44683 6817 44692 6851
rect 44640 6808 44692 6817
rect 45284 6851 45336 6860
rect 45284 6817 45293 6851
rect 45293 6817 45327 6851
rect 45327 6817 45336 6851
rect 45284 6808 45336 6817
rect 46388 6808 46440 6860
rect 46664 6851 46716 6860
rect 46664 6817 46673 6851
rect 46673 6817 46707 6851
rect 46707 6817 46716 6851
rect 46664 6808 46716 6817
rect 22100 6715 22152 6724
rect 22100 6681 22109 6715
rect 22109 6681 22143 6715
rect 22143 6681 22152 6715
rect 22100 6672 22152 6681
rect 23020 6672 23072 6724
rect 21180 6604 21232 6656
rect 28540 6604 28592 6656
rect 29184 6604 29236 6656
rect 31300 6672 31352 6724
rect 32680 6715 32732 6724
rect 32680 6681 32689 6715
rect 32689 6681 32723 6715
rect 32723 6681 32732 6715
rect 32680 6672 32732 6681
rect 33140 6672 33192 6724
rect 34888 6672 34940 6724
rect 36544 6672 36596 6724
rect 36728 6740 36780 6792
rect 36912 6740 36964 6792
rect 37188 6740 37240 6792
rect 37832 6783 37884 6792
rect 37832 6749 37841 6783
rect 37841 6749 37875 6783
rect 37875 6749 37884 6783
rect 37832 6740 37884 6749
rect 38384 6740 38436 6792
rect 39764 6740 39816 6792
rect 40868 6740 40920 6792
rect 43628 6783 43680 6792
rect 43628 6749 43637 6783
rect 43637 6749 43671 6783
rect 43671 6749 43680 6783
rect 43628 6740 43680 6749
rect 44364 6783 44416 6792
rect 44364 6749 44373 6783
rect 44373 6749 44407 6783
rect 44407 6749 44416 6783
rect 44364 6740 44416 6749
rect 42432 6715 42484 6724
rect 30840 6604 30892 6656
rect 31392 6604 31444 6656
rect 35900 6604 35952 6656
rect 36820 6604 36872 6656
rect 42432 6681 42441 6715
rect 42441 6681 42475 6715
rect 42475 6681 42484 6715
rect 42432 6672 42484 6681
rect 44088 6715 44140 6724
rect 44088 6681 44097 6715
rect 44097 6681 44131 6715
rect 44131 6681 44140 6715
rect 44088 6672 44140 6681
rect 45376 6672 45428 6724
rect 49976 6876 50028 6928
rect 55680 6876 55732 6928
rect 62028 6944 62080 6996
rect 62580 6944 62632 6996
rect 64604 6944 64656 6996
rect 64788 6944 64840 6996
rect 84844 6944 84896 6996
rect 59912 6876 59964 6928
rect 61108 6876 61160 6928
rect 61384 6876 61436 6928
rect 46848 6851 46900 6860
rect 46848 6817 46857 6851
rect 46857 6817 46891 6851
rect 46891 6817 46900 6851
rect 46848 6808 46900 6817
rect 47216 6808 47268 6860
rect 41144 6604 41196 6656
rect 44456 6604 44508 6656
rect 47124 6740 47176 6792
rect 48596 6851 48648 6860
rect 48596 6817 48630 6851
rect 48630 6817 48648 6851
rect 49424 6851 49476 6860
rect 48596 6808 48648 6817
rect 49424 6817 49433 6851
rect 49433 6817 49467 6851
rect 49467 6817 49476 6851
rect 49424 6808 49476 6817
rect 47952 6740 48004 6792
rect 48504 6783 48556 6792
rect 48504 6749 48513 6783
rect 48513 6749 48547 6783
rect 48547 6749 48556 6783
rect 48504 6740 48556 6749
rect 48780 6783 48832 6792
rect 48780 6749 48789 6783
rect 48789 6749 48823 6783
rect 48823 6749 48832 6783
rect 48780 6740 48832 6749
rect 48964 6740 49016 6792
rect 50068 6851 50120 6860
rect 50068 6817 50077 6851
rect 50077 6817 50111 6851
rect 50111 6817 50120 6851
rect 50252 6851 50304 6860
rect 50068 6808 50120 6817
rect 50252 6817 50261 6851
rect 50261 6817 50295 6851
rect 50295 6817 50304 6851
rect 50252 6808 50304 6817
rect 52828 6851 52880 6860
rect 52828 6817 52837 6851
rect 52837 6817 52871 6851
rect 52871 6817 52880 6851
rect 52828 6808 52880 6817
rect 53472 6851 53524 6860
rect 53472 6817 53481 6851
rect 53481 6817 53515 6851
rect 53515 6817 53524 6851
rect 53472 6808 53524 6817
rect 51816 6783 51868 6792
rect 48596 6604 48648 6656
rect 49516 6604 49568 6656
rect 51816 6749 51825 6783
rect 51825 6749 51859 6783
rect 51859 6749 51868 6783
rect 51816 6740 51868 6749
rect 52552 6783 52604 6792
rect 52552 6749 52561 6783
rect 52561 6749 52595 6783
rect 52595 6749 52604 6783
rect 52552 6740 52604 6749
rect 52184 6672 52236 6724
rect 54024 6740 54076 6792
rect 54944 6851 54996 6860
rect 54944 6817 54978 6851
rect 54978 6817 54996 6851
rect 54944 6808 54996 6817
rect 56232 6808 56284 6860
rect 56876 6808 56928 6860
rect 59176 6851 59228 6860
rect 59176 6817 59185 6851
rect 59185 6817 59219 6851
rect 59219 6817 59228 6851
rect 59176 6808 59228 6817
rect 54668 6740 54720 6792
rect 54852 6783 54904 6792
rect 54852 6749 54861 6783
rect 54861 6749 54895 6783
rect 54895 6749 54904 6783
rect 54852 6740 54904 6749
rect 55312 6740 55364 6792
rect 54576 6715 54628 6724
rect 54576 6681 54585 6715
rect 54585 6681 54619 6715
rect 54619 6681 54628 6715
rect 54576 6672 54628 6681
rect 54944 6604 54996 6656
rect 55128 6604 55180 6656
rect 58348 6740 58400 6792
rect 56048 6672 56100 6724
rect 57336 6672 57388 6724
rect 58716 6740 58768 6792
rect 60004 6808 60056 6860
rect 61660 6808 61712 6860
rect 62488 6808 62540 6860
rect 60464 6740 60516 6792
rect 61752 6740 61804 6792
rect 63592 6876 63644 6928
rect 65432 6876 65484 6928
rect 70952 6876 71004 6928
rect 74080 6876 74132 6928
rect 63684 6851 63736 6860
rect 63684 6817 63693 6851
rect 63693 6817 63727 6851
rect 63727 6817 63736 6851
rect 63684 6808 63736 6817
rect 64144 6740 64196 6792
rect 64420 6740 64472 6792
rect 64604 6783 64656 6792
rect 64604 6749 64613 6783
rect 64613 6749 64647 6783
rect 64647 6749 64656 6783
rect 64604 6740 64656 6749
rect 64788 6740 64840 6792
rect 70676 6808 70728 6860
rect 80520 6851 80572 6860
rect 80520 6817 80529 6851
rect 80529 6817 80563 6851
rect 80563 6817 80572 6851
rect 80520 6808 80572 6817
rect 82912 6851 82964 6860
rect 82912 6817 82921 6851
rect 82921 6817 82955 6851
rect 82955 6817 82964 6851
rect 82912 6808 82964 6817
rect 59360 6672 59412 6724
rect 57704 6604 57756 6656
rect 58072 6647 58124 6656
rect 58072 6613 58081 6647
rect 58081 6613 58115 6647
rect 58115 6613 58124 6647
rect 58072 6604 58124 6613
rect 61476 6672 61528 6724
rect 61660 6672 61712 6724
rect 63316 6672 63368 6724
rect 64880 6715 64932 6724
rect 64880 6681 64889 6715
rect 64889 6681 64923 6715
rect 64923 6681 64932 6715
rect 64880 6672 64932 6681
rect 65064 6672 65116 6724
rect 65156 6672 65208 6724
rect 65432 6740 65484 6792
rect 87328 6740 87380 6792
rect 60924 6604 60976 6656
rect 62764 6647 62816 6656
rect 62764 6613 62773 6647
rect 62773 6613 62807 6647
rect 62807 6613 62816 6647
rect 62764 6604 62816 6613
rect 63408 6604 63460 6656
rect 88892 6672 88944 6724
rect 65524 6604 65576 6656
rect 67088 6604 67140 6656
rect 69756 6604 69808 6656
rect 69848 6604 69900 6656
rect 80244 6604 80296 6656
rect 80336 6604 80388 6656
rect 83188 6604 83240 6656
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 34966 6502 35018 6554
rect 35030 6502 35082 6554
rect 35094 6502 35146 6554
rect 35158 6502 35210 6554
rect 65686 6502 65738 6554
rect 65750 6502 65802 6554
rect 65814 6502 65866 6554
rect 65878 6502 65930 6554
rect 96406 6502 96458 6554
rect 96470 6502 96522 6554
rect 96534 6502 96586 6554
rect 96598 6502 96650 6554
rect 127126 6502 127178 6554
rect 127190 6502 127242 6554
rect 127254 6502 127306 6554
rect 127318 6502 127370 6554
rect 157846 6502 157898 6554
rect 157910 6502 157962 6554
rect 157974 6502 158026 6554
rect 158038 6502 158090 6554
rect 17316 6239 17368 6248
rect 17316 6205 17325 6239
rect 17325 6205 17359 6239
rect 17359 6205 17368 6239
rect 17316 6196 17368 6205
rect 18052 6196 18104 6248
rect 21272 6400 21324 6452
rect 20628 6332 20680 6384
rect 30196 6400 30248 6452
rect 31760 6400 31812 6452
rect 32312 6400 32364 6452
rect 33048 6400 33100 6452
rect 34428 6400 34480 6452
rect 35348 6400 35400 6452
rect 36452 6400 36504 6452
rect 36544 6400 36596 6452
rect 37372 6443 37424 6452
rect 30380 6332 30432 6384
rect 31208 6332 31260 6384
rect 37372 6409 37381 6443
rect 37381 6409 37415 6443
rect 37415 6409 37424 6443
rect 37372 6400 37424 6409
rect 40592 6400 40644 6452
rect 42524 6443 42576 6452
rect 42524 6409 42533 6443
rect 42533 6409 42567 6443
rect 42567 6409 42576 6443
rect 42524 6400 42576 6409
rect 21180 6264 21232 6316
rect 19156 6239 19208 6248
rect 19156 6205 19165 6239
rect 19165 6205 19199 6239
rect 19199 6205 19208 6239
rect 19156 6196 19208 6205
rect 20720 6196 20772 6248
rect 20996 6239 21048 6248
rect 20996 6205 21005 6239
rect 21005 6205 21039 6239
rect 21039 6205 21048 6239
rect 20996 6196 21048 6205
rect 18788 6128 18840 6180
rect 23848 6196 23900 6248
rect 25044 6196 25096 6248
rect 27804 6239 27856 6248
rect 27804 6205 27813 6239
rect 27813 6205 27847 6239
rect 27847 6205 27856 6239
rect 27804 6196 27856 6205
rect 32680 6264 32732 6316
rect 35532 6307 35584 6316
rect 28908 6196 28960 6248
rect 31024 6196 31076 6248
rect 35532 6273 35541 6307
rect 35541 6273 35575 6307
rect 35575 6273 35584 6307
rect 35532 6264 35584 6273
rect 36176 6307 36228 6316
rect 36176 6273 36185 6307
rect 36185 6273 36219 6307
rect 36219 6273 36228 6307
rect 36176 6264 36228 6273
rect 37556 6332 37608 6384
rect 36912 6264 36964 6316
rect 37832 6264 37884 6316
rect 38292 6264 38344 6316
rect 40868 6264 40920 6316
rect 33140 6196 33192 6248
rect 29000 6128 29052 6180
rect 16580 6060 16632 6112
rect 18512 6060 18564 6112
rect 18604 6060 18656 6112
rect 19340 6060 19392 6112
rect 20444 6060 20496 6112
rect 21548 6103 21600 6112
rect 21548 6069 21557 6103
rect 21557 6069 21591 6103
rect 21591 6069 21600 6103
rect 21548 6060 21600 6069
rect 21824 6060 21876 6112
rect 26608 6060 26660 6112
rect 28540 6060 28592 6112
rect 30564 6128 30616 6180
rect 31208 6128 31260 6180
rect 35624 6196 35676 6248
rect 36452 6239 36504 6248
rect 36452 6205 36461 6239
rect 36461 6205 36495 6239
rect 36495 6205 36504 6239
rect 36452 6196 36504 6205
rect 33324 6128 33376 6180
rect 33784 6128 33836 6180
rect 34428 6060 34480 6112
rect 35348 6103 35400 6112
rect 35348 6069 35357 6103
rect 35357 6069 35391 6103
rect 35391 6069 35400 6103
rect 35348 6060 35400 6069
rect 38200 6128 38252 6180
rect 38752 6171 38804 6180
rect 38752 6137 38761 6171
rect 38761 6137 38795 6171
rect 38795 6137 38804 6171
rect 38752 6128 38804 6137
rect 35992 6060 36044 6112
rect 37832 6060 37884 6112
rect 39948 6128 40000 6180
rect 42064 6196 42116 6248
rect 45008 6400 45060 6452
rect 46204 6400 46256 6452
rect 43812 6264 43864 6316
rect 44088 6264 44140 6316
rect 46480 6400 46532 6452
rect 46664 6400 46716 6452
rect 47216 6375 47268 6384
rect 47216 6341 47225 6375
rect 47225 6341 47259 6375
rect 47259 6341 47268 6375
rect 47216 6332 47268 6341
rect 47400 6400 47452 6452
rect 48964 6400 49016 6452
rect 49056 6400 49108 6452
rect 57980 6443 58032 6452
rect 47584 6332 47636 6384
rect 48780 6332 48832 6384
rect 51632 6332 51684 6384
rect 52828 6332 52880 6384
rect 54760 6332 54812 6384
rect 55312 6332 55364 6384
rect 56048 6332 56100 6384
rect 57980 6409 57989 6443
rect 57989 6409 58023 6443
rect 58023 6409 58032 6443
rect 57980 6400 58032 6409
rect 61016 6400 61068 6452
rect 61844 6400 61896 6452
rect 62396 6400 62448 6452
rect 62672 6400 62724 6452
rect 63132 6400 63184 6452
rect 62948 6375 63000 6384
rect 46112 6264 46164 6316
rect 46664 6307 46716 6316
rect 46664 6273 46673 6307
rect 46673 6273 46707 6307
rect 46707 6273 46716 6307
rect 46664 6264 46716 6273
rect 46848 6307 46900 6316
rect 46848 6273 46866 6307
rect 46866 6273 46900 6307
rect 46848 6264 46900 6273
rect 47860 6307 47912 6316
rect 47860 6273 47869 6307
rect 47869 6273 47903 6307
rect 47903 6273 47912 6307
rect 47860 6264 47912 6273
rect 48596 6264 48648 6316
rect 41420 6128 41472 6180
rect 41696 6128 41748 6180
rect 44640 6239 44692 6248
rect 44640 6205 44649 6239
rect 44649 6205 44683 6239
rect 44683 6205 44692 6239
rect 44916 6239 44968 6248
rect 44640 6196 44692 6205
rect 44916 6205 44925 6239
rect 44925 6205 44959 6239
rect 44959 6205 44968 6239
rect 44916 6196 44968 6205
rect 46940 6239 46992 6248
rect 46940 6205 46949 6239
rect 46949 6205 46983 6239
rect 46983 6205 46992 6239
rect 46940 6196 46992 6205
rect 47676 6239 47728 6248
rect 47676 6205 47685 6239
rect 47685 6205 47719 6239
rect 47719 6205 47728 6239
rect 47676 6196 47728 6205
rect 48780 6239 48832 6248
rect 48780 6205 48789 6239
rect 48789 6205 48823 6239
rect 48823 6205 48832 6239
rect 48780 6196 48832 6205
rect 49792 6264 49844 6316
rect 49240 6196 49292 6248
rect 49424 6196 49476 6248
rect 50068 6196 50120 6248
rect 51080 6264 51132 6316
rect 52276 6264 52328 6316
rect 55680 6264 55732 6316
rect 54484 6196 54536 6248
rect 56692 6264 56744 6316
rect 62948 6341 62957 6375
rect 62957 6341 62991 6375
rect 62991 6341 63000 6375
rect 62948 6332 63000 6341
rect 64512 6375 64564 6384
rect 64512 6341 64521 6375
rect 64521 6341 64555 6375
rect 64555 6341 64564 6375
rect 64512 6332 64564 6341
rect 57244 6264 57296 6316
rect 57336 6307 57388 6316
rect 57336 6273 57345 6307
rect 57345 6273 57379 6307
rect 57379 6273 57388 6307
rect 59268 6307 59320 6316
rect 57336 6264 57388 6273
rect 59268 6273 59277 6307
rect 59277 6273 59311 6307
rect 59311 6273 59320 6307
rect 59268 6264 59320 6273
rect 60004 6264 60056 6316
rect 60648 6264 60700 6316
rect 62212 6264 62264 6316
rect 63408 6307 63460 6316
rect 39304 6060 39356 6112
rect 42432 6060 42484 6112
rect 43720 6060 43772 6112
rect 47860 6128 47912 6180
rect 48688 6128 48740 6180
rect 48964 6171 49016 6180
rect 48964 6137 48973 6171
rect 48973 6137 49007 6171
rect 49007 6137 49016 6171
rect 48964 6128 49016 6137
rect 53840 6128 53892 6180
rect 54576 6128 54628 6180
rect 55496 6128 55548 6180
rect 56232 6128 56284 6180
rect 57060 6239 57112 6248
rect 57060 6205 57069 6239
rect 57069 6205 57103 6239
rect 57103 6205 57112 6239
rect 57060 6196 57112 6205
rect 58164 6196 58216 6248
rect 59360 6196 59412 6248
rect 59636 6196 59688 6248
rect 60326 6239 60378 6248
rect 60326 6205 60335 6239
rect 60335 6205 60369 6239
rect 60369 6205 60378 6239
rect 61752 6239 61804 6248
rect 60326 6196 60378 6205
rect 61752 6205 61761 6239
rect 61761 6205 61795 6239
rect 61795 6205 61804 6239
rect 61752 6196 61804 6205
rect 62672 6239 62724 6248
rect 62672 6205 62681 6239
rect 62681 6205 62715 6239
rect 62715 6205 62724 6239
rect 62672 6196 62724 6205
rect 63408 6273 63417 6307
rect 63417 6273 63451 6307
rect 63451 6273 63460 6307
rect 63408 6264 63460 6273
rect 64420 6307 64472 6316
rect 64420 6273 64429 6307
rect 64429 6273 64463 6307
rect 64463 6273 64472 6307
rect 64420 6264 64472 6273
rect 57888 6128 57940 6180
rect 59268 6128 59320 6180
rect 64052 6196 64104 6248
rect 65800 6264 65852 6316
rect 69112 6332 69164 6384
rect 75092 6332 75144 6384
rect 75552 6400 75604 6452
rect 80612 6332 80664 6384
rect 69572 6264 69624 6316
rect 69756 6264 69808 6316
rect 65432 6239 65484 6248
rect 65432 6205 65441 6239
rect 65441 6205 65475 6239
rect 65475 6205 65484 6239
rect 65432 6196 65484 6205
rect 65984 6196 66036 6248
rect 66996 6239 67048 6248
rect 64604 6128 64656 6180
rect 66996 6205 67005 6239
rect 67005 6205 67039 6239
rect 67039 6205 67048 6239
rect 66996 6196 67048 6205
rect 68100 6239 68152 6248
rect 68100 6205 68109 6239
rect 68109 6205 68143 6239
rect 68143 6205 68152 6239
rect 68100 6196 68152 6205
rect 70308 6239 70360 6248
rect 70308 6205 70317 6239
rect 70317 6205 70351 6239
rect 70351 6205 70360 6239
rect 70308 6196 70360 6205
rect 71320 6239 71372 6248
rect 71320 6205 71329 6239
rect 71329 6205 71363 6239
rect 71363 6205 71372 6239
rect 71320 6196 71372 6205
rect 79140 6264 79192 6316
rect 85304 6264 85356 6316
rect 77208 6239 77260 6248
rect 77208 6205 77217 6239
rect 77217 6205 77251 6239
rect 77251 6205 77260 6239
rect 77208 6196 77260 6205
rect 78312 6239 78364 6248
rect 78312 6205 78321 6239
rect 78321 6205 78355 6239
rect 78355 6205 78364 6239
rect 78312 6196 78364 6205
rect 80060 6196 80112 6248
rect 80796 6196 80848 6248
rect 81624 6196 81676 6248
rect 81992 6196 82044 6248
rect 83096 6196 83148 6248
rect 83832 6196 83884 6248
rect 84844 6196 84896 6248
rect 89812 6196 89864 6248
rect 88708 6128 88760 6180
rect 44456 6060 44508 6112
rect 46572 6060 46624 6112
rect 46940 6060 46992 6112
rect 49792 6103 49844 6112
rect 49792 6069 49801 6103
rect 49801 6069 49835 6103
rect 49835 6069 49844 6103
rect 49792 6060 49844 6069
rect 50988 6060 51040 6112
rect 53104 6060 53156 6112
rect 54024 6103 54076 6112
rect 54024 6069 54033 6103
rect 54033 6069 54067 6103
rect 54067 6069 54076 6103
rect 54024 6060 54076 6069
rect 54208 6060 54260 6112
rect 61568 6060 61620 6112
rect 63408 6060 63460 6112
rect 63592 6060 63644 6112
rect 65248 6060 65300 6112
rect 65432 6060 65484 6112
rect 66812 6103 66864 6112
rect 66812 6069 66821 6103
rect 66821 6069 66855 6103
rect 66855 6069 66864 6103
rect 66812 6060 66864 6069
rect 67916 6103 67968 6112
rect 67916 6069 67925 6103
rect 67925 6069 67959 6103
rect 67959 6069 67968 6103
rect 67916 6060 67968 6069
rect 69020 6060 69072 6112
rect 71136 6103 71188 6112
rect 71136 6069 71145 6103
rect 71145 6069 71179 6103
rect 71179 6069 71188 6103
rect 71136 6060 71188 6069
rect 73620 6060 73672 6112
rect 77392 6103 77444 6112
rect 77392 6069 77401 6103
rect 77401 6069 77435 6103
rect 77435 6069 77444 6103
rect 77392 6060 77444 6069
rect 78588 6060 78640 6112
rect 80428 6103 80480 6112
rect 80428 6069 80437 6103
rect 80437 6069 80471 6103
rect 80471 6069 80480 6103
rect 80428 6060 80480 6069
rect 82084 6060 82136 6112
rect 82820 6103 82872 6112
rect 82820 6069 82829 6103
rect 82829 6069 82863 6103
rect 82863 6069 82872 6103
rect 82820 6060 82872 6069
rect 84016 6060 84068 6112
rect 19606 5958 19658 6010
rect 19670 5958 19722 6010
rect 19734 5958 19786 6010
rect 19798 5958 19850 6010
rect 50326 5958 50378 6010
rect 50390 5958 50442 6010
rect 50454 5958 50506 6010
rect 50518 5958 50570 6010
rect 81046 5958 81098 6010
rect 81110 5958 81162 6010
rect 81174 5958 81226 6010
rect 81238 5958 81290 6010
rect 111766 5958 111818 6010
rect 111830 5958 111882 6010
rect 111894 5958 111946 6010
rect 111958 5958 112010 6010
rect 142486 5958 142538 6010
rect 142550 5958 142602 6010
rect 142614 5958 142666 6010
rect 142678 5958 142730 6010
rect 173206 5958 173258 6010
rect 173270 5958 173322 6010
rect 173334 5958 173386 6010
rect 173398 5958 173450 6010
rect 15292 5856 15344 5908
rect 17408 5856 17460 5908
rect 18696 5856 18748 5908
rect 31576 5856 31628 5908
rect 31944 5856 31996 5908
rect 22100 5788 22152 5840
rect 23480 5788 23532 5840
rect 26332 5788 26384 5840
rect 27436 5788 27488 5840
rect 17316 5720 17368 5772
rect 20720 5720 20772 5772
rect 22284 5720 22336 5772
rect 17316 5516 17368 5568
rect 19156 5652 19208 5704
rect 20628 5695 20680 5704
rect 20628 5661 20637 5695
rect 20637 5661 20671 5695
rect 20671 5661 20680 5695
rect 20628 5652 20680 5661
rect 21640 5652 21692 5704
rect 23848 5720 23900 5772
rect 27804 5720 27856 5772
rect 29276 5720 29328 5772
rect 32036 5788 32088 5840
rect 33692 5856 33744 5908
rect 40500 5856 40552 5908
rect 43536 5856 43588 5908
rect 45836 5856 45888 5908
rect 46388 5856 46440 5908
rect 47216 5856 47268 5908
rect 47400 5856 47452 5908
rect 47492 5856 47544 5908
rect 49424 5856 49476 5908
rect 55036 5899 55088 5908
rect 31576 5652 31628 5704
rect 31852 5652 31904 5704
rect 18512 5516 18564 5568
rect 21640 5516 21692 5568
rect 22008 5559 22060 5568
rect 22008 5525 22017 5559
rect 22017 5525 22051 5559
rect 22051 5525 22060 5559
rect 22008 5516 22060 5525
rect 24216 5559 24268 5568
rect 24216 5525 24225 5559
rect 24225 5525 24259 5559
rect 24259 5525 24268 5559
rect 26608 5559 26660 5568
rect 24216 5516 24268 5525
rect 26608 5525 26617 5559
rect 26617 5525 26651 5559
rect 26651 5525 26660 5559
rect 26608 5516 26660 5525
rect 27804 5516 27856 5568
rect 27988 5516 28040 5568
rect 28724 5584 28776 5636
rect 33876 5720 33928 5772
rect 35440 5720 35492 5772
rect 36268 5720 36320 5772
rect 37188 5788 37240 5840
rect 41236 5788 41288 5840
rect 45928 5788 45980 5840
rect 38108 5720 38160 5772
rect 39488 5720 39540 5772
rect 30656 5516 30708 5568
rect 32036 5516 32088 5568
rect 32680 5516 32732 5568
rect 33692 5559 33744 5568
rect 33692 5525 33701 5559
rect 33701 5525 33735 5559
rect 33735 5525 33744 5559
rect 33692 5516 33744 5525
rect 34060 5584 34112 5636
rect 37556 5652 37608 5704
rect 43812 5720 43864 5772
rect 41880 5695 41932 5704
rect 41880 5661 41889 5695
rect 41889 5661 41923 5695
rect 41923 5661 41932 5695
rect 41880 5652 41932 5661
rect 43444 5652 43496 5704
rect 35440 5516 35492 5568
rect 36544 5516 36596 5568
rect 41788 5584 41840 5636
rect 43260 5627 43312 5636
rect 43260 5593 43269 5627
rect 43269 5593 43303 5627
rect 43303 5593 43312 5627
rect 43260 5584 43312 5593
rect 38660 5559 38712 5568
rect 38660 5525 38669 5559
rect 38669 5525 38703 5559
rect 38703 5525 38712 5559
rect 38660 5516 38712 5525
rect 41144 5516 41196 5568
rect 42616 5516 42668 5568
rect 42800 5516 42852 5568
rect 46020 5584 46072 5636
rect 45008 5516 45060 5568
rect 49516 5788 49568 5840
rect 46848 5763 46900 5772
rect 46848 5729 46857 5763
rect 46857 5729 46891 5763
rect 46891 5729 46900 5763
rect 47124 5763 47176 5772
rect 46848 5720 46900 5729
rect 47124 5729 47133 5763
rect 47133 5729 47167 5763
rect 47167 5729 47176 5763
rect 47124 5720 47176 5729
rect 48044 5763 48096 5772
rect 46664 5652 46716 5704
rect 48044 5729 48053 5763
rect 48053 5729 48087 5763
rect 48087 5729 48096 5763
rect 48044 5720 48096 5729
rect 49056 5720 49108 5772
rect 52092 5763 52144 5772
rect 52092 5729 52101 5763
rect 52101 5729 52135 5763
rect 52135 5729 52144 5763
rect 52092 5720 52144 5729
rect 53196 5763 53248 5772
rect 53196 5729 53205 5763
rect 53205 5729 53239 5763
rect 53239 5729 53248 5763
rect 53196 5720 53248 5729
rect 55036 5865 55045 5899
rect 55045 5865 55079 5899
rect 55079 5865 55088 5899
rect 55036 5856 55088 5865
rect 56692 5856 56744 5908
rect 54300 5720 54352 5772
rect 55680 5763 55732 5772
rect 55680 5729 55689 5763
rect 55689 5729 55723 5763
rect 55723 5729 55732 5763
rect 55680 5720 55732 5729
rect 47400 5627 47452 5636
rect 47400 5593 47409 5627
rect 47409 5593 47443 5627
rect 47443 5593 47452 5627
rect 47400 5584 47452 5593
rect 47492 5584 47544 5636
rect 52184 5652 52236 5704
rect 53840 5695 53892 5704
rect 53840 5661 53849 5695
rect 53849 5661 53883 5695
rect 53883 5661 53892 5695
rect 53840 5652 53892 5661
rect 54760 5652 54812 5704
rect 47308 5516 47360 5568
rect 47860 5516 47912 5568
rect 48044 5516 48096 5568
rect 49976 5516 50028 5568
rect 52828 5516 52880 5568
rect 52920 5516 52972 5568
rect 56048 5516 56100 5568
rect 58532 5856 58584 5908
rect 59544 5856 59596 5908
rect 59268 5788 59320 5840
rect 63132 5856 63184 5908
rect 58532 5763 58584 5772
rect 58532 5729 58566 5763
rect 58566 5729 58584 5763
rect 58716 5763 58768 5772
rect 58532 5720 58584 5729
rect 58716 5729 58725 5763
rect 58725 5729 58759 5763
rect 58759 5729 58768 5763
rect 58716 5720 58768 5729
rect 59452 5720 59504 5772
rect 60648 5763 60700 5772
rect 60648 5729 60665 5763
rect 60665 5729 60699 5763
rect 60699 5729 60700 5763
rect 60648 5720 60700 5729
rect 62120 5720 62172 5772
rect 62948 5720 63000 5772
rect 63408 5720 63460 5772
rect 64236 5763 64288 5772
rect 64236 5729 64254 5763
rect 64254 5729 64288 5763
rect 64236 5720 64288 5729
rect 57612 5652 57664 5704
rect 58256 5652 58308 5704
rect 62304 5652 62356 5704
rect 64052 5695 64104 5704
rect 64052 5661 64061 5695
rect 64061 5661 64095 5695
rect 64095 5661 64104 5695
rect 64052 5652 64104 5661
rect 64328 5695 64380 5704
rect 64328 5661 64337 5695
rect 64337 5661 64371 5695
rect 64371 5661 64380 5695
rect 64328 5652 64380 5661
rect 65248 5856 65300 5908
rect 68008 5856 68060 5908
rect 68928 5856 68980 5908
rect 73712 5856 73764 5908
rect 75092 5856 75144 5908
rect 77760 5856 77812 5908
rect 82820 5856 82872 5908
rect 89076 5856 89128 5908
rect 65524 5788 65576 5840
rect 72056 5788 72108 5840
rect 65340 5720 65392 5772
rect 68928 5720 68980 5772
rect 69664 5720 69716 5772
rect 72608 5763 72660 5772
rect 72608 5729 72617 5763
rect 72617 5729 72651 5763
rect 72651 5729 72660 5763
rect 73252 5763 73304 5772
rect 72608 5720 72660 5729
rect 73252 5729 73261 5763
rect 73261 5729 73295 5763
rect 73295 5729 73304 5763
rect 73252 5720 73304 5729
rect 74080 5763 74132 5772
rect 74080 5729 74089 5763
rect 74089 5729 74123 5763
rect 74123 5729 74132 5763
rect 74080 5720 74132 5729
rect 74632 5720 74684 5772
rect 77576 5720 77628 5772
rect 77668 5720 77720 5772
rect 78680 5720 78732 5772
rect 79416 5720 79468 5772
rect 58164 5627 58216 5636
rect 58164 5593 58173 5627
rect 58173 5593 58207 5627
rect 58207 5593 58216 5627
rect 58164 5584 58216 5593
rect 64604 5627 64656 5636
rect 59452 5516 59504 5568
rect 59912 5516 59964 5568
rect 63592 5516 63644 5568
rect 64604 5593 64613 5627
rect 64613 5593 64647 5627
rect 64647 5593 64656 5627
rect 64604 5584 64656 5593
rect 64880 5584 64932 5636
rect 65248 5695 65300 5704
rect 65248 5661 65257 5695
rect 65257 5661 65291 5695
rect 65291 5661 65300 5695
rect 65248 5652 65300 5661
rect 68192 5652 68244 5704
rect 70216 5652 70268 5704
rect 79140 5652 79192 5704
rect 79416 5584 79468 5636
rect 79876 5788 79928 5840
rect 79600 5720 79652 5772
rect 79784 5720 79836 5772
rect 81716 5763 81768 5772
rect 81716 5729 81725 5763
rect 81725 5729 81759 5763
rect 81759 5729 81768 5763
rect 81716 5720 81768 5729
rect 82820 5720 82872 5772
rect 84476 5763 84528 5772
rect 84476 5729 84485 5763
rect 84485 5729 84519 5763
rect 84519 5729 84528 5763
rect 84476 5720 84528 5729
rect 84936 5720 84988 5772
rect 86040 5763 86092 5772
rect 86040 5729 86049 5763
rect 86049 5729 86083 5763
rect 86083 5729 86092 5763
rect 86040 5720 86092 5729
rect 178684 5720 178736 5772
rect 79600 5584 79652 5636
rect 64788 5516 64840 5568
rect 65248 5516 65300 5568
rect 67824 5516 67876 5568
rect 73804 5516 73856 5568
rect 75184 5516 75236 5568
rect 79968 5516 80020 5568
rect 80244 5584 80296 5636
rect 89996 5652 90048 5704
rect 82176 5584 82228 5636
rect 80888 5516 80940 5568
rect 82452 5516 82504 5568
rect 83556 5516 83608 5568
rect 85120 5516 85172 5568
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 34966 5414 35018 5466
rect 35030 5414 35082 5466
rect 35094 5414 35146 5466
rect 35158 5414 35210 5466
rect 65686 5414 65738 5466
rect 65750 5414 65802 5466
rect 65814 5414 65866 5466
rect 65878 5414 65930 5466
rect 96406 5414 96458 5466
rect 96470 5414 96522 5466
rect 96534 5414 96586 5466
rect 96598 5414 96650 5466
rect 127126 5414 127178 5466
rect 127190 5414 127242 5466
rect 127254 5414 127306 5466
rect 127318 5414 127370 5466
rect 157846 5414 157898 5466
rect 157910 5414 157962 5466
rect 157974 5414 158026 5466
rect 158038 5414 158090 5466
rect 1952 5312 2004 5364
rect 23756 5312 23808 5364
rect 18696 5287 18748 5296
rect 18696 5253 18705 5287
rect 18705 5253 18739 5287
rect 18739 5253 18748 5287
rect 18696 5244 18748 5253
rect 20536 5287 20588 5296
rect 20536 5253 20545 5287
rect 20545 5253 20579 5287
rect 20579 5253 20588 5287
rect 20536 5244 20588 5253
rect 17316 5219 17368 5228
rect 17316 5185 17325 5219
rect 17325 5185 17359 5219
rect 17359 5185 17368 5219
rect 17316 5176 17368 5185
rect 19156 5219 19208 5228
rect 19156 5185 19165 5219
rect 19165 5185 19199 5219
rect 19199 5185 19208 5219
rect 19156 5176 19208 5185
rect 28816 5312 28868 5364
rect 28172 5176 28224 5228
rect 30564 5312 30616 5364
rect 30932 5312 30984 5364
rect 31576 5244 31628 5296
rect 29276 5219 29328 5228
rect 29276 5185 29285 5219
rect 29285 5185 29319 5219
rect 29319 5185 29328 5219
rect 29276 5176 29328 5185
rect 21088 5108 21140 5160
rect 24952 5108 25004 5160
rect 25412 5108 25464 5160
rect 34244 5312 34296 5364
rect 34336 5312 34388 5364
rect 32036 5176 32088 5228
rect 21548 5040 21600 5092
rect 27988 5040 28040 5092
rect 15660 4972 15712 5024
rect 20536 4972 20588 5024
rect 28356 4972 28408 5024
rect 33140 5040 33192 5092
rect 34796 5244 34848 5296
rect 35992 5312 36044 5364
rect 36084 5312 36136 5364
rect 37280 5244 37332 5296
rect 38292 5312 38344 5364
rect 39856 5244 39908 5296
rect 41512 5355 41564 5364
rect 41512 5321 41521 5355
rect 41521 5321 41555 5355
rect 41555 5321 41564 5355
rect 41512 5312 41564 5321
rect 42156 5312 42208 5364
rect 41880 5244 41932 5296
rect 43536 5244 43588 5296
rect 46756 5312 46808 5364
rect 47676 5312 47728 5364
rect 47216 5244 47268 5296
rect 63224 5312 63276 5364
rect 72056 5312 72108 5364
rect 76564 5312 76616 5364
rect 78772 5312 78824 5364
rect 81808 5312 81860 5364
rect 82452 5312 82504 5364
rect 84660 5312 84712 5364
rect 84752 5312 84804 5364
rect 88984 5312 89036 5364
rect 34520 5040 34572 5092
rect 38292 5151 38344 5160
rect 38292 5117 38301 5151
rect 38301 5117 38335 5151
rect 38335 5117 38344 5151
rect 38292 5108 38344 5117
rect 44824 5176 44876 5228
rect 45284 5176 45336 5228
rect 46388 5176 46440 5228
rect 47768 5176 47820 5228
rect 61660 5176 61712 5228
rect 61936 5219 61988 5228
rect 61936 5185 61945 5219
rect 61945 5185 61979 5219
rect 61979 5185 61988 5219
rect 61936 5176 61988 5185
rect 62396 5176 62448 5228
rect 43536 5151 43588 5160
rect 43536 5117 43545 5151
rect 43545 5117 43579 5151
rect 43579 5117 43588 5151
rect 43536 5108 43588 5117
rect 30472 4972 30524 5024
rect 30564 4972 30616 5024
rect 30748 4972 30800 5024
rect 31760 4972 31812 5024
rect 31852 4972 31904 5024
rect 38384 5040 38436 5092
rect 38476 5040 38528 5092
rect 38660 5040 38712 5092
rect 39212 5040 39264 5092
rect 36268 5015 36320 5024
rect 36268 4981 36277 5015
rect 36277 4981 36311 5015
rect 36311 4981 36320 5015
rect 36268 4972 36320 4981
rect 37096 4972 37148 5024
rect 39948 5040 40000 5092
rect 44180 5108 44232 5160
rect 47032 5108 47084 5160
rect 47400 5151 47452 5160
rect 47400 5117 47409 5151
rect 47409 5117 47443 5151
rect 47443 5117 47452 5151
rect 47400 5108 47452 5117
rect 62212 5151 62264 5160
rect 62212 5117 62221 5151
rect 62221 5117 62255 5151
rect 62255 5117 62264 5151
rect 62488 5151 62540 5160
rect 62212 5108 62264 5117
rect 62488 5117 62497 5151
rect 62497 5117 62531 5151
rect 62531 5117 62540 5151
rect 62488 5108 62540 5117
rect 50620 5040 50672 5092
rect 40040 4972 40092 5024
rect 41512 4972 41564 5024
rect 43996 4972 44048 5024
rect 45376 4972 45428 5024
rect 45468 4972 45520 5024
rect 46388 4972 46440 5024
rect 46480 4972 46532 5024
rect 47032 4972 47084 5024
rect 49884 4972 49936 5024
rect 60464 4972 60516 5024
rect 64788 5176 64840 5228
rect 63868 5108 63920 5160
rect 76104 5108 76156 5160
rect 76472 5108 76524 5160
rect 77576 5151 77628 5160
rect 77576 5117 77585 5151
rect 77585 5117 77619 5151
rect 77619 5117 77628 5151
rect 77576 5108 77628 5117
rect 71964 5040 72016 5092
rect 63500 4972 63552 5024
rect 75920 4972 75972 5024
rect 76380 4972 76432 5024
rect 78220 5176 78272 5228
rect 78772 5176 78824 5228
rect 78128 5108 78180 5160
rect 80244 5108 80296 5160
rect 80704 5176 80756 5228
rect 82636 5219 82688 5228
rect 82636 5185 82645 5219
rect 82645 5185 82679 5219
rect 82679 5185 82688 5219
rect 82636 5176 82688 5185
rect 79324 4972 79376 5024
rect 80336 4972 80388 5024
rect 82820 5108 82872 5160
rect 83372 5108 83424 5160
rect 83464 5151 83516 5160
rect 83464 5117 83473 5151
rect 83473 5117 83507 5151
rect 83507 5117 83516 5151
rect 83464 5108 83516 5117
rect 82268 5083 82320 5092
rect 82268 5049 82277 5083
rect 82277 5049 82311 5083
rect 82311 5049 82320 5083
rect 82268 5040 82320 5049
rect 86224 5176 86276 5228
rect 94412 5312 94464 5364
rect 85580 5108 85632 5160
rect 86776 5151 86828 5160
rect 86776 5117 86785 5151
rect 86785 5117 86819 5151
rect 86819 5117 86828 5151
rect 86776 5108 86828 5117
rect 87144 5108 87196 5160
rect 177580 5108 177632 5160
rect 179052 5108 179104 5160
rect 86684 5040 86736 5092
rect 81532 4972 81584 5024
rect 83280 5015 83332 5024
rect 83280 4981 83289 5015
rect 83289 4981 83323 5015
rect 83323 4981 83332 5015
rect 83280 4972 83332 4981
rect 83372 5015 83424 5024
rect 83372 4981 83381 5015
rect 83381 4981 83415 5015
rect 83415 4981 83424 5015
rect 83648 5015 83700 5024
rect 83372 4972 83424 4981
rect 83648 4981 83657 5015
rect 83657 4981 83691 5015
rect 83691 4981 83700 5015
rect 83648 4972 83700 4981
rect 84292 5015 84344 5024
rect 84292 4981 84301 5015
rect 84301 4981 84335 5015
rect 84335 4981 84344 5015
rect 84292 4972 84344 4981
rect 86224 4972 86276 5024
rect 86500 4972 86552 5024
rect 102784 4972 102836 5024
rect 19606 4870 19658 4922
rect 19670 4870 19722 4922
rect 19734 4870 19786 4922
rect 19798 4870 19850 4922
rect 50326 4870 50378 4922
rect 50390 4870 50442 4922
rect 50454 4870 50506 4922
rect 50518 4870 50570 4922
rect 81046 4870 81098 4922
rect 81110 4870 81162 4922
rect 81174 4870 81226 4922
rect 81238 4870 81290 4922
rect 111766 4870 111818 4922
rect 111830 4870 111882 4922
rect 111894 4870 111946 4922
rect 111958 4870 112010 4922
rect 142486 4870 142538 4922
rect 142550 4870 142602 4922
rect 142614 4870 142666 4922
rect 142678 4870 142730 4922
rect 173206 4870 173258 4922
rect 173270 4870 173322 4922
rect 173334 4870 173386 4922
rect 173398 4870 173450 4922
rect 20076 4768 20128 4820
rect 26608 4768 26660 4820
rect 28356 4811 28408 4820
rect 28356 4777 28365 4811
rect 28365 4777 28399 4811
rect 28399 4777 28408 4811
rect 28356 4768 28408 4777
rect 37004 4811 37056 4820
rect 37004 4777 37013 4811
rect 37013 4777 37047 4811
rect 37047 4777 37056 4811
rect 37004 4768 37056 4777
rect 37280 4768 37332 4820
rect 23756 4700 23808 4752
rect 27988 4700 28040 4752
rect 36636 4700 36688 4752
rect 11796 4675 11848 4684
rect 11796 4641 11805 4675
rect 11805 4641 11839 4675
rect 11839 4641 11848 4675
rect 11796 4632 11848 4641
rect 21548 4632 21600 4684
rect 27896 4632 27948 4684
rect 28080 4632 28132 4684
rect 28908 4632 28960 4684
rect 34244 4632 34296 4684
rect 14280 4496 14332 4548
rect 21916 4496 21968 4548
rect 28172 4564 28224 4616
rect 30472 4564 30524 4616
rect 31668 4564 31720 4616
rect 32404 4607 32456 4616
rect 32404 4573 32413 4607
rect 32413 4573 32447 4607
rect 32447 4573 32456 4607
rect 32404 4564 32456 4573
rect 33784 4564 33836 4616
rect 30748 4496 30800 4548
rect 33140 4496 33192 4548
rect 33692 4496 33744 4548
rect 36912 4564 36964 4616
rect 36084 4496 36136 4548
rect 37188 4496 37240 4548
rect 38292 4632 38344 4684
rect 38660 4768 38712 4820
rect 41972 4768 42024 4820
rect 45468 4768 45520 4820
rect 40224 4700 40276 4752
rect 48136 4768 48188 4820
rect 73896 4768 73948 4820
rect 81440 4768 81492 4820
rect 84108 4768 84160 4820
rect 102784 4811 102836 4820
rect 102784 4777 102793 4811
rect 102793 4777 102827 4811
rect 102827 4777 102836 4811
rect 102784 4768 102836 4777
rect 46112 4700 46164 4752
rect 52184 4700 52236 4752
rect 53932 4700 53984 4752
rect 39764 4632 39816 4684
rect 43536 4632 43588 4684
rect 45376 4632 45428 4684
rect 46296 4632 46348 4684
rect 46940 4632 46992 4684
rect 47032 4632 47084 4684
rect 49608 4632 49660 4684
rect 70584 4675 70636 4684
rect 70584 4641 70593 4675
rect 70593 4641 70627 4675
rect 70627 4641 70636 4675
rect 70584 4632 70636 4641
rect 71780 4632 71832 4684
rect 72792 4632 72844 4684
rect 75000 4632 75052 4684
rect 75368 4632 75420 4684
rect 75920 4632 75972 4684
rect 76656 4632 76708 4684
rect 77576 4700 77628 4752
rect 79232 4700 79284 4752
rect 80244 4743 80296 4752
rect 80244 4709 80253 4743
rect 80253 4709 80287 4743
rect 80287 4709 80296 4743
rect 80244 4700 80296 4709
rect 80888 4700 80940 4752
rect 83648 4700 83700 4752
rect 98092 4700 98144 4752
rect 82820 4632 82872 4684
rect 45284 4564 45336 4616
rect 45744 4564 45796 4616
rect 46020 4564 46072 4616
rect 59636 4564 59688 4616
rect 35900 4428 35952 4480
rect 36636 4428 36688 4480
rect 39212 4428 39264 4480
rect 39764 4428 39816 4480
rect 62120 4496 62172 4548
rect 68008 4496 68060 4548
rect 75460 4496 75512 4548
rect 80704 4496 80756 4548
rect 81348 4496 81400 4548
rect 82544 4564 82596 4616
rect 83004 4564 83056 4616
rect 83924 4632 83976 4684
rect 84016 4632 84068 4684
rect 83648 4564 83700 4616
rect 85488 4539 85540 4548
rect 85488 4505 85497 4539
rect 85497 4505 85531 4539
rect 85531 4505 85540 4539
rect 85488 4496 85540 4505
rect 87512 4632 87564 4684
rect 88340 4632 88392 4684
rect 89352 4632 89404 4684
rect 93768 4675 93820 4684
rect 93768 4641 93777 4675
rect 93777 4641 93811 4675
rect 93811 4641 93820 4675
rect 93768 4632 93820 4641
rect 102600 4675 102652 4684
rect 102600 4641 102609 4675
rect 102609 4641 102643 4675
rect 102643 4641 102652 4675
rect 102600 4632 102652 4641
rect 175372 4675 175424 4684
rect 175372 4641 175381 4675
rect 175381 4641 175415 4675
rect 175415 4641 175424 4675
rect 175372 4632 175424 4641
rect 86500 4564 86552 4616
rect 176660 4632 176712 4684
rect 177948 4675 178000 4684
rect 177948 4641 177957 4675
rect 177957 4641 177991 4675
rect 177991 4641 178000 4675
rect 177948 4632 178000 4641
rect 88156 4496 88208 4548
rect 88432 4496 88484 4548
rect 88984 4539 89036 4548
rect 88984 4505 88993 4539
rect 88993 4505 89027 4539
rect 89027 4505 89036 4539
rect 88984 4496 89036 4505
rect 179788 4564 179840 4616
rect 48320 4428 48372 4480
rect 48596 4428 48648 4480
rect 74724 4428 74776 4480
rect 75644 4428 75696 4480
rect 76748 4471 76800 4480
rect 76748 4437 76757 4471
rect 76757 4437 76791 4471
rect 76791 4437 76800 4471
rect 76748 4428 76800 4437
rect 77944 4428 77996 4480
rect 80152 4428 80204 4480
rect 80888 4428 80940 4480
rect 81716 4428 81768 4480
rect 82268 4428 82320 4480
rect 84660 4428 84712 4480
rect 86132 4471 86184 4480
rect 86132 4437 86141 4471
rect 86141 4437 86175 4471
rect 86175 4437 86184 4471
rect 86132 4428 86184 4437
rect 86960 4428 87012 4480
rect 89168 4428 89220 4480
rect 94504 4428 94556 4480
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 34966 4326 35018 4378
rect 35030 4326 35082 4378
rect 35094 4326 35146 4378
rect 35158 4326 35210 4378
rect 65686 4326 65738 4378
rect 65750 4326 65802 4378
rect 65814 4326 65866 4378
rect 65878 4326 65930 4378
rect 96406 4326 96458 4378
rect 96470 4326 96522 4378
rect 96534 4326 96586 4378
rect 96598 4326 96650 4378
rect 127126 4326 127178 4378
rect 127190 4326 127242 4378
rect 127254 4326 127306 4378
rect 127318 4326 127370 4378
rect 157846 4326 157898 4378
rect 157910 4326 157962 4378
rect 157974 4326 158026 4378
rect 158038 4326 158090 4378
rect 5816 4224 5868 4276
rect 32312 4224 32364 4276
rect 32404 4224 32456 4276
rect 46112 4224 46164 4276
rect 51816 4224 51868 4276
rect 78036 4224 78088 4276
rect 78404 4224 78456 4276
rect 78496 4224 78548 4276
rect 80888 4224 80940 4276
rect 82452 4224 82504 4276
rect 83924 4224 83976 4276
rect 84016 4224 84068 4276
rect 85212 4224 85264 4276
rect 19340 4156 19392 4208
rect 21916 4156 21968 4208
rect 34060 4156 34112 4208
rect 3148 4088 3200 4140
rect 12348 4088 12400 4140
rect 1124 4020 1176 4072
rect 1860 4020 1912 4072
rect 10968 4020 11020 4072
rect 12716 4020 12768 4072
rect 13636 4063 13688 4072
rect 13636 4029 13645 4063
rect 13645 4029 13679 4063
rect 13679 4029 13688 4063
rect 13636 4020 13688 4029
rect 14832 4088 14884 4140
rect 21824 4088 21876 4140
rect 15660 4020 15712 4072
rect 15844 4063 15896 4072
rect 15844 4029 15853 4063
rect 15853 4029 15887 4063
rect 15887 4029 15896 4063
rect 15844 4020 15896 4029
rect 16212 4020 16264 4072
rect 20076 4020 20128 4072
rect 20260 4063 20312 4072
rect 20260 4029 20269 4063
rect 20269 4029 20303 4063
rect 20303 4029 20312 4063
rect 20260 4020 20312 4029
rect 24952 4088 25004 4140
rect 25504 4088 25556 4140
rect 35992 4131 36044 4140
rect 12072 3952 12124 4004
rect 12256 3952 12308 4004
rect 12440 3952 12492 4004
rect 9956 3884 10008 3936
rect 10048 3884 10100 3936
rect 13728 3952 13780 4004
rect 22376 4020 22428 4072
rect 31944 4020 31996 4072
rect 35992 4097 36001 4131
rect 36001 4097 36035 4131
rect 36035 4097 36044 4131
rect 35992 4088 36044 4097
rect 38292 4131 38344 4140
rect 38292 4097 38301 4131
rect 38301 4097 38335 4131
rect 38335 4097 38344 4131
rect 38292 4088 38344 4097
rect 39580 4088 39632 4140
rect 39764 4156 39816 4208
rect 51632 4199 51684 4208
rect 40776 4088 40828 4140
rect 40960 4088 41012 4140
rect 43996 4088 44048 4140
rect 51632 4165 51641 4199
rect 51641 4165 51675 4199
rect 51675 4165 51684 4199
rect 51632 4156 51684 4165
rect 56232 4156 56284 4208
rect 36084 4020 36136 4072
rect 12624 3884 12676 3936
rect 18788 3884 18840 3936
rect 18880 3884 18932 3936
rect 22100 3884 22152 3936
rect 22192 3884 22244 3936
rect 34152 3952 34204 4004
rect 27896 3884 27948 3936
rect 38200 4020 38252 4072
rect 42248 4020 42300 4072
rect 45744 4063 45796 4072
rect 45744 4029 45753 4063
rect 45753 4029 45787 4063
rect 45787 4029 45796 4063
rect 45744 4020 45796 4029
rect 71044 4088 71096 4140
rect 73436 4088 73488 4140
rect 56968 4063 57020 4072
rect 56968 4029 56977 4063
rect 56977 4029 57011 4063
rect 57011 4029 57020 4063
rect 56968 4020 57020 4029
rect 66168 4063 66220 4072
rect 66168 4029 66177 4063
rect 66177 4029 66211 4063
rect 66211 4029 66220 4063
rect 66168 4020 66220 4029
rect 67272 4063 67324 4072
rect 67272 4029 67281 4063
rect 67281 4029 67315 4063
rect 67315 4029 67324 4063
rect 67272 4020 67324 4029
rect 68376 4063 68428 4072
rect 68376 4029 68385 4063
rect 68385 4029 68419 4063
rect 68419 4029 68428 4063
rect 68376 4020 68428 4029
rect 69480 4020 69532 4072
rect 70952 4020 71004 4072
rect 71228 4063 71280 4072
rect 71228 4029 71237 4063
rect 71237 4029 71271 4063
rect 71271 4029 71280 4063
rect 71228 4020 71280 4029
rect 72056 4063 72108 4072
rect 72056 4029 72065 4063
rect 72065 4029 72099 4063
rect 72099 4029 72108 4063
rect 72056 4020 72108 4029
rect 73160 4063 73212 4072
rect 73160 4029 73169 4063
rect 73169 4029 73203 4063
rect 73203 4029 73212 4063
rect 73160 4020 73212 4029
rect 73896 4063 73948 4072
rect 73896 4029 73905 4063
rect 73905 4029 73939 4063
rect 73939 4029 73948 4063
rect 73896 4020 73948 4029
rect 74264 4020 74316 4072
rect 76748 4063 76800 4072
rect 37464 3884 37516 3936
rect 38384 3952 38436 4004
rect 40132 3884 40184 3936
rect 49332 3952 49384 4004
rect 70860 3952 70912 4004
rect 71412 3952 71464 4004
rect 76748 4029 76757 4063
rect 76757 4029 76791 4063
rect 76791 4029 76800 4063
rect 76748 4020 76800 4029
rect 77576 4088 77628 4140
rect 78496 4088 78548 4140
rect 80244 4088 80296 4140
rect 80428 4156 80480 4208
rect 82360 4156 82412 4208
rect 81900 4088 81952 4140
rect 78128 4020 78180 4072
rect 79968 4020 80020 4072
rect 80428 4020 80480 4072
rect 80704 4020 80756 4072
rect 78220 3995 78272 4004
rect 48228 3884 48280 3936
rect 70400 3884 70452 3936
rect 71044 3884 71096 3936
rect 71504 3927 71556 3936
rect 71504 3893 71513 3927
rect 71513 3893 71547 3927
rect 71547 3893 71556 3927
rect 71504 3884 71556 3893
rect 75092 3884 75144 3936
rect 76840 3927 76892 3936
rect 76840 3893 76849 3927
rect 76849 3893 76883 3927
rect 76883 3893 76892 3927
rect 76840 3884 76892 3893
rect 78220 3961 78229 3995
rect 78229 3961 78263 3995
rect 78263 3961 78272 3995
rect 78220 3952 78272 3961
rect 79140 3952 79192 4004
rect 77576 3884 77628 3936
rect 79600 3884 79652 3936
rect 80060 3884 80112 3936
rect 80336 3884 80388 3936
rect 84108 4156 84160 4208
rect 84568 4199 84620 4208
rect 84568 4165 84577 4199
rect 84577 4165 84611 4199
rect 84611 4165 84620 4199
rect 84568 4156 84620 4165
rect 85028 4156 85080 4208
rect 86868 4224 86920 4276
rect 87052 4156 87104 4208
rect 83004 4088 83056 4140
rect 80888 3952 80940 4004
rect 83740 4020 83792 4072
rect 81808 3952 81860 4004
rect 82820 3952 82872 4004
rect 87604 4088 87656 4140
rect 88524 4224 88576 4276
rect 88708 4224 88760 4276
rect 89444 4267 89496 4276
rect 89444 4233 89453 4267
rect 89453 4233 89487 4267
rect 89487 4233 89496 4267
rect 89444 4224 89496 4233
rect 89536 4224 89588 4276
rect 109316 4224 109368 4276
rect 90824 4156 90876 4208
rect 84200 4063 84252 4072
rect 84200 4029 84209 4063
rect 84209 4029 84243 4063
rect 84243 4029 84252 4063
rect 84200 4020 84252 4029
rect 83924 3952 83976 4004
rect 84568 3952 84620 4004
rect 85396 3952 85448 4004
rect 86684 4020 86736 4072
rect 86960 4063 87012 4072
rect 86960 4029 86969 4063
rect 86969 4029 87003 4063
rect 87003 4029 87012 4063
rect 86960 4020 87012 4029
rect 87788 4020 87840 4072
rect 81716 3927 81768 3936
rect 81716 3893 81725 3927
rect 81725 3893 81759 3927
rect 81759 3893 81768 3927
rect 81716 3884 81768 3893
rect 81900 3927 81952 3936
rect 81900 3893 81909 3927
rect 81909 3893 81943 3927
rect 81943 3893 81952 3927
rect 81900 3884 81952 3893
rect 85028 3884 85080 3936
rect 85672 3884 85724 3936
rect 86224 3927 86276 3936
rect 86224 3893 86233 3927
rect 86233 3893 86267 3927
rect 86267 3893 86276 3927
rect 86224 3884 86276 3893
rect 86592 3884 86644 3936
rect 86776 3884 86828 3936
rect 88616 3995 88668 4004
rect 88616 3961 88625 3995
rect 88625 3961 88659 3995
rect 88659 3961 88668 3995
rect 88616 3952 88668 3961
rect 89720 4088 89772 4140
rect 91100 4156 91152 4208
rect 92388 4156 92440 4208
rect 91008 4088 91060 4140
rect 94504 4156 94556 4208
rect 109960 4156 110012 4208
rect 94412 4088 94464 4140
rect 90456 4020 90508 4072
rect 91560 4063 91612 4072
rect 91560 4029 91569 4063
rect 91569 4029 91603 4063
rect 91603 4029 91612 4063
rect 91560 4020 91612 4029
rect 91652 4020 91704 4072
rect 92664 4020 92716 4072
rect 93032 4063 93084 4072
rect 93032 4029 93041 4063
rect 93041 4029 93075 4063
rect 93075 4029 93084 4063
rect 93032 4020 93084 4029
rect 94136 4063 94188 4072
rect 94136 4029 94145 4063
rect 94145 4029 94179 4063
rect 94179 4029 94188 4063
rect 94136 4020 94188 4029
rect 94872 4063 94924 4072
rect 94872 4029 94881 4063
rect 94881 4029 94915 4063
rect 94915 4029 94924 4063
rect 94872 4020 94924 4029
rect 95976 4063 96028 4072
rect 95976 4029 95985 4063
rect 95985 4029 96019 4063
rect 96019 4029 96028 4063
rect 95976 4020 96028 4029
rect 98000 4088 98052 4140
rect 102876 4088 102928 4140
rect 97080 4063 97132 4072
rect 97080 4029 97089 4063
rect 97089 4029 97123 4063
rect 97123 4029 97132 4063
rect 97080 4020 97132 4029
rect 98184 4063 98236 4072
rect 98184 4029 98193 4063
rect 98193 4029 98227 4063
rect 98227 4029 98236 4063
rect 98184 4020 98236 4029
rect 99288 4063 99340 4072
rect 99288 4029 99297 4063
rect 99297 4029 99331 4063
rect 99331 4029 99340 4063
rect 99288 4020 99340 4029
rect 100392 4020 100444 4072
rect 101496 4020 101548 4072
rect 102968 4063 103020 4072
rect 102968 4029 102977 4063
rect 102977 4029 103011 4063
rect 103011 4029 103020 4063
rect 102968 4020 103020 4029
rect 91652 3884 91704 3936
rect 91836 3884 91888 3936
rect 93216 3927 93268 3936
rect 93216 3893 93225 3927
rect 93225 3893 93259 3927
rect 93259 3893 93268 3927
rect 93216 3884 93268 3893
rect 95056 3927 95108 3936
rect 95056 3893 95065 3927
rect 95065 3893 95099 3927
rect 95099 3893 95108 3927
rect 95056 3884 95108 3893
rect 97264 3927 97316 3936
rect 97264 3893 97273 3927
rect 97273 3893 97307 3927
rect 97307 3893 97316 3927
rect 97264 3884 97316 3893
rect 98368 3927 98420 3936
rect 98368 3893 98377 3927
rect 98377 3893 98411 3927
rect 98411 3893 98420 3927
rect 98368 3884 98420 3893
rect 101036 3952 101088 4004
rect 103796 4020 103848 4072
rect 104808 4063 104860 4072
rect 104808 4029 104817 4063
rect 104817 4029 104851 4063
rect 104851 4029 104860 4063
rect 104808 4020 104860 4029
rect 105912 4020 105964 4072
rect 107016 4020 107068 4072
rect 111432 4020 111484 4072
rect 112536 4063 112588 4072
rect 112536 4029 112545 4063
rect 112545 4029 112579 4063
rect 112579 4029 112588 4063
rect 112536 4020 112588 4029
rect 113640 4063 113692 4072
rect 113640 4029 113649 4063
rect 113649 4029 113683 4063
rect 113683 4029 113692 4063
rect 113640 4020 113692 4029
rect 114744 4063 114796 4072
rect 114744 4029 114753 4063
rect 114753 4029 114787 4063
rect 114787 4029 114796 4063
rect 114744 4020 114796 4029
rect 115848 4063 115900 4072
rect 115848 4029 115857 4063
rect 115857 4029 115891 4063
rect 115891 4029 115900 4063
rect 115848 4020 115900 4029
rect 116952 4063 117004 4072
rect 116952 4029 116961 4063
rect 116961 4029 116995 4063
rect 116995 4029 117004 4063
rect 116952 4020 117004 4029
rect 118056 4063 118108 4072
rect 118056 4029 118065 4063
rect 118065 4029 118099 4063
rect 118099 4029 118108 4063
rect 118056 4020 118108 4029
rect 119160 4063 119212 4072
rect 119160 4029 119169 4063
rect 119169 4029 119203 4063
rect 119203 4029 119212 4063
rect 119160 4020 119212 4029
rect 120172 4063 120224 4072
rect 120172 4029 120181 4063
rect 120181 4029 120215 4063
rect 120215 4029 120224 4063
rect 120172 4020 120224 4029
rect 121276 4020 121328 4072
rect 122288 4020 122340 4072
rect 123484 4063 123536 4072
rect 123484 4029 123493 4063
rect 123493 4029 123527 4063
rect 123527 4029 123536 4063
rect 123484 4020 123536 4029
rect 124588 4063 124640 4072
rect 124588 4029 124597 4063
rect 124597 4029 124631 4063
rect 124631 4029 124640 4063
rect 124588 4020 124640 4029
rect 125692 4063 125744 4072
rect 125692 4029 125701 4063
rect 125701 4029 125735 4063
rect 125735 4029 125744 4063
rect 125692 4020 125744 4029
rect 126796 4020 126848 4072
rect 127900 4020 127952 4072
rect 131212 4063 131264 4072
rect 131212 4029 131221 4063
rect 131221 4029 131255 4063
rect 131255 4029 131264 4063
rect 131212 4020 131264 4029
rect 133420 4063 133472 4072
rect 133420 4029 133429 4063
rect 133429 4029 133463 4063
rect 133463 4029 133472 4063
rect 133420 4020 133472 4029
rect 134524 4063 134576 4072
rect 134524 4029 134533 4063
rect 134533 4029 134567 4063
rect 134567 4029 134576 4063
rect 134524 4020 134576 4029
rect 136732 4063 136784 4072
rect 136732 4029 136741 4063
rect 136741 4029 136775 4063
rect 136775 4029 136784 4063
rect 136732 4020 136784 4029
rect 137836 4020 137888 4072
rect 138940 4063 138992 4072
rect 138940 4029 138949 4063
rect 138949 4029 138983 4063
rect 138983 4029 138992 4063
rect 138940 4020 138992 4029
rect 140044 4063 140096 4072
rect 140044 4029 140053 4063
rect 140053 4029 140087 4063
rect 140087 4029 140096 4063
rect 140044 4020 140096 4029
rect 141148 4063 141200 4072
rect 141148 4029 141157 4063
rect 141157 4029 141191 4063
rect 141191 4029 141200 4063
rect 141148 4020 141200 4029
rect 142252 4020 142304 4072
rect 143448 4020 143500 4072
rect 144460 4063 144512 4072
rect 144460 4029 144469 4063
rect 144469 4029 144503 4063
rect 144503 4029 144512 4063
rect 144460 4020 144512 4029
rect 145564 4063 145616 4072
rect 145564 4029 145573 4063
rect 145573 4029 145607 4063
rect 145607 4029 145616 4063
rect 145564 4020 145616 4029
rect 146668 4063 146720 4072
rect 146668 4029 146677 4063
rect 146677 4029 146711 4063
rect 146711 4029 146720 4063
rect 146668 4020 146720 4029
rect 147772 4020 147824 4072
rect 148876 4020 148928 4072
rect 152188 4063 152240 4072
rect 152188 4029 152197 4063
rect 152197 4029 152231 4063
rect 152231 4029 152240 4063
rect 152188 4020 152240 4029
rect 153292 4020 153344 4072
rect 154396 4063 154448 4072
rect 154396 4029 154405 4063
rect 154405 4029 154439 4063
rect 154439 4029 154448 4063
rect 154396 4020 154448 4029
rect 155500 4063 155552 4072
rect 155500 4029 155509 4063
rect 155509 4029 155543 4063
rect 155543 4029 155552 4063
rect 155500 4020 155552 4029
rect 157708 4063 157760 4072
rect 157708 4029 157717 4063
rect 157717 4029 157751 4063
rect 157751 4029 157760 4063
rect 157708 4020 157760 4029
rect 158812 4020 158864 4072
rect 159916 4063 159968 4072
rect 159916 4029 159925 4063
rect 159925 4029 159959 4063
rect 159959 4029 159968 4063
rect 159916 4020 159968 4029
rect 161020 4063 161072 4072
rect 161020 4029 161029 4063
rect 161029 4029 161063 4063
rect 161063 4029 161072 4063
rect 161020 4020 161072 4029
rect 162124 4063 162176 4072
rect 162124 4029 162133 4063
rect 162133 4029 162167 4063
rect 162167 4029 162176 4063
rect 162124 4020 162176 4029
rect 165436 4063 165488 4072
rect 165436 4029 165445 4063
rect 165445 4029 165479 4063
rect 165479 4029 165488 4063
rect 165436 4020 165488 4029
rect 166540 4063 166592 4072
rect 166540 4029 166549 4063
rect 166549 4029 166583 4063
rect 166583 4029 166592 4063
rect 166540 4020 166592 4029
rect 167644 4063 167696 4072
rect 167644 4029 167653 4063
rect 167653 4029 167687 4063
rect 167687 4029 167696 4063
rect 167644 4020 167696 4029
rect 168748 4020 168800 4072
rect 169852 4020 169904 4072
rect 173072 4020 173124 4072
rect 174268 4020 174320 4072
rect 175740 4063 175792 4072
rect 175740 4029 175749 4063
rect 175749 4029 175783 4063
rect 175783 4029 175792 4063
rect 175740 4020 175792 4029
rect 177304 4020 177356 4072
rect 103520 3952 103572 4004
rect 101404 3927 101456 3936
rect 101404 3893 101413 3927
rect 101413 3893 101447 3927
rect 101447 3893 101456 3927
rect 101404 3884 101456 3893
rect 102048 3927 102100 3936
rect 102048 3893 102057 3927
rect 102057 3893 102091 3927
rect 102091 3893 102100 3927
rect 102048 3884 102100 3893
rect 103060 3884 103112 3936
rect 103888 3927 103940 3936
rect 103888 3893 103897 3927
rect 103897 3893 103931 3927
rect 103931 3893 103940 3927
rect 103888 3884 103940 3893
rect 176844 3952 176896 4004
rect 107292 3927 107344 3936
rect 107292 3893 107301 3927
rect 107301 3893 107335 3927
rect 107335 3893 107344 3927
rect 107292 3884 107344 3893
rect 107476 3884 107528 3936
rect 19606 3782 19658 3834
rect 19670 3782 19722 3834
rect 19734 3782 19786 3834
rect 19798 3782 19850 3834
rect 50326 3782 50378 3834
rect 50390 3782 50442 3834
rect 50454 3782 50506 3834
rect 50518 3782 50570 3834
rect 81046 3782 81098 3834
rect 81110 3782 81162 3834
rect 81174 3782 81226 3834
rect 81238 3782 81290 3834
rect 111766 3782 111818 3834
rect 111830 3782 111882 3834
rect 111894 3782 111946 3834
rect 111958 3782 112010 3834
rect 142486 3782 142538 3834
rect 142550 3782 142602 3834
rect 142614 3782 142666 3834
rect 142678 3782 142730 3834
rect 173206 3782 173258 3834
rect 173270 3782 173322 3834
rect 173334 3782 173386 3834
rect 173398 3782 173450 3834
rect 3148 3723 3200 3732
rect 3148 3689 3157 3723
rect 3157 3689 3191 3723
rect 3191 3689 3200 3723
rect 3148 3680 3200 3689
rect 1952 3655 2004 3664
rect 1952 3621 1961 3655
rect 1961 3621 1995 3655
rect 1995 3621 2004 3655
rect 1952 3612 2004 3621
rect 9956 3612 10008 3664
rect 12256 3655 12308 3664
rect 3332 3587 3384 3596
rect 1492 3476 1544 3528
rect 3332 3553 3341 3587
rect 3341 3553 3375 3587
rect 3375 3553 3384 3587
rect 3332 3544 3384 3553
rect 4804 3544 4856 3596
rect 6276 3544 6328 3596
rect 9588 3587 9640 3596
rect 9588 3553 9597 3587
rect 9597 3553 9631 3587
rect 9631 3553 9640 3587
rect 9588 3544 9640 3553
rect 10324 3587 10376 3596
rect 10324 3553 10333 3587
rect 10333 3553 10367 3587
rect 10367 3553 10376 3587
rect 10324 3544 10376 3553
rect 10692 3544 10744 3596
rect 12256 3621 12265 3655
rect 12265 3621 12299 3655
rect 12299 3621 12308 3655
rect 12256 3612 12308 3621
rect 12348 3612 12400 3664
rect 13728 3655 13780 3664
rect 13360 3587 13412 3596
rect 13360 3553 13369 3587
rect 13369 3553 13403 3587
rect 13403 3553 13412 3587
rect 13360 3544 13412 3553
rect 13728 3621 13737 3655
rect 13737 3621 13771 3655
rect 13771 3621 13780 3655
rect 13728 3612 13780 3621
rect 14832 3655 14884 3664
rect 14832 3621 14841 3655
rect 14841 3621 14875 3655
rect 14875 3621 14884 3655
rect 14832 3612 14884 3621
rect 15660 3612 15712 3664
rect 18880 3655 18932 3664
rect 756 3408 808 3460
rect 10140 3476 10192 3528
rect 14740 3476 14792 3528
rect 16580 3544 16632 3596
rect 16764 3544 16816 3596
rect 16948 3544 17000 3596
rect 18052 3587 18104 3596
rect 18052 3553 18061 3587
rect 18061 3553 18095 3587
rect 18095 3553 18104 3587
rect 18052 3544 18104 3553
rect 18880 3621 18889 3655
rect 18889 3621 18923 3655
rect 18923 3621 18932 3655
rect 18880 3612 18932 3621
rect 19156 3544 19208 3596
rect 33140 3680 33192 3732
rect 33232 3680 33284 3732
rect 45468 3680 45520 3732
rect 21272 3544 21324 3596
rect 21364 3544 21416 3596
rect 22468 3587 22520 3596
rect 22468 3553 22477 3587
rect 22477 3553 22511 3587
rect 22511 3553 22520 3587
rect 22468 3544 22520 3553
rect 23572 3587 23624 3596
rect 23572 3553 23581 3587
rect 23581 3553 23615 3587
rect 23615 3553 23624 3587
rect 23572 3544 23624 3553
rect 28816 3612 28868 3664
rect 40040 3612 40092 3664
rect 41420 3612 41472 3664
rect 62212 3612 62264 3664
rect 70676 3680 70728 3732
rect 70768 3680 70820 3732
rect 72700 3680 72752 3732
rect 73252 3680 73304 3732
rect 75276 3680 75328 3732
rect 75828 3680 75880 3732
rect 79048 3680 79100 3732
rect 79416 3723 79468 3732
rect 79416 3689 79425 3723
rect 79425 3689 79459 3723
rect 79459 3689 79468 3723
rect 79416 3680 79468 3689
rect 80060 3680 80112 3732
rect 68284 3655 68336 3664
rect 24676 3544 24728 3596
rect 25780 3544 25832 3596
rect 26884 3587 26936 3596
rect 26884 3553 26893 3587
rect 26893 3553 26927 3587
rect 26927 3553 26936 3587
rect 26884 3544 26936 3553
rect 27988 3587 28040 3596
rect 27988 3553 27997 3587
rect 27997 3553 28031 3587
rect 28031 3553 28040 3587
rect 27988 3544 28040 3553
rect 28172 3544 28224 3596
rect 30380 3544 30432 3596
rect 31300 3587 31352 3596
rect 31300 3553 31309 3587
rect 31309 3553 31343 3587
rect 31343 3553 31352 3587
rect 31300 3544 31352 3553
rect 32404 3587 32456 3596
rect 32404 3553 32413 3587
rect 32413 3553 32447 3587
rect 32447 3553 32456 3587
rect 32404 3544 32456 3553
rect 33508 3587 33560 3596
rect 33508 3553 33517 3587
rect 33517 3553 33551 3587
rect 33551 3553 33560 3587
rect 33508 3544 33560 3553
rect 34612 3587 34664 3596
rect 34612 3553 34621 3587
rect 34621 3553 34655 3587
rect 34655 3553 34664 3587
rect 34612 3544 34664 3553
rect 35716 3587 35768 3596
rect 35716 3553 35725 3587
rect 35725 3553 35759 3587
rect 35759 3553 35768 3587
rect 35716 3544 35768 3553
rect 21548 3476 21600 3528
rect 22284 3476 22336 3528
rect 24124 3476 24176 3528
rect 25320 3476 25372 3528
rect 37464 3544 37516 3596
rect 37924 3587 37976 3596
rect 37924 3553 37933 3587
rect 37933 3553 37967 3587
rect 37967 3553 37976 3587
rect 37924 3544 37976 3553
rect 38200 3544 38252 3596
rect 39580 3544 39632 3596
rect 39764 3587 39816 3596
rect 39764 3553 39773 3587
rect 39773 3553 39807 3587
rect 39807 3553 39816 3587
rect 39764 3544 39816 3553
rect 40868 3544 40920 3596
rect 41972 3587 42024 3596
rect 41972 3553 41981 3587
rect 41981 3553 42015 3587
rect 42015 3553 42024 3587
rect 41972 3544 42024 3553
rect 43076 3587 43128 3596
rect 43076 3553 43085 3587
rect 43085 3553 43119 3587
rect 43119 3553 43128 3587
rect 43076 3544 43128 3553
rect 44180 3587 44232 3596
rect 44180 3553 44189 3587
rect 44189 3553 44223 3587
rect 44223 3553 44232 3587
rect 44180 3544 44232 3553
rect 45284 3544 45336 3596
rect 46388 3587 46440 3596
rect 46388 3553 46397 3587
rect 46397 3553 46431 3587
rect 46431 3553 46440 3587
rect 46388 3544 46440 3553
rect 47492 3587 47544 3596
rect 47492 3553 47501 3587
rect 47501 3553 47535 3587
rect 47535 3553 47544 3587
rect 47492 3544 47544 3553
rect 48596 3587 48648 3596
rect 48596 3553 48605 3587
rect 48605 3553 48639 3587
rect 48639 3553 48648 3587
rect 48596 3544 48648 3553
rect 49700 3587 49752 3596
rect 49700 3553 49709 3587
rect 49709 3553 49743 3587
rect 49743 3553 49752 3587
rect 49700 3544 49752 3553
rect 54116 3587 54168 3596
rect 54116 3553 54125 3587
rect 54125 3553 54159 3587
rect 54159 3553 54168 3587
rect 54116 3544 54168 3553
rect 55220 3587 55272 3596
rect 55220 3553 55229 3587
rect 55229 3553 55263 3587
rect 55263 3553 55272 3587
rect 55220 3544 55272 3553
rect 56324 3544 56376 3596
rect 57428 3587 57480 3596
rect 57428 3553 57437 3587
rect 57437 3553 57471 3587
rect 57471 3553 57480 3587
rect 57428 3544 57480 3553
rect 58532 3587 58584 3596
rect 58532 3553 58541 3587
rect 58541 3553 58575 3587
rect 58575 3553 58584 3587
rect 58532 3544 58584 3553
rect 59636 3587 59688 3596
rect 59636 3553 59645 3587
rect 59645 3553 59679 3587
rect 59679 3553 59688 3587
rect 59636 3544 59688 3553
rect 60648 3587 60700 3596
rect 60648 3553 60657 3587
rect 60657 3553 60691 3587
rect 60691 3553 60700 3587
rect 60648 3544 60700 3553
rect 61752 3544 61804 3596
rect 62856 3587 62908 3596
rect 62856 3553 62865 3587
rect 62865 3553 62899 3587
rect 62899 3553 62908 3587
rect 62856 3544 62908 3553
rect 63960 3587 64012 3596
rect 63960 3553 63969 3587
rect 63969 3553 64003 3587
rect 64003 3553 64012 3587
rect 63960 3544 64012 3553
rect 65064 3587 65116 3596
rect 65064 3553 65073 3587
rect 65073 3553 65107 3587
rect 65107 3553 65116 3587
rect 65064 3544 65116 3553
rect 66536 3544 66588 3596
rect 67732 3544 67784 3596
rect 68284 3621 68293 3655
rect 68293 3621 68327 3655
rect 68327 3621 68336 3655
rect 68284 3612 68336 3621
rect 69664 3612 69716 3664
rect 69848 3612 69900 3664
rect 69940 3612 69992 3664
rect 72424 3612 72476 3664
rect 76288 3655 76340 3664
rect 76288 3621 76297 3655
rect 76297 3621 76331 3655
rect 76331 3621 76340 3655
rect 76288 3612 76340 3621
rect 76748 3612 76800 3664
rect 80428 3655 80480 3664
rect 69112 3544 69164 3596
rect 69388 3587 69440 3596
rect 69388 3553 69406 3587
rect 69406 3553 69440 3587
rect 69388 3544 69440 3553
rect 69572 3544 69624 3596
rect 70860 3544 70912 3596
rect 71228 3544 71280 3596
rect 73436 3587 73488 3596
rect 73436 3553 73445 3587
rect 73445 3553 73479 3587
rect 73479 3553 73488 3587
rect 73436 3544 73488 3553
rect 75736 3544 75788 3596
rect 76012 3544 76064 3596
rect 78220 3544 78272 3596
rect 36452 3476 36504 3528
rect 45008 3476 45060 3528
rect 75828 3476 75880 3528
rect 80060 3544 80112 3596
rect 80428 3621 80437 3655
rect 80437 3621 80471 3655
rect 80471 3621 80480 3655
rect 80428 3612 80480 3621
rect 80612 3723 80664 3732
rect 80612 3689 80621 3723
rect 80621 3689 80655 3723
rect 80655 3689 80664 3723
rect 80612 3680 80664 3689
rect 81440 3680 81492 3732
rect 81808 3680 81860 3732
rect 83464 3680 83516 3732
rect 85028 3723 85080 3732
rect 80980 3544 81032 3596
rect 81532 3587 81584 3596
rect 80888 3476 80940 3528
rect 22008 3408 22060 3460
rect 35348 3408 35400 3460
rect 35440 3408 35492 3460
rect 46204 3408 46256 3460
rect 61568 3408 61620 3460
rect 72700 3408 72752 3460
rect 74724 3408 74776 3460
rect 78864 3408 78916 3460
rect 79048 3451 79100 3460
rect 79048 3417 79057 3451
rect 79057 3417 79091 3451
rect 79091 3417 79100 3451
rect 79048 3408 79100 3417
rect 79232 3408 79284 3460
rect 2688 3383 2740 3392
rect 2688 3349 2697 3383
rect 2697 3349 2731 3383
rect 2731 3349 2740 3383
rect 2688 3340 2740 3349
rect 11980 3340 12032 3392
rect 12164 3340 12216 3392
rect 13084 3340 13136 3392
rect 14372 3340 14424 3392
rect 15384 3340 15436 3392
rect 18696 3340 18748 3392
rect 18788 3340 18840 3392
rect 19064 3340 19116 3392
rect 20904 3340 20956 3392
rect 20996 3340 21048 3392
rect 22652 3340 22704 3392
rect 34244 3340 34296 3392
rect 34336 3340 34388 3392
rect 45376 3340 45428 3392
rect 67548 3383 67600 3392
rect 67548 3349 67557 3383
rect 67557 3349 67591 3383
rect 67591 3349 67600 3383
rect 67548 3340 67600 3349
rect 69756 3383 69808 3392
rect 69756 3349 69765 3383
rect 69765 3349 69799 3383
rect 69799 3349 69808 3383
rect 69756 3340 69808 3349
rect 70032 3340 70084 3392
rect 70492 3340 70544 3392
rect 71228 3340 71280 3392
rect 72332 3340 72384 3392
rect 72976 3383 73028 3392
rect 72976 3349 72985 3383
rect 72985 3349 73019 3383
rect 73019 3349 73028 3383
rect 72976 3340 73028 3349
rect 75092 3340 75144 3392
rect 75276 3340 75328 3392
rect 76288 3383 76340 3392
rect 76288 3349 76297 3383
rect 76297 3349 76331 3383
rect 76331 3349 76340 3383
rect 76288 3340 76340 3349
rect 76656 3340 76708 3392
rect 77852 3340 77904 3392
rect 79324 3340 79376 3392
rect 80612 3408 80664 3460
rect 81532 3553 81541 3587
rect 81541 3553 81575 3587
rect 81575 3553 81584 3587
rect 81532 3544 81584 3553
rect 82176 3612 82228 3664
rect 82360 3612 82412 3664
rect 81808 3544 81860 3596
rect 81900 3476 81952 3528
rect 84108 3544 84160 3596
rect 84384 3544 84436 3596
rect 85028 3689 85037 3723
rect 85037 3689 85071 3723
rect 85071 3689 85080 3723
rect 85028 3680 85080 3689
rect 85764 3680 85816 3732
rect 87328 3680 87380 3732
rect 88708 3680 88760 3732
rect 88892 3680 88944 3732
rect 91652 3723 91704 3732
rect 91652 3689 91661 3723
rect 91661 3689 91695 3723
rect 91695 3689 91704 3723
rect 91652 3680 91704 3689
rect 101680 3680 101732 3732
rect 101772 3680 101824 3732
rect 109316 3723 109368 3732
rect 85212 3612 85264 3664
rect 86868 3612 86920 3664
rect 83556 3476 83608 3528
rect 84660 3519 84712 3528
rect 84660 3485 84669 3519
rect 84669 3485 84703 3519
rect 84703 3485 84712 3519
rect 84660 3476 84712 3485
rect 85488 3587 85540 3596
rect 85488 3553 85497 3587
rect 85497 3553 85531 3587
rect 85531 3553 85540 3587
rect 85488 3544 85540 3553
rect 85672 3587 85724 3596
rect 85672 3553 85681 3587
rect 85681 3553 85715 3587
rect 85715 3553 85724 3587
rect 85672 3544 85724 3553
rect 86500 3544 86552 3596
rect 85396 3476 85448 3528
rect 89536 3655 89588 3664
rect 89536 3621 89545 3655
rect 89545 3621 89579 3655
rect 89579 3621 89588 3655
rect 89536 3612 89588 3621
rect 89720 3612 89772 3664
rect 93952 3655 94004 3664
rect 87328 3544 87380 3596
rect 89168 3587 89220 3596
rect 89168 3553 89177 3587
rect 89177 3553 89211 3587
rect 89211 3553 89220 3587
rect 89168 3544 89220 3553
rect 90180 3587 90232 3596
rect 90180 3553 90189 3587
rect 90189 3553 90223 3587
rect 90223 3553 90232 3587
rect 90180 3544 90232 3553
rect 93952 3621 93961 3655
rect 93961 3621 93995 3655
rect 93995 3621 94004 3655
rect 93952 3612 94004 3621
rect 95608 3612 95660 3664
rect 101404 3612 101456 3664
rect 101864 3612 101916 3664
rect 90916 3544 90968 3596
rect 91928 3544 91980 3596
rect 94688 3544 94740 3596
rect 95516 3544 95568 3596
rect 96252 3544 96304 3596
rect 97448 3587 97500 3596
rect 97448 3553 97457 3587
rect 97457 3553 97491 3587
rect 97491 3553 97500 3587
rect 97448 3544 97500 3553
rect 98552 3544 98604 3596
rect 99656 3587 99708 3596
rect 99656 3553 99665 3587
rect 99665 3553 99699 3587
rect 99699 3553 99708 3587
rect 99656 3544 99708 3553
rect 100760 3544 100812 3596
rect 101956 3544 102008 3596
rect 104072 3587 104124 3596
rect 104072 3553 104081 3587
rect 104081 3553 104115 3587
rect 104115 3553 104124 3587
rect 104072 3544 104124 3553
rect 105176 3587 105228 3596
rect 105176 3553 105185 3587
rect 105185 3553 105219 3587
rect 105219 3553 105228 3587
rect 105176 3544 105228 3553
rect 106280 3587 106332 3596
rect 106280 3553 106289 3587
rect 106289 3553 106323 3587
rect 106323 3553 106332 3587
rect 106280 3544 106332 3553
rect 107384 3587 107436 3596
rect 107384 3553 107393 3587
rect 107393 3553 107427 3587
rect 107427 3553 107436 3587
rect 107384 3544 107436 3553
rect 81440 3408 81492 3460
rect 81532 3408 81584 3460
rect 82544 3408 82596 3460
rect 81072 3340 81124 3392
rect 81164 3340 81216 3392
rect 83740 3340 83792 3392
rect 84292 3408 84344 3460
rect 93308 3476 93360 3528
rect 101404 3476 101456 3528
rect 101588 3476 101640 3528
rect 109316 3689 109325 3723
rect 109325 3689 109359 3723
rect 109359 3689 109368 3723
rect 109316 3680 109368 3689
rect 109960 3723 110012 3732
rect 109960 3689 109969 3723
rect 109969 3689 110003 3723
rect 110003 3689 110012 3723
rect 109960 3680 110012 3689
rect 108488 3544 108540 3596
rect 109224 3544 109276 3596
rect 110696 3587 110748 3596
rect 110696 3553 110705 3587
rect 110705 3553 110739 3587
rect 110739 3553 110748 3587
rect 110696 3544 110748 3553
rect 112076 3544 112128 3596
rect 112904 3587 112956 3596
rect 112904 3553 112913 3587
rect 112913 3553 112947 3587
rect 112947 3553 112956 3587
rect 112904 3544 112956 3553
rect 114008 3544 114060 3596
rect 115112 3587 115164 3596
rect 115112 3553 115121 3587
rect 115121 3553 115155 3587
rect 115155 3553 115164 3587
rect 115112 3544 115164 3553
rect 116216 3587 116268 3596
rect 116216 3553 116225 3587
rect 116225 3553 116259 3587
rect 116259 3553 116268 3587
rect 116216 3544 116268 3553
rect 117320 3587 117372 3596
rect 117320 3553 117329 3587
rect 117329 3553 117363 3587
rect 117363 3553 117372 3587
rect 117320 3544 117372 3553
rect 118424 3587 118476 3596
rect 118424 3553 118433 3587
rect 118433 3553 118467 3587
rect 118467 3553 118476 3587
rect 118424 3544 118476 3553
rect 119528 3544 119580 3596
rect 120540 3587 120592 3596
rect 120540 3553 120549 3587
rect 120549 3553 120583 3587
rect 120583 3553 120592 3587
rect 120540 3544 120592 3553
rect 121644 3587 121696 3596
rect 121644 3553 121653 3587
rect 121653 3553 121687 3587
rect 121687 3553 121696 3587
rect 121644 3544 121696 3553
rect 122748 3587 122800 3596
rect 122748 3553 122757 3587
rect 122757 3553 122791 3587
rect 122791 3553 122800 3587
rect 122748 3544 122800 3553
rect 123852 3544 123904 3596
rect 124956 3587 125008 3596
rect 124956 3553 124965 3587
rect 124965 3553 124999 3587
rect 124999 3553 125008 3587
rect 124956 3544 125008 3553
rect 126060 3587 126112 3596
rect 126060 3553 126069 3587
rect 126069 3553 126103 3587
rect 126103 3553 126112 3587
rect 126060 3544 126112 3553
rect 126980 3544 127032 3596
rect 128268 3587 128320 3596
rect 128268 3553 128277 3587
rect 128277 3553 128311 3587
rect 128311 3553 128320 3587
rect 128268 3544 128320 3553
rect 129004 3587 129056 3596
rect 129004 3553 129013 3587
rect 129013 3553 129047 3587
rect 129047 3553 129056 3587
rect 129004 3544 129056 3553
rect 129372 3544 129424 3596
rect 130200 3544 130252 3596
rect 131580 3544 131632 3596
rect 133788 3587 133840 3596
rect 132316 3476 132368 3528
rect 133788 3553 133797 3587
rect 133797 3553 133831 3587
rect 133831 3553 133840 3587
rect 133788 3544 133840 3553
rect 134892 3544 134944 3596
rect 135628 3544 135680 3596
rect 137100 3587 137152 3596
rect 137100 3553 137109 3587
rect 137109 3553 137143 3587
rect 137143 3553 137152 3587
rect 137100 3544 137152 3553
rect 138204 3587 138256 3596
rect 138204 3553 138213 3587
rect 138213 3553 138247 3587
rect 138247 3553 138256 3587
rect 138204 3544 138256 3553
rect 139308 3587 139360 3596
rect 139308 3553 139317 3587
rect 139317 3553 139351 3587
rect 139351 3553 139360 3587
rect 139308 3544 139360 3553
rect 140412 3544 140464 3596
rect 141516 3587 141568 3596
rect 141516 3553 141525 3587
rect 141525 3553 141559 3587
rect 141559 3553 141568 3587
rect 141516 3544 141568 3553
rect 142804 3544 142856 3596
rect 143724 3587 143776 3596
rect 143724 3553 143733 3587
rect 143733 3553 143767 3587
rect 143767 3553 143776 3587
rect 143724 3544 143776 3553
rect 144828 3544 144880 3596
rect 145932 3587 145984 3596
rect 145932 3553 145941 3587
rect 145941 3553 145975 3587
rect 145975 3553 145984 3587
rect 145932 3544 145984 3553
rect 147036 3587 147088 3596
rect 147036 3553 147045 3587
rect 147045 3553 147079 3587
rect 147079 3553 147088 3587
rect 147036 3544 147088 3553
rect 148140 3587 148192 3596
rect 148140 3553 148149 3587
rect 148149 3553 148183 3587
rect 148183 3553 148192 3587
rect 148140 3544 148192 3553
rect 149244 3587 149296 3596
rect 149244 3553 149253 3587
rect 149253 3553 149287 3587
rect 149287 3553 149296 3587
rect 149244 3544 149296 3553
rect 149980 3587 150032 3596
rect 149980 3553 149989 3587
rect 149989 3553 150023 3587
rect 150023 3553 150032 3587
rect 149980 3544 150032 3553
rect 150348 3544 150400 3596
rect 151176 3544 151228 3596
rect 153660 3587 153712 3596
rect 153660 3553 153669 3587
rect 153669 3553 153703 3587
rect 153703 3553 153712 3587
rect 153660 3544 153712 3553
rect 154764 3587 154816 3596
rect 154764 3553 154773 3587
rect 154773 3553 154807 3587
rect 154807 3553 154816 3587
rect 154764 3544 154816 3553
rect 155868 3544 155920 3596
rect 156604 3544 156656 3596
rect 158168 3544 158220 3596
rect 159180 3587 159232 3596
rect 159180 3553 159189 3587
rect 159189 3553 159223 3587
rect 159223 3553 159232 3587
rect 159180 3544 159232 3553
rect 160284 3587 160336 3596
rect 160284 3553 160293 3587
rect 160293 3553 160327 3587
rect 160327 3553 160336 3587
rect 160284 3544 160336 3553
rect 161388 3544 161440 3596
rect 162492 3587 162544 3596
rect 162492 3553 162501 3587
rect 162501 3553 162535 3587
rect 162535 3553 162544 3587
rect 162492 3544 162544 3553
rect 163596 3587 163648 3596
rect 163596 3553 163605 3587
rect 163605 3553 163639 3587
rect 163639 3553 163648 3587
rect 163596 3544 163648 3553
rect 163228 3476 163280 3528
rect 164424 3544 164476 3596
rect 165804 3544 165856 3596
rect 166908 3587 166960 3596
rect 166908 3553 166917 3587
rect 166917 3553 166951 3587
rect 166951 3553 166960 3587
rect 166908 3544 166960 3553
rect 168012 3587 168064 3596
rect 168012 3553 168021 3587
rect 168021 3553 168055 3587
rect 168055 3553 168064 3587
rect 168012 3544 168064 3553
rect 169116 3587 169168 3596
rect 169116 3553 169125 3587
rect 169125 3553 169159 3587
rect 169159 3553 169168 3587
rect 169116 3544 169168 3553
rect 170220 3587 170272 3596
rect 170220 3553 170229 3587
rect 170229 3553 170263 3587
rect 170263 3553 170272 3587
rect 170220 3544 170272 3553
rect 170956 3587 171008 3596
rect 170956 3553 170965 3587
rect 170965 3553 170999 3587
rect 170999 3553 171008 3587
rect 170956 3544 171008 3553
rect 171324 3544 171376 3596
rect 172152 3544 172204 3596
rect 173532 3544 173584 3596
rect 174636 3544 174688 3596
rect 84568 3340 84620 3392
rect 86776 3408 86828 3460
rect 88064 3408 88116 3460
rect 86592 3340 86644 3392
rect 87052 3383 87104 3392
rect 87052 3349 87061 3383
rect 87061 3349 87095 3383
rect 87095 3349 87104 3383
rect 88524 3383 88576 3392
rect 87052 3340 87104 3349
rect 88524 3349 88533 3383
rect 88533 3349 88567 3383
rect 88567 3349 88576 3383
rect 88524 3340 88576 3349
rect 89076 3340 89128 3392
rect 89168 3340 89220 3392
rect 90824 3408 90876 3460
rect 95148 3408 95200 3460
rect 98092 3408 98144 3460
rect 89628 3340 89680 3392
rect 89812 3340 89864 3392
rect 93492 3340 93544 3392
rect 97632 3383 97684 3392
rect 97632 3349 97641 3383
rect 97641 3349 97675 3383
rect 97675 3349 97684 3383
rect 97632 3340 97684 3349
rect 98828 3383 98880 3392
rect 98828 3349 98837 3383
rect 98837 3349 98871 3383
rect 98871 3349 98880 3383
rect 98828 3340 98880 3349
rect 98920 3340 98972 3392
rect 102048 3408 102100 3460
rect 102324 3408 102376 3460
rect 179420 3408 179472 3460
rect 100484 3383 100536 3392
rect 100484 3349 100493 3383
rect 100493 3349 100527 3383
rect 100527 3349 100536 3383
rect 100484 3340 100536 3349
rect 101864 3340 101916 3392
rect 102232 3383 102284 3392
rect 102232 3349 102241 3383
rect 102241 3349 102275 3383
rect 102275 3349 102284 3383
rect 102232 3340 102284 3349
rect 102876 3383 102928 3392
rect 102876 3349 102885 3383
rect 102885 3349 102919 3383
rect 102919 3349 102928 3383
rect 102876 3340 102928 3349
rect 106464 3383 106516 3392
rect 106464 3349 106473 3383
rect 106473 3349 106507 3383
rect 106507 3349 106516 3383
rect 106464 3340 106516 3349
rect 131948 3383 132000 3392
rect 131948 3349 131957 3383
rect 131957 3349 131991 3383
rect 131991 3349 132000 3383
rect 131948 3340 132000 3349
rect 153752 3340 153804 3392
rect 173900 3383 173952 3392
rect 173900 3349 173909 3383
rect 173909 3349 173943 3383
rect 173943 3349 173952 3383
rect 173900 3340 173952 3349
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 34966 3238 35018 3290
rect 35030 3238 35082 3290
rect 35094 3238 35146 3290
rect 35158 3238 35210 3290
rect 65686 3238 65738 3290
rect 65750 3238 65802 3290
rect 65814 3238 65866 3290
rect 65878 3238 65930 3290
rect 96406 3238 96458 3290
rect 96470 3238 96522 3290
rect 96534 3238 96586 3290
rect 96598 3238 96650 3290
rect 127126 3238 127178 3290
rect 127190 3238 127242 3290
rect 127254 3238 127306 3290
rect 127318 3238 127370 3290
rect 157846 3238 157898 3290
rect 157910 3238 157962 3290
rect 157974 3238 158026 3290
rect 158038 3238 158090 3290
rect 2688 3136 2740 3188
rect 1676 3043 1728 3052
rect 1676 3009 1685 3043
rect 1685 3009 1719 3043
rect 1719 3009 1728 3043
rect 1676 3000 1728 3009
rect 388 2932 440 2984
rect 2228 2932 2280 2984
rect 9956 3068 10008 3120
rect 11888 3068 11940 3120
rect 3700 2975 3752 2984
rect 3700 2941 3709 2975
rect 3709 2941 3743 2975
rect 3743 2941 3752 2975
rect 3700 2932 3752 2941
rect 5172 2975 5224 2984
rect 5172 2941 5181 2975
rect 5181 2941 5215 2975
rect 5215 2941 5224 2975
rect 5172 2932 5224 2941
rect 6644 2932 6696 2984
rect 7748 2932 7800 2984
rect 9220 2975 9272 2984
rect 9220 2941 9229 2975
rect 9229 2941 9263 2975
rect 9263 2941 9272 2975
rect 9220 2932 9272 2941
rect 10048 2907 10100 2916
rect 10048 2873 10057 2907
rect 10057 2873 10091 2907
rect 10091 2873 10100 2907
rect 10048 2864 10100 2873
rect 10968 2907 11020 2916
rect 10968 2873 10977 2907
rect 10977 2873 11011 2907
rect 11011 2873 11020 2907
rect 10968 2864 11020 2873
rect 2964 2796 3016 2848
rect 4620 2839 4672 2848
rect 4620 2805 4629 2839
rect 4629 2805 4663 2839
rect 4663 2805 4672 2839
rect 4620 2796 4672 2805
rect 9864 2796 9916 2848
rect 9956 2796 10008 2848
rect 11060 2839 11112 2848
rect 11060 2805 11069 2839
rect 11069 2805 11103 2839
rect 11103 2805 11112 2839
rect 11060 2796 11112 2805
rect 12072 2975 12124 2984
rect 12072 2941 12081 2975
rect 12081 2941 12115 2975
rect 12115 2941 12124 2975
rect 12072 2932 12124 2941
rect 13176 3136 13228 3188
rect 15384 3136 15436 3188
rect 15476 3136 15528 3188
rect 16396 3136 16448 3188
rect 12532 3068 12584 3120
rect 17684 3111 17736 3120
rect 13360 3000 13412 3052
rect 15200 3000 15252 3052
rect 17684 3077 17693 3111
rect 17693 3077 17727 3111
rect 17727 3077 17736 3111
rect 17684 3068 17736 3077
rect 21088 3068 21140 3120
rect 21272 3136 21324 3188
rect 24308 3136 24360 3188
rect 24492 3179 24544 3188
rect 24492 3145 24501 3179
rect 24501 3145 24535 3179
rect 24535 3145 24544 3179
rect 24492 3136 24544 3145
rect 24584 3136 24636 3188
rect 22376 3068 22428 3120
rect 38660 3136 38712 3188
rect 28080 3068 28132 3120
rect 28172 3068 28224 3120
rect 30656 3068 30708 3120
rect 31576 3068 31628 3120
rect 14004 2975 14056 2984
rect 13084 2864 13136 2916
rect 14004 2941 14013 2975
rect 14013 2941 14047 2975
rect 14047 2941 14056 2975
rect 14004 2932 14056 2941
rect 14280 2975 14332 2984
rect 14280 2941 14289 2975
rect 14289 2941 14323 2975
rect 14323 2941 14332 2975
rect 14280 2932 14332 2941
rect 15660 2932 15712 2984
rect 16396 2932 16448 2984
rect 17500 2975 17552 2984
rect 17500 2941 17509 2975
rect 17509 2941 17543 2975
rect 17543 2941 17552 2975
rect 25412 3000 25464 3052
rect 17500 2932 17552 2941
rect 16212 2907 16264 2916
rect 13176 2796 13228 2848
rect 13268 2796 13320 2848
rect 16212 2873 16221 2907
rect 16221 2873 16255 2907
rect 16255 2873 16264 2907
rect 16212 2864 16264 2873
rect 15568 2796 15620 2848
rect 18512 2864 18564 2916
rect 18972 2864 19024 2916
rect 19892 2932 19944 2984
rect 20628 2975 20680 2984
rect 20628 2941 20637 2975
rect 20637 2941 20671 2975
rect 20671 2941 20680 2975
rect 20628 2932 20680 2941
rect 20904 2975 20956 2984
rect 20904 2941 20913 2975
rect 20913 2941 20947 2975
rect 20947 2941 20956 2975
rect 20904 2932 20956 2941
rect 22652 2975 22704 2984
rect 22652 2941 22661 2975
rect 22661 2941 22695 2975
rect 22695 2941 22704 2975
rect 22652 2932 22704 2941
rect 24308 2932 24360 2984
rect 22008 2864 22060 2916
rect 24584 2932 24636 2984
rect 25320 2864 25372 2916
rect 25504 2907 25556 2916
rect 25504 2873 25513 2907
rect 25513 2873 25547 2907
rect 25547 2873 25556 2907
rect 25504 2864 25556 2873
rect 27896 2907 27948 2916
rect 27896 2873 27905 2907
rect 27905 2873 27939 2907
rect 27939 2873 27948 2907
rect 27896 2864 27948 2873
rect 28816 2907 28868 2916
rect 28816 2873 28825 2907
rect 28825 2873 28859 2907
rect 28859 2873 28868 2907
rect 28816 2864 28868 2873
rect 29092 2932 29144 2984
rect 30196 2975 30248 2984
rect 30196 2941 30205 2975
rect 30205 2941 30239 2975
rect 30239 2941 30248 2975
rect 30196 2932 30248 2941
rect 36452 3068 36504 3120
rect 40960 3136 41012 3188
rect 41052 3136 41104 3188
rect 45100 3136 45152 3188
rect 67548 3179 67600 3188
rect 67548 3145 67557 3179
rect 67557 3145 67591 3179
rect 67591 3145 67600 3179
rect 67548 3136 67600 3145
rect 67640 3136 67692 3188
rect 39120 3068 39172 3120
rect 48044 3068 48096 3120
rect 39028 3000 39080 3052
rect 33232 2975 33284 2984
rect 33232 2941 33241 2975
rect 33241 2941 33275 2975
rect 33275 2941 33284 2975
rect 33232 2932 33284 2941
rect 34336 2975 34388 2984
rect 34336 2941 34345 2975
rect 34345 2941 34379 2975
rect 34379 2941 34388 2975
rect 34336 2932 34388 2941
rect 35440 2975 35492 2984
rect 35440 2941 35449 2975
rect 35449 2941 35483 2975
rect 35483 2941 35492 2975
rect 35440 2932 35492 2941
rect 36820 2932 36872 2984
rect 44272 3000 44324 3052
rect 61568 3000 61620 3052
rect 36268 2864 36320 2916
rect 38384 2907 38436 2916
rect 38384 2873 38393 2907
rect 38393 2873 38427 2907
rect 38427 2873 38436 2907
rect 39120 2907 39172 2916
rect 38384 2864 38436 2873
rect 39120 2873 39129 2907
rect 39129 2873 39163 2907
rect 39163 2873 39172 2907
rect 39120 2864 39172 2873
rect 40132 2932 40184 2984
rect 41236 2975 41288 2984
rect 41236 2941 41245 2975
rect 41245 2941 41279 2975
rect 41279 2941 41288 2975
rect 41236 2932 41288 2941
rect 42340 2975 42392 2984
rect 42340 2941 42349 2975
rect 42349 2941 42383 2975
rect 42383 2941 42392 2975
rect 42340 2932 42392 2941
rect 43444 2932 43496 2984
rect 44548 2975 44600 2984
rect 44548 2941 44557 2975
rect 44557 2941 44591 2975
rect 44591 2941 44600 2975
rect 44548 2932 44600 2941
rect 45652 2975 45704 2984
rect 45652 2941 45661 2975
rect 45661 2941 45695 2975
rect 45695 2941 45704 2975
rect 45652 2932 45704 2941
rect 46756 2975 46808 2984
rect 46756 2941 46765 2975
rect 46765 2941 46799 2975
rect 46799 2941 46808 2975
rect 46756 2932 46808 2941
rect 47860 2932 47912 2984
rect 48964 2975 49016 2984
rect 48964 2941 48973 2975
rect 48973 2941 49007 2975
rect 49007 2941 49016 2975
rect 48964 2932 49016 2941
rect 50068 2975 50120 2984
rect 50068 2941 50077 2975
rect 50077 2941 50111 2975
rect 50111 2941 50120 2975
rect 50068 2932 50120 2941
rect 50804 2975 50856 2984
rect 50804 2941 50813 2975
rect 50813 2941 50847 2975
rect 50847 2941 50856 2975
rect 50804 2932 50856 2941
rect 51908 2932 51960 2984
rect 52276 2975 52328 2984
rect 52276 2941 52285 2975
rect 52285 2941 52319 2975
rect 52319 2941 52328 2975
rect 52276 2932 52328 2941
rect 53012 2932 53064 2984
rect 53380 2932 53432 2984
rect 54484 2932 54536 2984
rect 55588 2975 55640 2984
rect 55588 2941 55597 2975
rect 55597 2941 55631 2975
rect 55631 2941 55640 2975
rect 55588 2932 55640 2941
rect 56692 2975 56744 2984
rect 56692 2941 56701 2975
rect 56701 2941 56735 2975
rect 56735 2941 56744 2975
rect 56692 2932 56744 2941
rect 57796 2975 57848 2984
rect 57796 2941 57805 2975
rect 57805 2941 57839 2975
rect 57839 2941 57848 2975
rect 57796 2932 57848 2941
rect 58900 2932 58952 2984
rect 60004 2975 60056 2984
rect 60004 2941 60013 2975
rect 60013 2941 60047 2975
rect 60047 2941 60056 2975
rect 60004 2932 60056 2941
rect 61016 2975 61068 2984
rect 61016 2941 61025 2975
rect 61025 2941 61059 2975
rect 61059 2941 61068 2975
rect 61016 2932 61068 2941
rect 62120 2975 62172 2984
rect 62120 2941 62129 2975
rect 62129 2941 62163 2975
rect 62163 2941 62172 2975
rect 62120 2932 62172 2941
rect 63224 2975 63276 2984
rect 63224 2941 63233 2975
rect 63233 2941 63267 2975
rect 63267 2941 63276 2975
rect 63224 2932 63276 2941
rect 64328 2932 64380 2984
rect 65432 2975 65484 2984
rect 65432 2941 65441 2975
rect 65441 2941 65475 2975
rect 65475 2941 65484 2975
rect 65432 2932 65484 2941
rect 66628 2932 66680 2984
rect 48320 2864 48372 2916
rect 68008 3000 68060 3052
rect 68560 3136 68612 3188
rect 69940 3136 69992 3188
rect 71872 3136 71924 3188
rect 72332 3179 72384 3188
rect 72332 3145 72341 3179
rect 72341 3145 72375 3179
rect 72375 3145 72384 3179
rect 72332 3136 72384 3145
rect 72516 3179 72568 3188
rect 72516 3145 72525 3179
rect 72525 3145 72559 3179
rect 72559 3145 72568 3179
rect 72516 3136 72568 3145
rect 72608 3136 72660 3188
rect 74540 3136 74592 3188
rect 75092 3136 75144 3188
rect 76288 3136 76340 3188
rect 76564 3179 76616 3188
rect 76564 3145 76573 3179
rect 76573 3145 76607 3179
rect 76607 3145 76616 3179
rect 76564 3136 76616 3145
rect 77852 3136 77904 3188
rect 78128 3136 78180 3188
rect 79324 3136 79376 3188
rect 70032 3068 70084 3120
rect 70308 3111 70360 3120
rect 70308 3077 70317 3111
rect 70317 3077 70351 3111
rect 70351 3077 70360 3111
rect 70308 3068 70360 3077
rect 70400 3068 70452 3120
rect 75920 3068 75972 3120
rect 76748 3068 76800 3120
rect 81164 3136 81216 3188
rect 81808 3136 81860 3188
rect 83280 3136 83332 3188
rect 83924 3136 83976 3188
rect 80704 3111 80756 3120
rect 80704 3077 80713 3111
rect 80713 3077 80747 3111
rect 80747 3077 80756 3111
rect 80704 3068 80756 3077
rect 80888 3068 80940 3120
rect 81532 3068 81584 3120
rect 82728 3068 82780 3120
rect 83740 3068 83792 3120
rect 85764 3136 85816 3188
rect 84844 3068 84896 3120
rect 87696 3136 87748 3188
rect 88524 3136 88576 3188
rect 87236 3068 87288 3120
rect 98920 3136 98972 3188
rect 70768 3000 70820 3052
rect 74908 3000 74960 3052
rect 78864 3000 78916 3052
rect 21272 2796 21324 2848
rect 22100 2796 22152 2848
rect 23204 2796 23256 2848
rect 25412 2796 25464 2848
rect 26516 2796 26568 2848
rect 27620 2796 27672 2848
rect 28724 2796 28776 2848
rect 30932 2796 30984 2848
rect 32036 2839 32088 2848
rect 32036 2805 32045 2839
rect 32045 2805 32079 2839
rect 32079 2805 32088 2839
rect 32036 2796 32088 2805
rect 33140 2796 33192 2848
rect 34244 2796 34296 2848
rect 35348 2796 35400 2848
rect 36452 2796 36504 2848
rect 37556 2796 37608 2848
rect 38660 2796 38712 2848
rect 68652 2907 68704 2916
rect 68652 2873 68661 2907
rect 68661 2873 68695 2907
rect 68695 2873 68704 2907
rect 68652 2864 68704 2873
rect 68836 2839 68888 2848
rect 68836 2805 68845 2839
rect 68845 2805 68879 2839
rect 68879 2805 68888 2839
rect 68836 2796 68888 2805
rect 70216 2864 70268 2916
rect 71320 2864 71372 2916
rect 71596 2932 71648 2984
rect 72148 2932 72200 2984
rect 73620 2975 73672 2984
rect 73620 2941 73629 2975
rect 73629 2941 73663 2975
rect 73663 2941 73672 2975
rect 73620 2932 73672 2941
rect 75460 2864 75512 2916
rect 76656 2864 76708 2916
rect 71596 2796 71648 2848
rect 73436 2796 73488 2848
rect 73528 2796 73580 2848
rect 75552 2839 75604 2848
rect 75552 2805 75561 2839
rect 75561 2805 75595 2839
rect 75595 2805 75604 2839
rect 75552 2796 75604 2805
rect 77576 2932 77628 2984
rect 78956 2932 79008 2984
rect 78772 2864 78824 2916
rect 79048 2907 79100 2916
rect 79048 2873 79057 2907
rect 79057 2873 79091 2907
rect 79091 2873 79100 2907
rect 79048 2864 79100 2873
rect 80060 2932 80112 2984
rect 80336 2932 80388 2984
rect 80704 2932 80756 2984
rect 80888 2932 80940 2984
rect 82084 3000 82136 3052
rect 82360 3000 82412 3052
rect 81532 2975 81584 2984
rect 81532 2941 81541 2975
rect 81541 2941 81575 2975
rect 81575 2941 81584 2975
rect 81532 2932 81584 2941
rect 82176 2932 82228 2984
rect 82268 2975 82320 2984
rect 82268 2941 82277 2975
rect 82277 2941 82311 2975
rect 82311 2941 82320 2975
rect 82268 2932 82320 2941
rect 82544 2975 82596 2984
rect 82544 2941 82553 2975
rect 82553 2941 82587 2975
rect 82587 2941 82596 2975
rect 82544 2932 82596 2941
rect 82820 2975 82872 2984
rect 82820 2941 82829 2975
rect 82829 2941 82863 2975
rect 82863 2941 82872 2975
rect 82820 2932 82872 2941
rect 83740 2975 83792 2984
rect 79324 2796 79376 2848
rect 79692 2796 79744 2848
rect 82728 2864 82780 2916
rect 83004 2864 83056 2916
rect 80428 2796 80480 2848
rect 82084 2796 82136 2848
rect 82176 2796 82228 2848
rect 82636 2796 82688 2848
rect 83740 2941 83749 2975
rect 83749 2941 83783 2975
rect 83783 2941 83792 2975
rect 83740 2932 83792 2941
rect 84016 2932 84068 2984
rect 84292 2932 84344 2984
rect 84660 2932 84712 2984
rect 85304 2864 85356 2916
rect 85856 2932 85908 2984
rect 86592 2975 86644 2984
rect 86592 2941 86601 2975
rect 86601 2941 86635 2975
rect 86635 2941 86644 2975
rect 86592 2932 86644 2941
rect 86776 2975 86828 2984
rect 86776 2941 86785 2975
rect 86785 2941 86819 2975
rect 86819 2941 86828 2975
rect 86776 2932 86828 2941
rect 93124 3068 93176 3120
rect 93308 3068 93360 3120
rect 100484 3136 100536 3188
rect 101680 3136 101732 3188
rect 93216 3000 93268 3052
rect 93584 3000 93636 3052
rect 87696 2975 87748 2984
rect 87696 2941 87705 2975
rect 87705 2941 87739 2975
rect 87739 2941 87748 2975
rect 87972 2975 88024 2984
rect 87696 2932 87748 2941
rect 87972 2941 87997 2975
rect 87997 2941 88024 2975
rect 87972 2932 88024 2941
rect 88156 2932 88208 2984
rect 88340 2932 88392 2984
rect 89444 2932 89496 2984
rect 93308 2932 93360 2984
rect 94412 2932 94464 2984
rect 96068 2932 96120 2984
rect 96620 2932 96672 2984
rect 98460 3000 98512 3052
rect 103888 3068 103940 3120
rect 101312 3043 101364 3052
rect 86500 2864 86552 2916
rect 86868 2864 86920 2916
rect 92204 2864 92256 2916
rect 84292 2796 84344 2848
rect 85488 2796 85540 2848
rect 86592 2796 86644 2848
rect 86684 2796 86736 2848
rect 87696 2796 87748 2848
rect 88432 2796 88484 2848
rect 88892 2796 88944 2848
rect 89168 2796 89220 2848
rect 90088 2796 90140 2848
rect 92572 2796 92624 2848
rect 92756 2864 92808 2916
rect 97264 2864 97316 2916
rect 98736 2932 98788 2984
rect 101312 3009 101321 3043
rect 101321 3009 101355 3043
rect 101355 3009 101364 3043
rect 101312 3000 101364 3009
rect 102140 3000 102192 3052
rect 107476 3000 107528 3052
rect 109132 3000 109184 3052
rect 111616 3000 111668 3052
rect 99932 2932 99984 2984
rect 101128 2932 101180 2984
rect 103704 2975 103756 2984
rect 103704 2941 103713 2975
rect 103713 2941 103747 2975
rect 103747 2941 103756 2975
rect 103704 2932 103756 2941
rect 104440 2975 104492 2984
rect 104440 2941 104449 2975
rect 104449 2941 104483 2975
rect 104483 2941 104492 2975
rect 104440 2932 104492 2941
rect 105544 2975 105596 2984
rect 105544 2941 105553 2975
rect 105553 2941 105587 2975
rect 105587 2941 105596 2975
rect 105544 2932 105596 2941
rect 106648 2975 106700 2984
rect 106648 2941 106657 2975
rect 106657 2941 106691 2975
rect 106691 2941 106700 2975
rect 106648 2932 106700 2941
rect 109868 2932 109920 2984
rect 102876 2864 102928 2916
rect 107200 2864 107252 2916
rect 109592 2864 109644 2916
rect 112444 2932 112496 2984
rect 113180 2932 113232 2984
rect 114284 2932 114336 2984
rect 115204 2932 115256 2984
rect 116400 2932 116452 2984
rect 117136 2975 117188 2984
rect 117136 2941 117145 2975
rect 117145 2941 117179 2975
rect 117179 2941 117188 2975
rect 117136 2932 117188 2941
rect 117780 2975 117832 2984
rect 117780 2941 117789 2975
rect 117789 2941 117823 2975
rect 117823 2941 117832 2975
rect 117780 2932 117832 2941
rect 118792 2975 118844 2984
rect 118792 2941 118801 2975
rect 118801 2941 118835 2975
rect 118835 2941 118844 2975
rect 118792 2932 118844 2941
rect 119896 2975 119948 2984
rect 119896 2941 119905 2975
rect 119905 2941 119939 2975
rect 119939 2941 119948 2975
rect 119896 2932 119948 2941
rect 121736 2932 121788 2984
rect 122380 2975 122432 2984
rect 122380 2941 122389 2975
rect 122389 2941 122423 2975
rect 122423 2941 122432 2975
rect 122380 2932 122432 2941
rect 123116 2975 123168 2984
rect 123116 2941 123125 2975
rect 123125 2941 123159 2975
rect 123159 2941 123168 2975
rect 123116 2932 123168 2941
rect 124220 2975 124272 2984
rect 124220 2941 124229 2975
rect 124229 2941 124263 2975
rect 124263 2941 124272 2975
rect 124220 2932 124272 2941
rect 125324 2975 125376 2984
rect 125324 2941 125333 2975
rect 125333 2941 125367 2975
rect 125367 2941 125376 2975
rect 125324 2932 125376 2941
rect 127072 2932 127124 2984
rect 127624 2975 127676 2984
rect 127624 2941 127633 2975
rect 127633 2941 127667 2975
rect 127667 2941 127676 2975
rect 127624 2932 127676 2941
rect 128636 2975 128688 2984
rect 128636 2941 128645 2975
rect 128645 2941 128679 2975
rect 128679 2941 128688 2975
rect 128636 2932 128688 2941
rect 129740 2975 129792 2984
rect 129740 2941 129749 2975
rect 129749 2941 129783 2975
rect 129783 2941 129792 2975
rect 129740 2932 129792 2941
rect 130844 2975 130896 2984
rect 130844 2941 130853 2975
rect 130853 2941 130887 2975
rect 130887 2941 130896 2975
rect 130844 2932 130896 2941
rect 133052 2975 133104 2984
rect 130476 2864 130528 2916
rect 133052 2941 133061 2975
rect 133061 2941 133095 2975
rect 133095 2941 133104 2975
rect 133052 2932 133104 2941
rect 134156 2975 134208 2984
rect 134156 2941 134165 2975
rect 134165 2941 134199 2975
rect 134199 2941 134208 2975
rect 134156 2932 134208 2941
rect 135260 2975 135312 2984
rect 135260 2941 135269 2975
rect 135269 2941 135303 2975
rect 135303 2941 135312 2975
rect 135260 2932 135312 2941
rect 136364 2975 136416 2984
rect 136364 2941 136373 2975
rect 136373 2941 136407 2975
rect 136407 2941 136416 2975
rect 136364 2932 136416 2941
rect 138112 2975 138164 2984
rect 135996 2864 136048 2916
rect 138112 2941 138121 2975
rect 138121 2941 138155 2975
rect 138155 2941 138164 2975
rect 138112 2932 138164 2941
rect 138756 2975 138808 2984
rect 138756 2941 138765 2975
rect 138765 2941 138799 2975
rect 138799 2941 138808 2975
rect 138756 2932 138808 2941
rect 139676 2975 139728 2984
rect 139676 2941 139685 2975
rect 139685 2941 139719 2975
rect 139719 2941 139728 2975
rect 139676 2932 139728 2941
rect 140780 2975 140832 2984
rect 140780 2941 140789 2975
rect 140789 2941 140823 2975
rect 140823 2941 140832 2975
rect 140780 2932 140832 2941
rect 141884 2975 141936 2984
rect 141884 2941 141893 2975
rect 141893 2941 141927 2975
rect 141927 2941 141936 2975
rect 141884 2932 141936 2941
rect 143356 2975 143408 2984
rect 143356 2941 143365 2975
rect 143365 2941 143399 2975
rect 143399 2941 143408 2975
rect 143356 2932 143408 2941
rect 144092 2975 144144 2984
rect 144092 2941 144101 2975
rect 144101 2941 144135 2975
rect 144135 2941 144144 2975
rect 144092 2932 144144 2941
rect 145196 2975 145248 2984
rect 145196 2941 145205 2975
rect 145205 2941 145239 2975
rect 145239 2941 145248 2975
rect 145196 2932 145248 2941
rect 146300 2975 146352 2984
rect 146300 2941 146309 2975
rect 146309 2941 146343 2975
rect 146343 2941 146352 2975
rect 146300 2932 146352 2941
rect 147404 2975 147456 2984
rect 147404 2941 147413 2975
rect 147413 2941 147447 2975
rect 147447 2941 147456 2975
rect 147404 2932 147456 2941
rect 148600 2975 148652 2984
rect 148600 2941 148609 2975
rect 148609 2941 148643 2975
rect 148643 2941 148652 2975
rect 148600 2932 148652 2941
rect 149612 2975 149664 2984
rect 149612 2941 149621 2975
rect 149621 2941 149655 2975
rect 149655 2941 149664 2975
rect 149612 2932 149664 2941
rect 150716 2975 150768 2984
rect 150716 2941 150725 2975
rect 150725 2941 150759 2975
rect 150759 2941 150768 2975
rect 150716 2932 150768 2941
rect 151820 2975 151872 2984
rect 151820 2941 151829 2975
rect 151829 2941 151863 2975
rect 151863 2941 151872 2975
rect 152556 2975 152608 2984
rect 151820 2932 151872 2941
rect 152556 2941 152565 2975
rect 152565 2941 152599 2975
rect 152599 2941 152608 2975
rect 152556 2932 152608 2941
rect 154028 2975 154080 2984
rect 154028 2941 154037 2975
rect 154037 2941 154071 2975
rect 154071 2941 154080 2975
rect 154028 2932 154080 2941
rect 155132 2975 155184 2984
rect 155132 2941 155141 2975
rect 155141 2941 155175 2975
rect 155175 2941 155184 2975
rect 155132 2932 155184 2941
rect 156236 2975 156288 2984
rect 156236 2941 156245 2975
rect 156245 2941 156279 2975
rect 156279 2941 156288 2975
rect 156236 2932 156288 2941
rect 157340 2975 157392 2984
rect 157340 2941 157349 2975
rect 157349 2941 157383 2975
rect 157383 2941 157392 2975
rect 157340 2932 157392 2941
rect 159088 2975 159140 2984
rect 156972 2864 157024 2916
rect 159088 2941 159097 2975
rect 159097 2941 159131 2975
rect 159131 2941 159140 2975
rect 159088 2932 159140 2941
rect 159732 2975 159784 2984
rect 159732 2941 159741 2975
rect 159741 2941 159775 2975
rect 159775 2941 159784 2975
rect 159732 2932 159784 2941
rect 160652 2975 160704 2984
rect 160652 2941 160661 2975
rect 160661 2941 160695 2975
rect 160695 2941 160704 2975
rect 160652 2932 160704 2941
rect 161756 2975 161808 2984
rect 161756 2941 161765 2975
rect 161765 2941 161799 2975
rect 161799 2941 161808 2975
rect 161756 2932 161808 2941
rect 162860 2975 162912 2984
rect 162860 2941 162869 2975
rect 162869 2941 162903 2975
rect 162903 2941 162912 2975
rect 162860 2932 162912 2941
rect 164332 2975 164384 2984
rect 164332 2941 164341 2975
rect 164341 2941 164375 2975
rect 164375 2941 164384 2975
rect 164332 2932 164384 2941
rect 165068 2975 165120 2984
rect 165068 2941 165077 2975
rect 165077 2941 165111 2975
rect 165111 2941 165120 2975
rect 165068 2932 165120 2941
rect 167092 2932 167144 2984
rect 167276 2975 167328 2984
rect 167276 2941 167285 2975
rect 167285 2941 167319 2975
rect 167319 2941 167328 2975
rect 167276 2932 167328 2941
rect 168380 2975 168432 2984
rect 168380 2941 168389 2975
rect 168389 2941 168423 2975
rect 168423 2941 168432 2975
rect 168380 2932 168432 2941
rect 169760 2932 169812 2984
rect 170588 2975 170640 2984
rect 170588 2941 170597 2975
rect 170597 2941 170631 2975
rect 170631 2941 170640 2975
rect 170588 2932 170640 2941
rect 171692 2975 171744 2984
rect 171692 2941 171701 2975
rect 171701 2941 171735 2975
rect 171735 2941 171744 2975
rect 171692 2932 171744 2941
rect 172796 2975 172848 2984
rect 172796 2941 172805 2975
rect 172805 2941 172839 2975
rect 172839 2941 172848 2975
rect 172796 2932 172848 2941
rect 175004 2975 175056 2984
rect 172428 2864 172480 2916
rect 175004 2941 175013 2975
rect 175013 2941 175047 2975
rect 175047 2941 175056 2975
rect 175004 2932 175056 2941
rect 176108 2975 176160 2984
rect 176108 2941 176117 2975
rect 176117 2941 176151 2975
rect 176151 2941 176160 2975
rect 176108 2932 176160 2941
rect 176936 2975 176988 2984
rect 176936 2941 176945 2975
rect 176945 2941 176979 2975
rect 176979 2941 176988 2975
rect 176936 2932 176988 2941
rect 177304 2932 177356 2984
rect 178316 2864 178368 2916
rect 98828 2796 98880 2848
rect 102324 2839 102376 2848
rect 102324 2805 102333 2839
rect 102333 2805 102367 2839
rect 102367 2805 102376 2839
rect 102324 2796 102376 2805
rect 102508 2796 102560 2848
rect 107292 2796 107344 2848
rect 19606 2694 19658 2746
rect 19670 2694 19722 2746
rect 19734 2694 19786 2746
rect 19798 2694 19850 2746
rect 50326 2694 50378 2746
rect 50390 2694 50442 2746
rect 50454 2694 50506 2746
rect 50518 2694 50570 2746
rect 81046 2694 81098 2746
rect 81110 2694 81162 2746
rect 81174 2694 81226 2746
rect 81238 2694 81290 2746
rect 111766 2694 111818 2746
rect 111830 2694 111882 2746
rect 111894 2694 111946 2746
rect 111958 2694 112010 2746
rect 142486 2694 142538 2746
rect 142550 2694 142602 2746
rect 142614 2694 142666 2746
rect 142678 2694 142730 2746
rect 173206 2694 173258 2746
rect 173270 2694 173322 2746
rect 173334 2694 173386 2746
rect 173398 2694 173450 2746
rect 7380 2592 7432 2644
rect 5816 2567 5868 2576
rect 5816 2533 5825 2567
rect 5825 2533 5859 2567
rect 5859 2533 5868 2567
rect 5816 2524 5868 2533
rect 18604 2592 18656 2644
rect 37280 2592 37332 2644
rect 65340 2592 65392 2644
rect 112 2456 164 2508
rect 1676 2499 1728 2508
rect 1676 2465 1685 2499
rect 1685 2465 1719 2499
rect 1719 2465 1728 2499
rect 1676 2456 1728 2465
rect 2596 2456 2648 2508
rect 4068 2456 4120 2508
rect 5540 2456 5592 2508
rect 7012 2456 7064 2508
rect 8116 2456 8168 2508
rect 8484 2499 8536 2508
rect 8484 2465 8493 2499
rect 8493 2465 8527 2499
rect 8527 2465 8536 2499
rect 8484 2456 8536 2465
rect 9680 2499 9732 2508
rect 9680 2465 9689 2499
rect 9689 2465 9723 2499
rect 9723 2465 9732 2499
rect 9680 2456 9732 2465
rect 11428 2456 11480 2508
rect 5908 2388 5960 2440
rect 12900 2431 12952 2440
rect 12900 2397 12909 2431
rect 12909 2397 12943 2431
rect 12943 2397 12952 2431
rect 12900 2388 12952 2397
rect 32128 2524 32180 2576
rect 36544 2524 36596 2576
rect 40500 2567 40552 2576
rect 40500 2533 40509 2567
rect 40509 2533 40543 2567
rect 40543 2533 40552 2567
rect 40500 2524 40552 2533
rect 41144 2524 41196 2576
rect 45100 2567 45152 2576
rect 15108 2456 15160 2508
rect 16212 2456 16264 2508
rect 17316 2456 17368 2508
rect 17960 2388 18012 2440
rect 18420 2431 18472 2440
rect 18420 2397 18429 2431
rect 18429 2397 18463 2431
rect 18463 2397 18472 2431
rect 18420 2388 18472 2397
rect 19524 2388 19576 2440
rect 20536 2431 20588 2440
rect 20536 2397 20545 2431
rect 20545 2397 20579 2431
rect 20579 2397 20588 2431
rect 20536 2388 20588 2397
rect 21732 2456 21784 2508
rect 22836 2456 22888 2508
rect 23940 2456 23992 2508
rect 25044 2456 25096 2508
rect 26148 2456 26200 2508
rect 27252 2456 27304 2508
rect 28356 2456 28408 2508
rect 29460 2456 29512 2508
rect 30564 2456 30616 2508
rect 31668 2456 31720 2508
rect 32496 2499 32548 2508
rect 32496 2465 32505 2499
rect 32505 2465 32539 2499
rect 32539 2465 32548 2499
rect 32496 2456 32548 2465
rect 32772 2456 32824 2508
rect 33876 2456 33928 2508
rect 35256 2456 35308 2508
rect 36084 2456 36136 2508
rect 37188 2456 37240 2508
rect 38292 2456 38344 2508
rect 39948 2456 40000 2508
rect 41788 2456 41840 2508
rect 45100 2533 45109 2567
rect 45109 2533 45143 2567
rect 45143 2533 45152 2567
rect 45100 2524 45152 2533
rect 45192 2524 45244 2576
rect 47216 2567 47268 2576
rect 47216 2533 47225 2567
rect 47225 2533 47259 2567
rect 47259 2533 47268 2567
rect 47216 2524 47268 2533
rect 49792 2524 49844 2576
rect 50988 2524 51040 2576
rect 52828 2524 52880 2576
rect 54024 2524 54076 2576
rect 44456 2456 44508 2508
rect 48320 2499 48372 2508
rect 33784 2388 33836 2440
rect 26608 2363 26660 2372
rect 2780 2295 2832 2304
rect 2780 2261 2789 2295
rect 2789 2261 2823 2295
rect 2823 2261 2832 2295
rect 2780 2252 2832 2261
rect 7196 2295 7248 2304
rect 7196 2261 7205 2295
rect 7205 2261 7239 2295
rect 7239 2261 7248 2295
rect 7196 2252 7248 2261
rect 8576 2295 8628 2304
rect 8576 2261 8585 2295
rect 8585 2261 8619 2295
rect 8619 2261 8628 2295
rect 8576 2252 8628 2261
rect 8852 2252 8904 2304
rect 15292 2295 15344 2304
rect 15292 2261 15301 2295
rect 15301 2261 15335 2295
rect 15335 2261 15344 2295
rect 15292 2252 15344 2261
rect 16396 2295 16448 2304
rect 16396 2261 16405 2295
rect 16405 2261 16439 2295
rect 16439 2261 16448 2295
rect 16396 2252 16448 2261
rect 17776 2295 17828 2304
rect 17776 2261 17785 2295
rect 17785 2261 17819 2295
rect 17819 2261 17828 2295
rect 17776 2252 17828 2261
rect 21916 2295 21968 2304
rect 21916 2261 21925 2295
rect 21925 2261 21959 2295
rect 21959 2261 21968 2295
rect 21916 2252 21968 2261
rect 23112 2295 23164 2304
rect 23112 2261 23121 2295
rect 23121 2261 23155 2295
rect 23155 2261 23164 2295
rect 23112 2252 23164 2261
rect 24124 2295 24176 2304
rect 24124 2261 24133 2295
rect 24133 2261 24167 2295
rect 24167 2261 24176 2295
rect 24124 2252 24176 2261
rect 25964 2252 26016 2304
rect 26608 2329 26617 2363
rect 26617 2329 26651 2363
rect 26651 2329 26660 2363
rect 26608 2320 26660 2329
rect 27344 2363 27396 2372
rect 27344 2329 27353 2363
rect 27353 2329 27387 2363
rect 27387 2329 27396 2363
rect 27344 2320 27396 2329
rect 28632 2363 28684 2372
rect 28632 2329 28641 2363
rect 28641 2329 28675 2363
rect 28675 2329 28684 2363
rect 28632 2320 28684 2329
rect 29736 2363 29788 2372
rect 29736 2329 29745 2363
rect 29745 2329 29779 2363
rect 29779 2329 29788 2363
rect 29736 2320 29788 2329
rect 29828 2320 29880 2372
rect 47032 2388 47084 2440
rect 48320 2465 48329 2499
rect 48329 2465 48363 2499
rect 48363 2465 48372 2499
rect 48320 2456 48372 2465
rect 49884 2456 49936 2508
rect 51172 2499 51224 2508
rect 51172 2465 51181 2499
rect 51181 2465 51215 2499
rect 51215 2465 51224 2499
rect 51172 2456 51224 2465
rect 53104 2499 53156 2508
rect 53104 2465 53113 2499
rect 53113 2465 53147 2499
rect 53147 2465 53156 2499
rect 53104 2456 53156 2465
rect 61292 2524 61344 2576
rect 62764 2524 62816 2576
rect 63500 2524 63552 2576
rect 65248 2524 65300 2576
rect 56048 2499 56100 2508
rect 56048 2465 56057 2499
rect 56057 2465 56091 2499
rect 56091 2465 56100 2499
rect 56048 2456 56100 2465
rect 57704 2499 57756 2508
rect 57704 2465 57713 2499
rect 57713 2465 57747 2499
rect 57747 2465 57756 2499
rect 57704 2456 57756 2465
rect 59084 2456 59136 2508
rect 59912 2456 59964 2508
rect 60924 2456 60976 2508
rect 66812 2524 66864 2576
rect 67824 2524 67876 2576
rect 69020 2524 69072 2576
rect 71136 2592 71188 2644
rect 71320 2592 71372 2644
rect 77760 2592 77812 2644
rect 81900 2592 81952 2644
rect 83372 2592 83424 2644
rect 73436 2524 73488 2576
rect 73712 2567 73764 2576
rect 73712 2533 73721 2567
rect 73721 2533 73755 2567
rect 73755 2533 73764 2567
rect 73712 2524 73764 2533
rect 73804 2524 73856 2576
rect 75184 2567 75236 2576
rect 75184 2533 75193 2567
rect 75193 2533 75227 2567
rect 75227 2533 75236 2567
rect 75184 2524 75236 2533
rect 77116 2524 77168 2576
rect 77576 2524 77628 2576
rect 80612 2524 80664 2576
rect 81808 2524 81860 2576
rect 84108 2592 84160 2644
rect 84292 2635 84344 2644
rect 84292 2601 84301 2635
rect 84301 2601 84335 2635
rect 84335 2601 84344 2635
rect 84292 2592 84344 2601
rect 84384 2592 84436 2644
rect 85488 2592 85540 2644
rect 83648 2524 83700 2576
rect 67916 2456 67968 2508
rect 68008 2456 68060 2508
rect 69940 2456 69992 2508
rect 75828 2456 75880 2508
rect 80244 2456 80296 2508
rect 82176 2499 82228 2508
rect 53288 2388 53340 2440
rect 30840 2252 30892 2304
rect 31116 2295 31168 2304
rect 31116 2261 31125 2295
rect 31125 2261 31159 2295
rect 31159 2261 31168 2295
rect 31116 2252 31168 2261
rect 34520 2295 34572 2304
rect 34520 2261 34529 2295
rect 34529 2261 34563 2295
rect 34563 2261 34572 2295
rect 34520 2252 34572 2261
rect 37280 2252 37332 2304
rect 37372 2252 37424 2304
rect 38844 2252 38896 2304
rect 39120 2295 39172 2304
rect 39120 2261 39129 2295
rect 39129 2261 39163 2295
rect 39163 2261 39172 2295
rect 39120 2252 39172 2261
rect 39396 2252 39448 2304
rect 40500 2252 40552 2304
rect 41604 2252 41656 2304
rect 42708 2252 42760 2304
rect 43812 2252 43864 2304
rect 44916 2252 44968 2304
rect 46020 2252 46072 2304
rect 47124 2252 47176 2304
rect 48228 2252 48280 2304
rect 49332 2252 49384 2304
rect 50436 2252 50488 2304
rect 51540 2252 51592 2304
rect 52644 2252 52696 2304
rect 53748 2252 53800 2304
rect 54852 2252 54904 2304
rect 55956 2252 56008 2304
rect 57060 2252 57112 2304
rect 58164 2252 58216 2304
rect 59268 2320 59320 2372
rect 64236 2320 64288 2372
rect 64696 2363 64748 2372
rect 64696 2329 64705 2363
rect 64705 2329 64739 2363
rect 64739 2329 64748 2363
rect 64696 2320 64748 2329
rect 71412 2320 71464 2372
rect 60280 2252 60332 2304
rect 61384 2252 61436 2304
rect 62488 2252 62540 2304
rect 63592 2252 63644 2304
rect 65984 2295 66036 2304
rect 65984 2261 65993 2295
rect 65993 2261 66027 2295
rect 66027 2261 66036 2295
rect 65984 2252 66036 2261
rect 66904 2252 66956 2304
rect 68008 2252 68060 2304
rect 69112 2252 69164 2304
rect 70216 2252 70268 2304
rect 71872 2295 71924 2304
rect 71872 2261 71881 2295
rect 71881 2261 71915 2295
rect 71915 2261 71924 2295
rect 71872 2252 71924 2261
rect 71964 2252 72016 2304
rect 72424 2252 72476 2304
rect 81808 2388 81860 2440
rect 82176 2465 82185 2499
rect 82185 2465 82219 2499
rect 82219 2465 82228 2499
rect 82176 2456 82228 2465
rect 82268 2456 82320 2508
rect 82544 2499 82596 2508
rect 82544 2465 82553 2499
rect 82553 2465 82587 2499
rect 82587 2465 82596 2499
rect 82544 2456 82596 2465
rect 82636 2388 82688 2440
rect 76288 2320 76340 2372
rect 77024 2320 77076 2372
rect 82820 2456 82872 2508
rect 84568 2499 84620 2508
rect 84568 2465 84577 2499
rect 84577 2465 84611 2499
rect 84611 2465 84620 2499
rect 84844 2499 84896 2508
rect 84568 2456 84620 2465
rect 84844 2465 84853 2499
rect 84853 2465 84887 2499
rect 84887 2465 84896 2499
rect 84844 2456 84896 2465
rect 85488 2499 85540 2508
rect 85488 2465 85497 2499
rect 85497 2465 85531 2499
rect 85531 2465 85540 2499
rect 85488 2456 85540 2465
rect 85856 2499 85908 2508
rect 85856 2465 85865 2499
rect 85865 2465 85899 2499
rect 85899 2465 85908 2499
rect 85856 2456 85908 2465
rect 86132 2592 86184 2644
rect 89812 2635 89864 2644
rect 86592 2524 86644 2576
rect 86776 2524 86828 2576
rect 87328 2524 87380 2576
rect 88156 2567 88208 2576
rect 88156 2533 88165 2567
rect 88165 2533 88199 2567
rect 88199 2533 88208 2567
rect 88156 2524 88208 2533
rect 89812 2601 89821 2635
rect 89821 2601 89855 2635
rect 89855 2601 89864 2635
rect 89812 2592 89864 2601
rect 93400 2592 93452 2644
rect 87236 2456 87288 2508
rect 87420 2456 87472 2508
rect 88064 2456 88116 2508
rect 83004 2320 83056 2372
rect 86224 2388 86276 2440
rect 87696 2388 87748 2440
rect 87880 2388 87932 2440
rect 88524 2499 88576 2508
rect 88524 2465 88533 2499
rect 88533 2465 88567 2499
rect 88567 2465 88576 2499
rect 88524 2456 88576 2465
rect 92388 2567 92440 2576
rect 92388 2533 92397 2567
rect 92397 2533 92431 2567
rect 92431 2533 92440 2567
rect 92388 2524 92440 2533
rect 93124 2567 93176 2576
rect 93124 2533 93133 2567
rect 93133 2533 93167 2567
rect 93167 2533 93176 2567
rect 93124 2524 93176 2533
rect 93216 2524 93268 2576
rect 94412 2524 94464 2576
rect 96068 2524 96120 2576
rect 96620 2524 96672 2576
rect 98460 2567 98512 2576
rect 98460 2533 98469 2567
rect 98469 2533 98503 2567
rect 98503 2533 98512 2567
rect 98460 2524 98512 2533
rect 98736 2524 98788 2576
rect 99932 2524 99984 2576
rect 101128 2567 101180 2576
rect 101128 2533 101137 2567
rect 101137 2533 101171 2567
rect 101171 2533 101180 2567
rect 101128 2524 101180 2533
rect 101864 2567 101916 2576
rect 101864 2533 101873 2567
rect 101873 2533 101907 2567
rect 101907 2533 101916 2567
rect 101864 2524 101916 2533
rect 102232 2524 102284 2576
rect 103152 2524 103204 2576
rect 106464 2592 106516 2644
rect 107200 2592 107252 2644
rect 103704 2524 103756 2576
rect 104440 2524 104492 2576
rect 105544 2524 105596 2576
rect 106648 2524 106700 2576
rect 109132 2567 109184 2576
rect 109132 2533 109141 2567
rect 109141 2533 109175 2567
rect 109175 2533 109184 2567
rect 109132 2524 109184 2533
rect 109868 2567 109920 2576
rect 109868 2533 109877 2567
rect 109877 2533 109911 2567
rect 109911 2533 109920 2567
rect 109868 2524 109920 2533
rect 111616 2524 111668 2576
rect 112444 2524 112496 2576
rect 113180 2524 113232 2576
rect 114284 2524 114336 2576
rect 115204 2567 115256 2576
rect 115204 2533 115213 2567
rect 115213 2533 115247 2567
rect 115247 2533 115256 2567
rect 115204 2524 115256 2533
rect 116400 2567 116452 2576
rect 116400 2533 116409 2567
rect 116409 2533 116443 2567
rect 116443 2533 116452 2567
rect 116400 2524 116452 2533
rect 117136 2567 117188 2576
rect 117136 2533 117145 2567
rect 117145 2533 117179 2567
rect 117179 2533 117188 2567
rect 117136 2524 117188 2533
rect 117780 2524 117832 2576
rect 118792 2524 118844 2576
rect 119896 2524 119948 2576
rect 121736 2567 121788 2576
rect 121736 2533 121745 2567
rect 121745 2533 121779 2567
rect 121779 2533 121788 2567
rect 121736 2524 121788 2533
rect 122380 2524 122432 2576
rect 123116 2524 123168 2576
rect 124220 2524 124272 2576
rect 125324 2524 125376 2576
rect 127072 2567 127124 2576
rect 127072 2533 127081 2567
rect 127081 2533 127115 2567
rect 127115 2533 127124 2567
rect 127072 2524 127124 2533
rect 127624 2524 127676 2576
rect 128636 2524 128688 2576
rect 129740 2524 129792 2576
rect 130844 2524 130896 2576
rect 131948 2524 132000 2576
rect 133052 2524 133104 2576
rect 134156 2524 134208 2576
rect 135260 2524 135312 2576
rect 136364 2524 136416 2576
rect 138112 2524 138164 2576
rect 138756 2524 138808 2576
rect 139676 2524 139728 2576
rect 140780 2524 140832 2576
rect 141884 2567 141936 2576
rect 141884 2533 141893 2567
rect 141893 2533 141927 2567
rect 141927 2533 141936 2567
rect 141884 2524 141936 2533
rect 143356 2524 143408 2576
rect 144092 2524 144144 2576
rect 145196 2524 145248 2576
rect 146300 2524 146352 2576
rect 147404 2524 147456 2576
rect 148600 2567 148652 2576
rect 148600 2533 148609 2567
rect 148609 2533 148643 2567
rect 148643 2533 148652 2567
rect 148600 2524 148652 2533
rect 149612 2524 149664 2576
rect 150716 2524 150768 2576
rect 151820 2524 151872 2576
rect 153752 2567 153804 2576
rect 153752 2533 153761 2567
rect 153761 2533 153795 2567
rect 153795 2533 153804 2567
rect 153752 2524 153804 2533
rect 154028 2524 154080 2576
rect 155132 2524 155184 2576
rect 156236 2524 156288 2576
rect 157340 2524 157392 2576
rect 159088 2567 159140 2576
rect 159088 2533 159097 2567
rect 159097 2533 159131 2567
rect 159131 2533 159140 2567
rect 159088 2524 159140 2533
rect 159732 2524 159784 2576
rect 160652 2524 160704 2576
rect 161756 2524 161808 2576
rect 162860 2524 162912 2576
rect 164332 2524 164384 2576
rect 165068 2524 165120 2576
rect 167092 2567 167144 2576
rect 167092 2533 167101 2567
rect 167101 2533 167135 2567
rect 167135 2533 167144 2567
rect 167092 2524 167144 2533
rect 167276 2524 167328 2576
rect 168380 2524 168432 2576
rect 169760 2567 169812 2576
rect 169760 2533 169769 2567
rect 169769 2533 169803 2567
rect 169803 2533 169812 2567
rect 169760 2524 169812 2533
rect 170588 2524 170640 2576
rect 171692 2524 171744 2576
rect 172796 2524 172848 2576
rect 173900 2567 173952 2576
rect 173900 2533 173909 2567
rect 173909 2533 173943 2567
rect 173943 2533 173952 2567
rect 173900 2524 173952 2533
rect 175004 2524 175056 2576
rect 176108 2524 176160 2576
rect 176936 2524 176988 2576
rect 89996 2456 90048 2508
rect 90272 2456 90324 2508
rect 92296 2456 92348 2508
rect 93308 2456 93360 2508
rect 95148 2456 95200 2508
rect 102508 2456 102560 2508
rect 108120 2456 108172 2508
rect 110328 2456 110380 2508
rect 132684 2456 132736 2508
rect 151452 2456 151504 2508
rect 164700 2456 164752 2508
rect 95608 2388 95660 2440
rect 98000 2388 98052 2440
rect 100024 2388 100076 2440
rect 107752 2388 107804 2440
rect 109960 2388 110012 2440
rect 76932 2252 76984 2304
rect 80244 2252 80296 2304
rect 80336 2295 80388 2304
rect 80336 2261 80345 2295
rect 80345 2261 80379 2295
rect 80379 2261 80388 2295
rect 80336 2252 80388 2261
rect 82452 2252 82504 2304
rect 82636 2252 82688 2304
rect 84568 2252 84620 2304
rect 86960 2295 87012 2304
rect 86960 2261 86969 2295
rect 86969 2261 87003 2295
rect 87003 2261 87012 2295
rect 86960 2252 87012 2261
rect 87052 2252 87104 2304
rect 87420 2252 87472 2304
rect 87972 2295 88024 2304
rect 87972 2261 87981 2295
rect 87981 2261 88015 2295
rect 88015 2261 88024 2295
rect 87972 2252 88024 2261
rect 88064 2252 88116 2304
rect 90364 2320 90416 2372
rect 90640 2363 90692 2372
rect 90640 2329 90649 2363
rect 90649 2329 90683 2363
rect 90683 2329 90692 2363
rect 90640 2320 90692 2329
rect 91376 2320 91428 2372
rect 94504 2320 94556 2372
rect 90272 2252 90324 2304
rect 91284 2295 91336 2304
rect 91284 2261 91293 2295
rect 91293 2261 91327 2295
rect 91327 2261 91336 2295
rect 91284 2252 91336 2261
rect 92572 2252 92624 2304
rect 96712 2320 96764 2372
rect 98920 2320 98972 2372
rect 101128 2320 101180 2372
rect 108856 2320 108908 2372
rect 111064 2320 111116 2372
rect 102232 2252 102284 2304
rect 103336 2252 103388 2304
rect 104440 2252 104492 2304
rect 105544 2252 105596 2304
rect 106648 2252 106700 2304
rect 106924 2252 106976 2304
rect 112168 2320 112220 2372
rect 114376 2320 114428 2372
rect 116584 2320 116636 2372
rect 125324 2320 125376 2372
rect 130844 2320 130896 2372
rect 147404 2363 147456 2372
rect 147404 2329 147413 2363
rect 147413 2329 147447 2363
rect 147447 2329 147456 2363
rect 147404 2320 147456 2329
rect 175004 2320 175056 2372
rect 113272 2252 113324 2304
rect 115480 2252 115532 2304
rect 117688 2252 117740 2304
rect 118792 2252 118844 2304
rect 119896 2252 119948 2304
rect 120908 2252 120960 2304
rect 122012 2252 122064 2304
rect 123116 2252 123168 2304
rect 124220 2252 124272 2304
rect 126428 2252 126480 2304
rect 127532 2252 127584 2304
rect 128636 2295 128688 2304
rect 128636 2261 128645 2295
rect 128645 2261 128679 2295
rect 128679 2261 128688 2295
rect 128636 2252 128688 2261
rect 129740 2252 129792 2304
rect 131948 2252 132000 2304
rect 133052 2252 133104 2304
rect 134156 2252 134208 2304
rect 135260 2252 135312 2304
rect 136364 2252 136416 2304
rect 137468 2252 137520 2304
rect 138572 2252 138624 2304
rect 139676 2252 139728 2304
rect 140780 2252 140832 2304
rect 141884 2252 141936 2304
rect 142988 2252 143040 2304
rect 144092 2252 144144 2304
rect 145196 2252 145248 2304
rect 146300 2252 146352 2304
rect 148508 2252 148560 2304
rect 149612 2252 149664 2304
rect 150716 2252 150768 2304
rect 151820 2252 151872 2304
rect 152924 2252 152976 2304
rect 154028 2252 154080 2304
rect 155132 2252 155184 2304
rect 156236 2252 156288 2304
rect 157340 2252 157392 2304
rect 158444 2252 158496 2304
rect 159548 2252 159600 2304
rect 160652 2295 160704 2304
rect 160652 2261 160661 2295
rect 160661 2261 160695 2295
rect 160695 2261 160704 2295
rect 160652 2252 160704 2261
rect 161756 2252 161808 2304
rect 162860 2252 162912 2304
rect 163964 2252 164016 2304
rect 165068 2252 165120 2304
rect 166172 2252 166224 2304
rect 167276 2252 167328 2304
rect 168380 2252 168432 2304
rect 169484 2252 169536 2304
rect 170588 2252 170640 2304
rect 171692 2252 171744 2304
rect 172796 2252 172848 2304
rect 173900 2252 173952 2304
rect 176108 2252 176160 2304
rect 177212 2252 177264 2304
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 34966 2150 35018 2202
rect 35030 2150 35082 2202
rect 35094 2150 35146 2202
rect 35158 2150 35210 2202
rect 65686 2150 65738 2202
rect 65750 2150 65802 2202
rect 65814 2150 65866 2202
rect 65878 2150 65930 2202
rect 96406 2150 96458 2202
rect 96470 2150 96522 2202
rect 96534 2150 96586 2202
rect 96598 2150 96650 2202
rect 127126 2150 127178 2202
rect 127190 2150 127242 2202
rect 127254 2150 127306 2202
rect 127318 2150 127370 2202
rect 157846 2150 157898 2202
rect 157910 2150 157962 2202
rect 157974 2150 158026 2202
rect 158038 2150 158090 2202
rect 8576 2048 8628 2100
rect 33416 2048 33468 2100
rect 39120 2048 39172 2100
rect 61292 2048 61344 2100
rect 72976 2048 73028 2100
rect 77116 2091 77168 2100
rect 77116 2057 77125 2091
rect 77125 2057 77159 2091
rect 77159 2057 77168 2091
rect 77116 2048 77168 2057
rect 78588 2048 78640 2100
rect 82268 2048 82320 2100
rect 82820 2048 82872 2100
rect 90364 2048 90416 2100
rect 95148 2048 95200 2100
rect 9680 1980 9732 2032
rect 15384 1980 15436 2032
rect 33784 1980 33836 2032
rect 46940 1980 46992 2032
rect 47032 1980 47084 2032
rect 2780 1912 2832 1964
rect 38752 1912 38804 1964
rect 42616 1912 42668 1964
rect 45192 1912 45244 1964
rect 45376 1912 45428 1964
rect 48320 1912 48372 1964
rect 71964 1980 72016 2032
rect 74540 1980 74592 2032
rect 80336 1980 80388 2032
rect 84200 1980 84252 2032
rect 87696 1980 87748 2032
rect 88340 1980 88392 2032
rect 89628 1980 89680 2032
rect 63684 1912 63736 1964
rect 65156 1912 65208 1964
rect 87972 1912 88024 1964
rect 88156 1912 88208 1964
rect 103152 1912 103204 1964
rect 7196 1844 7248 1896
rect 33324 1844 33376 1896
rect 34520 1844 34572 1896
rect 62672 1844 62724 1896
rect 71596 1844 71648 1896
rect 76380 1844 76432 1896
rect 84016 1844 84068 1896
rect 85396 1844 85448 1896
rect 88524 1844 88576 1896
rect 92756 1844 92808 1896
rect 32496 1776 32548 1828
rect 43260 1776 43312 1828
rect 44732 1776 44784 1828
rect 45376 1776 45428 1828
rect 47952 1776 48004 1828
rect 53288 1776 53340 1828
rect 57612 1776 57664 1828
rect 80244 1776 80296 1828
rect 37280 1708 37332 1760
rect 62580 1708 62632 1760
rect 80060 1708 80112 1760
rect 82176 1776 82228 1828
rect 83188 1776 83240 1828
rect 85856 1776 85908 1828
rect 87328 1776 87380 1828
rect 103060 1776 103112 1828
rect 80612 1708 80664 1760
rect 98368 1708 98420 1760
rect 20536 1640 20588 1692
rect 47584 1640 47636 1692
rect 66076 1640 66128 1692
rect 31116 1572 31168 1624
rect 41420 1572 41472 1624
rect 45836 1572 45888 1624
rect 63040 1572 63092 1624
rect 86960 1640 87012 1692
rect 93492 1640 93544 1692
rect 73436 1572 73488 1624
rect 85120 1572 85172 1624
rect 85212 1572 85264 1624
rect 71412 1504 71464 1556
rect 81440 1504 81492 1556
rect 82084 1504 82136 1556
rect 87236 1572 87288 1624
rect 87788 1572 87840 1624
rect 106924 1640 106976 1692
rect 97632 1504 97684 1556
rect 75736 1436 75788 1488
rect 77024 1436 77076 1488
rect 91652 1436 91704 1488
rect 74632 1368 74684 1420
rect 76932 1368 76984 1420
rect 84568 1368 84620 1420
rect 90640 1368 90692 1420
rect 35624 1300 35676 1352
rect 70308 1300 70360 1352
rect 85672 1300 85724 1352
rect 91284 1300 91336 1352
rect 36728 1232 36780 1284
rect 71504 1232 71556 1284
rect 83464 1232 83516 1284
rect 89812 1232 89864 1284
rect 32956 1164 33008 1216
rect 66628 1164 66680 1216
rect 34428 1096 34480 1148
rect 67732 1096 67784 1148
rect 68744 1096 68796 1148
rect 69572 1096 69624 1148
rect 15292 1028 15344 1080
rect 41512 1028 41564 1080
rect 43628 1028 43680 1080
rect 75552 1028 75604 1080
rect 43904 960 43956 1012
rect 75276 960 75328 1012
rect 88616 960 88668 1012
rect 90180 960 90232 1012
rect 27344 892 27396 944
rect 58256 892 58308 944
rect 24124 824 24176 876
rect 54760 824 54812 876
rect 28632 756 28684 808
rect 58072 756 58124 808
rect 26608 688 26660 740
rect 57152 688 57204 740
rect 29736 620 29788 672
rect 59820 620 59872 672
rect 39304 552 39356 604
rect 68836 552 68888 604
rect 31576 484 31628 536
rect 56968 484 57020 536
rect 23112 416 23164 468
rect 52920 416 52972 468
rect 20904 348 20956 400
rect 48412 348 48464 400
rect 21916 280 21968 332
rect 52552 280 52604 332
rect 25964 212 26016 264
rect 55772 212 55824 264
rect 17776 144 17828 196
rect 44640 144 44692 196
rect 16396 76 16448 128
rect 44364 76 44416 128
<< metal2 >>
rect 754 119200 810 120000
rect 2318 119200 2374 120000
rect 3882 119200 3938 120000
rect 5446 119200 5502 120000
rect 7010 119200 7066 120000
rect 8574 119200 8630 120000
rect 10138 119200 10194 120000
rect 11702 119200 11758 120000
rect 13266 119200 13322 120000
rect 14830 119200 14886 120000
rect 16394 119200 16450 120000
rect 17958 119200 18014 120000
rect 19522 119200 19578 120000
rect 21086 119200 21142 120000
rect 22650 119200 22706 120000
rect 24214 119200 24270 120000
rect 25778 119200 25834 120000
rect 27342 119200 27398 120000
rect 28906 119200 28962 120000
rect 30470 119200 30526 120000
rect 32034 119200 32090 120000
rect 33598 119200 33654 120000
rect 35162 119200 35218 120000
rect 36726 119200 36782 120000
rect 38290 119200 38346 120000
rect 39854 119200 39910 120000
rect 41418 119200 41474 120000
rect 42982 119200 43038 120000
rect 44546 119200 44602 120000
rect 46110 119200 46166 120000
rect 47674 119200 47730 120000
rect 49238 119200 49294 120000
rect 50802 119200 50858 120000
rect 52366 119200 52422 120000
rect 53930 119200 53986 120000
rect 55494 119200 55550 120000
rect 57058 119200 57114 120000
rect 58622 119200 58678 120000
rect 60186 119200 60242 120000
rect 61750 119200 61806 120000
rect 63314 119200 63370 120000
rect 64878 119200 64934 120000
rect 66442 119200 66498 120000
rect 68006 119200 68062 120000
rect 69570 119200 69626 120000
rect 71134 119200 71190 120000
rect 72698 119200 72754 120000
rect 74262 119200 74318 120000
rect 75826 119200 75882 120000
rect 77390 119200 77446 120000
rect 78954 119200 79010 120000
rect 80518 119200 80574 120000
rect 82082 119200 82138 120000
rect 83646 119200 83702 120000
rect 85210 119200 85266 120000
rect 86774 119200 86830 120000
rect 88338 119200 88394 120000
rect 89902 119200 89958 120000
rect 91558 119200 91614 120000
rect 93122 119200 93178 120000
rect 94686 119200 94742 120000
rect 96250 119200 96306 120000
rect 97814 119200 97870 120000
rect 99378 119200 99434 120000
rect 100942 119200 100998 120000
rect 102506 119200 102562 120000
rect 104070 119200 104126 120000
rect 105634 119200 105690 120000
rect 107198 119200 107254 120000
rect 108762 119200 108818 120000
rect 110326 119200 110382 120000
rect 111890 119200 111946 120000
rect 113454 119200 113510 120000
rect 115018 119200 115074 120000
rect 116582 119200 116638 120000
rect 118146 119200 118202 120000
rect 119710 119200 119766 120000
rect 121274 119200 121330 120000
rect 122838 119200 122894 120000
rect 124402 119200 124458 120000
rect 125966 119200 126022 120000
rect 127530 119200 127586 120000
rect 129094 119200 129150 120000
rect 130658 119200 130714 120000
rect 132222 119200 132278 120000
rect 133786 119200 133842 120000
rect 135350 119200 135406 120000
rect 136914 119200 136970 120000
rect 138478 119200 138534 120000
rect 140042 119200 140098 120000
rect 141606 119200 141662 120000
rect 143170 119200 143226 120000
rect 144734 119200 144790 120000
rect 146298 119200 146354 120000
rect 147862 119200 147918 120000
rect 149426 119200 149482 120000
rect 150990 119200 151046 120000
rect 152554 119200 152610 120000
rect 154118 119200 154174 120000
rect 155682 119200 155738 120000
rect 157246 119200 157302 120000
rect 158810 119200 158866 120000
rect 160374 119200 160430 120000
rect 161938 119200 161994 120000
rect 163502 119200 163558 120000
rect 165066 119200 165122 120000
rect 166630 119200 166686 120000
rect 168194 119200 168250 120000
rect 169758 119200 169814 120000
rect 171322 119200 171378 120000
rect 172886 119200 172942 120000
rect 174450 119200 174506 120000
rect 176014 119200 176070 120000
rect 177578 119200 177634 120000
rect 179142 119200 179198 120000
rect 768 117230 796 119200
rect 2332 117298 2360 119200
rect 3896 117298 3924 119200
rect 4220 117532 4516 117552
rect 4276 117530 4300 117532
rect 4356 117530 4380 117532
rect 4436 117530 4460 117532
rect 4298 117478 4300 117530
rect 4362 117478 4374 117530
rect 4436 117478 4438 117530
rect 4276 117476 4300 117478
rect 4356 117476 4380 117478
rect 4436 117476 4460 117478
rect 4220 117456 4516 117476
rect 2320 117292 2372 117298
rect 2320 117234 2372 117240
rect 3884 117292 3936 117298
rect 3884 117234 3936 117240
rect 5460 117230 5488 119200
rect 7024 117298 7052 119200
rect 8588 117298 8616 119200
rect 7012 117292 7064 117298
rect 7012 117234 7064 117240
rect 8576 117292 8628 117298
rect 8576 117234 8628 117240
rect 10152 117230 10180 119200
rect 11716 117298 11744 119200
rect 13280 117298 13308 119200
rect 11704 117292 11756 117298
rect 11704 117234 11756 117240
rect 13268 117292 13320 117298
rect 13268 117234 13320 117240
rect 14844 117230 14872 119200
rect 16408 117314 16436 119200
rect 16408 117298 16620 117314
rect 17972 117298 18000 119200
rect 16408 117292 16632 117298
rect 16408 117286 16580 117292
rect 16580 117234 16632 117240
rect 17960 117292 18012 117298
rect 17960 117234 18012 117240
rect 19536 117230 19564 119200
rect 21100 117298 21128 119200
rect 22664 117298 22692 119200
rect 21088 117292 21140 117298
rect 21088 117234 21140 117240
rect 22652 117292 22704 117298
rect 22652 117234 22704 117240
rect 24228 117230 24256 119200
rect 25792 117298 25820 119200
rect 27356 117298 27384 119200
rect 25780 117292 25832 117298
rect 25780 117234 25832 117240
rect 27344 117292 27396 117298
rect 27344 117234 27396 117240
rect 28920 117230 28948 119200
rect 30484 117298 30512 119200
rect 32048 117298 32076 119200
rect 30472 117292 30524 117298
rect 30472 117234 30524 117240
rect 32036 117292 32088 117298
rect 32036 117234 32088 117240
rect 33612 117230 33640 119200
rect 35176 118130 35204 119200
rect 35176 118102 35388 118130
rect 34940 117532 35236 117552
rect 34996 117530 35020 117532
rect 35076 117530 35100 117532
rect 35156 117530 35180 117532
rect 35018 117478 35020 117530
rect 35082 117478 35094 117530
rect 35156 117478 35158 117530
rect 34996 117476 35020 117478
rect 35076 117476 35100 117478
rect 35156 117476 35180 117478
rect 34940 117456 35236 117476
rect 35360 117298 35388 118102
rect 36740 117298 36768 119200
rect 35348 117292 35400 117298
rect 35348 117234 35400 117240
rect 36728 117292 36780 117298
rect 36728 117234 36780 117240
rect 38304 117230 38332 119200
rect 39868 117314 39896 119200
rect 39868 117298 40080 117314
rect 41432 117298 41460 119200
rect 39868 117292 40092 117298
rect 39868 117286 40040 117292
rect 40040 117234 40092 117240
rect 41420 117292 41472 117298
rect 41420 117234 41472 117240
rect 42996 117230 43024 119200
rect 44560 117298 44588 119200
rect 46124 117298 46152 119200
rect 44548 117292 44600 117298
rect 44548 117234 44600 117240
rect 46112 117292 46164 117298
rect 46112 117234 46164 117240
rect 47688 117230 47716 119200
rect 49252 117298 49280 119200
rect 50816 117314 50844 119200
rect 50816 117298 51120 117314
rect 49240 117292 49292 117298
rect 50816 117292 51132 117298
rect 50816 117286 51080 117292
rect 49240 117234 49292 117240
rect 51080 117234 51132 117240
rect 52380 117230 52408 119200
rect 53944 117298 53972 119200
rect 55508 117298 55536 119200
rect 53932 117292 53984 117298
rect 53932 117234 53984 117240
rect 55496 117292 55548 117298
rect 55496 117234 55548 117240
rect 57072 117230 57100 119200
rect 58636 117298 58664 119200
rect 60200 117298 60228 119200
rect 58624 117292 58676 117298
rect 58624 117234 58676 117240
rect 60188 117292 60240 117298
rect 60188 117234 60240 117240
rect 61764 117230 61792 119200
rect 63328 117314 63356 119200
rect 63328 117298 63540 117314
rect 64892 117298 64920 119200
rect 65660 117532 65956 117552
rect 65716 117530 65740 117532
rect 65796 117530 65820 117532
rect 65876 117530 65900 117532
rect 65738 117478 65740 117530
rect 65802 117478 65814 117530
rect 65876 117478 65878 117530
rect 65716 117476 65740 117478
rect 65796 117476 65820 117478
rect 65876 117476 65900 117478
rect 65660 117456 65956 117476
rect 63328 117292 63552 117298
rect 63328 117286 63500 117292
rect 63500 117234 63552 117240
rect 64880 117292 64932 117298
rect 64880 117234 64932 117240
rect 66456 117230 66484 119200
rect 68020 117298 68048 119200
rect 69584 117298 69612 119200
rect 68008 117292 68060 117298
rect 68008 117234 68060 117240
rect 69572 117292 69624 117298
rect 69572 117234 69624 117240
rect 71148 117230 71176 119200
rect 72712 117298 72740 119200
rect 74276 117298 74304 119200
rect 72700 117292 72752 117298
rect 72700 117234 72752 117240
rect 74264 117292 74316 117298
rect 74264 117234 74316 117240
rect 75840 117230 75868 119200
rect 77404 117298 77432 119200
rect 78968 117298 78996 119200
rect 77392 117292 77444 117298
rect 77392 117234 77444 117240
rect 78956 117292 79008 117298
rect 78956 117234 79008 117240
rect 80532 117230 80560 119200
rect 82096 117298 82124 119200
rect 83660 117298 83688 119200
rect 82084 117292 82136 117298
rect 82084 117234 82136 117240
rect 83648 117292 83700 117298
rect 83648 117234 83700 117240
rect 85224 117230 85252 119200
rect 86788 117314 86816 119200
rect 86788 117298 87000 117314
rect 88352 117298 88380 119200
rect 86788 117292 87012 117298
rect 86788 117286 86960 117292
rect 86960 117234 87012 117240
rect 88340 117292 88392 117298
rect 88340 117234 88392 117240
rect 89916 117230 89944 119200
rect 91572 117298 91600 119200
rect 93136 117298 93164 119200
rect 91560 117292 91612 117298
rect 91560 117234 91612 117240
rect 93124 117292 93176 117298
rect 93124 117234 93176 117240
rect 94700 117230 94728 119200
rect 96264 117298 96292 119200
rect 96380 117532 96676 117552
rect 96436 117530 96460 117532
rect 96516 117530 96540 117532
rect 96596 117530 96620 117532
rect 96458 117478 96460 117530
rect 96522 117478 96534 117530
rect 96596 117478 96598 117530
rect 96436 117476 96460 117478
rect 96516 117476 96540 117478
rect 96596 117476 96620 117478
rect 96380 117456 96676 117476
rect 97828 117298 97856 119200
rect 96252 117292 96304 117298
rect 96252 117234 96304 117240
rect 97816 117292 97868 117298
rect 97816 117234 97868 117240
rect 99392 117230 99420 119200
rect 100956 117298 100984 119200
rect 102520 117298 102548 119200
rect 100944 117292 100996 117298
rect 100944 117234 100996 117240
rect 102508 117292 102560 117298
rect 102508 117234 102560 117240
rect 104084 117230 104112 119200
rect 105648 117298 105676 119200
rect 107212 117298 107240 119200
rect 105636 117292 105688 117298
rect 105636 117234 105688 117240
rect 107200 117292 107252 117298
rect 107200 117234 107252 117240
rect 108776 117230 108804 119200
rect 110340 117314 110368 119200
rect 110340 117298 110460 117314
rect 111904 117298 111932 119200
rect 110340 117292 110472 117298
rect 110340 117286 110420 117292
rect 110420 117234 110472 117240
rect 111892 117292 111944 117298
rect 111892 117234 111944 117240
rect 113468 117230 113496 119200
rect 115032 117298 115060 119200
rect 116596 117298 116624 119200
rect 115020 117292 115072 117298
rect 115020 117234 115072 117240
rect 116584 117292 116636 117298
rect 116584 117234 116636 117240
rect 118160 117230 118188 119200
rect 119724 117298 119752 119200
rect 121288 117314 121316 119200
rect 121288 117298 121500 117314
rect 119712 117292 119764 117298
rect 121288 117292 121512 117298
rect 121288 117286 121460 117292
rect 119712 117234 119764 117240
rect 121460 117234 121512 117240
rect 122852 117230 122880 119200
rect 124416 117298 124444 119200
rect 125980 117298 126008 119200
rect 127100 117532 127396 117552
rect 127156 117530 127180 117532
rect 127236 117530 127260 117532
rect 127316 117530 127340 117532
rect 127178 117478 127180 117530
rect 127242 117478 127254 117530
rect 127316 117478 127318 117530
rect 127156 117476 127180 117478
rect 127236 117476 127260 117478
rect 127316 117476 127340 117478
rect 127100 117456 127396 117476
rect 124404 117292 124456 117298
rect 124404 117234 124456 117240
rect 125968 117292 126020 117298
rect 125968 117234 126020 117240
rect 127544 117230 127572 119200
rect 129108 117298 129136 119200
rect 130672 117298 130700 119200
rect 129096 117292 129148 117298
rect 129096 117234 129148 117240
rect 130660 117292 130712 117298
rect 130660 117234 130712 117240
rect 132236 117230 132264 119200
rect 133800 117314 133828 119200
rect 133800 117298 133920 117314
rect 135364 117298 135392 119200
rect 133800 117292 133932 117298
rect 133800 117286 133880 117292
rect 133880 117234 133932 117240
rect 135352 117292 135404 117298
rect 135352 117234 135404 117240
rect 136928 117230 136956 119200
rect 138492 117298 138520 119200
rect 140056 117298 140084 119200
rect 138480 117292 138532 117298
rect 138480 117234 138532 117240
rect 140044 117292 140096 117298
rect 140044 117234 140096 117240
rect 141620 117230 141648 119200
rect 143184 117298 143212 119200
rect 144748 117298 144776 119200
rect 143172 117292 143224 117298
rect 143172 117234 143224 117240
rect 144736 117292 144788 117298
rect 144736 117234 144788 117240
rect 146312 117230 146340 119200
rect 147876 117298 147904 119200
rect 149440 117298 149468 119200
rect 147864 117292 147916 117298
rect 147864 117234 147916 117240
rect 149428 117292 149480 117298
rect 149428 117234 149480 117240
rect 151004 117230 151032 119200
rect 152568 117298 152596 119200
rect 154132 117298 154160 119200
rect 152556 117292 152608 117298
rect 152556 117234 152608 117240
rect 154120 117292 154172 117298
rect 154120 117234 154172 117240
rect 155696 117230 155724 119200
rect 157260 117314 157288 119200
rect 157820 117532 158116 117552
rect 157876 117530 157900 117532
rect 157956 117530 157980 117532
rect 158036 117530 158060 117532
rect 157898 117478 157900 117530
rect 157962 117478 157974 117530
rect 158036 117478 158038 117530
rect 157876 117476 157900 117478
rect 157956 117476 157980 117478
rect 158036 117476 158060 117478
rect 157820 117456 158116 117476
rect 157260 117298 157380 117314
rect 158824 117298 158852 119200
rect 157260 117292 157392 117298
rect 157260 117286 157340 117292
rect 157340 117234 157392 117240
rect 158812 117292 158864 117298
rect 158812 117234 158864 117240
rect 160388 117230 160416 119200
rect 161952 117298 161980 119200
rect 163516 117298 163544 119200
rect 161940 117292 161992 117298
rect 161940 117234 161992 117240
rect 163504 117292 163556 117298
rect 163504 117234 163556 117240
rect 165080 117230 165108 119200
rect 166644 117298 166672 119200
rect 168208 117314 168236 119200
rect 168208 117298 168420 117314
rect 166632 117292 166684 117298
rect 168208 117292 168432 117298
rect 168208 117286 168380 117292
rect 166632 117234 166684 117240
rect 168380 117234 168432 117240
rect 169772 117230 169800 119200
rect 171336 117298 171364 119200
rect 172900 117298 172928 119200
rect 171324 117292 171376 117298
rect 171324 117234 171376 117240
rect 172888 117292 172940 117298
rect 172888 117234 172940 117240
rect 174464 117230 174492 119200
rect 176028 117298 176056 119200
rect 177592 117298 177620 119200
rect 176016 117292 176068 117298
rect 176016 117234 176068 117240
rect 177580 117292 177632 117298
rect 177580 117234 177632 117240
rect 179156 117230 179184 119200
rect 756 117224 808 117230
rect 756 117166 808 117172
rect 5448 117224 5500 117230
rect 5448 117166 5500 117172
rect 10140 117224 10192 117230
rect 10140 117166 10192 117172
rect 14832 117224 14884 117230
rect 14832 117166 14884 117172
rect 19524 117224 19576 117230
rect 19524 117166 19576 117172
rect 24216 117224 24268 117230
rect 24216 117166 24268 117172
rect 28908 117224 28960 117230
rect 28908 117166 28960 117172
rect 33600 117224 33652 117230
rect 33600 117166 33652 117172
rect 35256 117224 35308 117230
rect 35256 117166 35308 117172
rect 38292 117224 38344 117230
rect 38292 117166 38344 117172
rect 42984 117224 43036 117230
rect 42984 117166 43036 117172
rect 47676 117224 47728 117230
rect 47676 117166 47728 117172
rect 52368 117224 52420 117230
rect 52368 117166 52420 117172
rect 57060 117224 57112 117230
rect 57060 117166 57112 117172
rect 61752 117224 61804 117230
rect 61752 117166 61804 117172
rect 66444 117224 66496 117230
rect 66444 117166 66496 117172
rect 71136 117224 71188 117230
rect 71136 117166 71188 117172
rect 75828 117224 75880 117230
rect 75828 117166 75880 117172
rect 76932 117224 76984 117230
rect 76932 117166 76984 117172
rect 80520 117224 80572 117230
rect 80520 117166 80572 117172
rect 85212 117224 85264 117230
rect 85212 117166 85264 117172
rect 89904 117224 89956 117230
rect 89904 117166 89956 117172
rect 94688 117224 94740 117230
rect 94688 117166 94740 117172
rect 97632 117224 97684 117230
rect 97632 117166 97684 117172
rect 99380 117224 99432 117230
rect 99380 117166 99432 117172
rect 104072 117224 104124 117230
rect 104072 117166 104124 117172
rect 108764 117224 108816 117230
rect 108764 117166 108816 117172
rect 113456 117224 113508 117230
rect 113456 117166 113508 117172
rect 118148 117224 118200 117230
rect 118148 117166 118200 117172
rect 122840 117224 122892 117230
rect 122840 117166 122892 117172
rect 127532 117224 127584 117230
rect 127532 117166 127584 117172
rect 132224 117224 132276 117230
rect 132224 117166 132276 117172
rect 136916 117224 136968 117230
rect 136916 117166 136968 117172
rect 141608 117224 141660 117230
rect 141608 117166 141660 117172
rect 146300 117224 146352 117230
rect 146300 117166 146352 117172
rect 150992 117224 151044 117230
rect 150992 117166 151044 117172
rect 155684 117224 155736 117230
rect 155684 117166 155736 117172
rect 160376 117224 160428 117230
rect 160376 117166 160428 117172
rect 165068 117224 165120 117230
rect 165068 117166 165120 117172
rect 169760 117224 169812 117230
rect 169760 117166 169812 117172
rect 174452 117224 174504 117230
rect 174452 117166 174504 117172
rect 179144 117224 179196 117230
rect 179144 117166 179196 117172
rect 2412 117156 2464 117162
rect 2412 117098 2464 117104
rect 4344 117156 4396 117162
rect 4344 117098 4396 117104
rect 8300 117156 8352 117162
rect 8300 117098 8352 117104
rect 8484 117156 8536 117162
rect 8484 117098 8536 117104
rect 12348 117156 12400 117162
rect 12348 117098 12400 117104
rect 13360 117156 13412 117162
rect 13360 117098 13412 117104
rect 16488 117156 16540 117162
rect 16488 117098 16540 117104
rect 18052 117156 18104 117162
rect 18052 117098 18104 117104
rect 22560 117156 22612 117162
rect 22560 117098 22612 117104
rect 23020 117156 23072 117162
rect 23020 117098 23072 117104
rect 26516 117156 26568 117162
rect 26516 117098 26568 117104
rect 30840 117156 30892 117162
rect 30840 117098 30892 117104
rect 32128 117156 32180 117162
rect 32128 117098 32180 117104
rect 2424 116346 2452 117098
rect 4356 116754 4384 117098
rect 4344 116748 4396 116754
rect 4344 116690 4396 116696
rect 4220 116444 4516 116464
rect 4276 116442 4300 116444
rect 4356 116442 4380 116444
rect 4436 116442 4460 116444
rect 4298 116390 4300 116442
rect 4362 116390 4374 116442
rect 4436 116390 4438 116442
rect 4276 116388 4300 116390
rect 4356 116388 4380 116390
rect 4436 116388 4460 116390
rect 4220 116368 4516 116388
rect 8312 116346 8340 117098
rect 8496 116618 8524 117098
rect 8484 116612 8536 116618
rect 8484 116554 8536 116560
rect 12360 116346 12388 117098
rect 13372 116890 13400 117098
rect 13360 116884 13412 116890
rect 13360 116826 13412 116832
rect 16500 116346 16528 117098
rect 18064 116822 18092 117098
rect 19580 116988 19876 117008
rect 19636 116986 19660 116988
rect 19716 116986 19740 116988
rect 19796 116986 19820 116988
rect 19658 116934 19660 116986
rect 19722 116934 19734 116986
rect 19796 116934 19798 116986
rect 19636 116932 19660 116934
rect 19716 116932 19740 116934
rect 19796 116932 19820 116934
rect 19580 116912 19876 116932
rect 18052 116816 18104 116822
rect 18052 116758 18104 116764
rect 22572 116346 22600 117098
rect 23032 116686 23060 117098
rect 26424 116748 26476 116754
rect 26424 116690 26476 116696
rect 23020 116680 23072 116686
rect 23020 116622 23072 116628
rect 2412 116340 2464 116346
rect 2412 116282 2464 116288
rect 8300 116340 8352 116346
rect 8300 116282 8352 116288
rect 12348 116340 12400 116346
rect 12348 116282 12400 116288
rect 16488 116340 16540 116346
rect 16488 116282 16540 116288
rect 22560 116340 22612 116346
rect 22560 116282 22612 116288
rect 19580 115900 19876 115920
rect 19636 115898 19660 115900
rect 19716 115898 19740 115900
rect 19796 115898 19820 115900
rect 19658 115846 19660 115898
rect 19722 115846 19734 115898
rect 19796 115846 19798 115898
rect 19636 115844 19660 115846
rect 19716 115844 19740 115846
rect 19796 115844 19820 115846
rect 19580 115824 19876 115844
rect 4220 115356 4516 115376
rect 4276 115354 4300 115356
rect 4356 115354 4380 115356
rect 4436 115354 4460 115356
rect 4298 115302 4300 115354
rect 4362 115302 4374 115354
rect 4436 115302 4438 115354
rect 4276 115300 4300 115302
rect 4356 115300 4380 115302
rect 4436 115300 4460 115302
rect 4220 115280 4516 115300
rect 19580 114812 19876 114832
rect 19636 114810 19660 114812
rect 19716 114810 19740 114812
rect 19796 114810 19820 114812
rect 19658 114758 19660 114810
rect 19722 114758 19734 114810
rect 19796 114758 19798 114810
rect 19636 114756 19660 114758
rect 19716 114756 19740 114758
rect 19796 114756 19820 114758
rect 19580 114736 19876 114756
rect 4220 114268 4516 114288
rect 4276 114266 4300 114268
rect 4356 114266 4380 114268
rect 4436 114266 4460 114268
rect 4298 114214 4300 114266
rect 4362 114214 4374 114266
rect 4436 114214 4438 114266
rect 4276 114212 4300 114214
rect 4356 114212 4380 114214
rect 4436 114212 4460 114214
rect 4220 114192 4516 114212
rect 19580 113724 19876 113744
rect 19636 113722 19660 113724
rect 19716 113722 19740 113724
rect 19796 113722 19820 113724
rect 19658 113670 19660 113722
rect 19722 113670 19734 113722
rect 19796 113670 19798 113722
rect 19636 113668 19660 113670
rect 19716 113668 19740 113670
rect 19796 113668 19820 113670
rect 19580 113648 19876 113668
rect 4220 113180 4516 113200
rect 4276 113178 4300 113180
rect 4356 113178 4380 113180
rect 4436 113178 4460 113180
rect 4298 113126 4300 113178
rect 4362 113126 4374 113178
rect 4436 113126 4438 113178
rect 4276 113124 4300 113126
rect 4356 113124 4380 113126
rect 4436 113124 4460 113126
rect 4220 113104 4516 113124
rect 19580 112636 19876 112656
rect 19636 112634 19660 112636
rect 19716 112634 19740 112636
rect 19796 112634 19820 112636
rect 19658 112582 19660 112634
rect 19722 112582 19734 112634
rect 19796 112582 19798 112634
rect 19636 112580 19660 112582
rect 19716 112580 19740 112582
rect 19796 112580 19820 112582
rect 19580 112560 19876 112580
rect 4220 112092 4516 112112
rect 4276 112090 4300 112092
rect 4356 112090 4380 112092
rect 4436 112090 4460 112092
rect 4298 112038 4300 112090
rect 4362 112038 4374 112090
rect 4436 112038 4438 112090
rect 4276 112036 4300 112038
rect 4356 112036 4380 112038
rect 4436 112036 4460 112038
rect 4220 112016 4516 112036
rect 19580 111548 19876 111568
rect 19636 111546 19660 111548
rect 19716 111546 19740 111548
rect 19796 111546 19820 111548
rect 19658 111494 19660 111546
rect 19722 111494 19734 111546
rect 19796 111494 19798 111546
rect 19636 111492 19660 111494
rect 19716 111492 19740 111494
rect 19796 111492 19820 111494
rect 19580 111472 19876 111492
rect 4220 111004 4516 111024
rect 4276 111002 4300 111004
rect 4356 111002 4380 111004
rect 4436 111002 4460 111004
rect 4298 110950 4300 111002
rect 4362 110950 4374 111002
rect 4436 110950 4438 111002
rect 4276 110948 4300 110950
rect 4356 110948 4380 110950
rect 4436 110948 4460 110950
rect 4220 110928 4516 110948
rect 19580 110460 19876 110480
rect 19636 110458 19660 110460
rect 19716 110458 19740 110460
rect 19796 110458 19820 110460
rect 19658 110406 19660 110458
rect 19722 110406 19734 110458
rect 19796 110406 19798 110458
rect 19636 110404 19660 110406
rect 19716 110404 19740 110406
rect 19796 110404 19820 110406
rect 19580 110384 19876 110404
rect 4220 109916 4516 109936
rect 4276 109914 4300 109916
rect 4356 109914 4380 109916
rect 4436 109914 4460 109916
rect 4298 109862 4300 109914
rect 4362 109862 4374 109914
rect 4436 109862 4438 109914
rect 4276 109860 4300 109862
rect 4356 109860 4380 109862
rect 4436 109860 4460 109862
rect 4220 109840 4516 109860
rect 19580 109372 19876 109392
rect 19636 109370 19660 109372
rect 19716 109370 19740 109372
rect 19796 109370 19820 109372
rect 19658 109318 19660 109370
rect 19722 109318 19734 109370
rect 19796 109318 19798 109370
rect 19636 109316 19660 109318
rect 19716 109316 19740 109318
rect 19796 109316 19820 109318
rect 19580 109296 19876 109316
rect 4220 108828 4516 108848
rect 4276 108826 4300 108828
rect 4356 108826 4380 108828
rect 4436 108826 4460 108828
rect 4298 108774 4300 108826
rect 4362 108774 4374 108826
rect 4436 108774 4438 108826
rect 4276 108772 4300 108774
rect 4356 108772 4380 108774
rect 4436 108772 4460 108774
rect 4220 108752 4516 108772
rect 19580 108284 19876 108304
rect 19636 108282 19660 108284
rect 19716 108282 19740 108284
rect 19796 108282 19820 108284
rect 19658 108230 19660 108282
rect 19722 108230 19734 108282
rect 19796 108230 19798 108282
rect 19636 108228 19660 108230
rect 19716 108228 19740 108230
rect 19796 108228 19820 108230
rect 19580 108208 19876 108228
rect 4220 107740 4516 107760
rect 4276 107738 4300 107740
rect 4356 107738 4380 107740
rect 4436 107738 4460 107740
rect 4298 107686 4300 107738
rect 4362 107686 4374 107738
rect 4436 107686 4438 107738
rect 4276 107684 4300 107686
rect 4356 107684 4380 107686
rect 4436 107684 4460 107686
rect 4220 107664 4516 107684
rect 19580 107196 19876 107216
rect 19636 107194 19660 107196
rect 19716 107194 19740 107196
rect 19796 107194 19820 107196
rect 19658 107142 19660 107194
rect 19722 107142 19734 107194
rect 19796 107142 19798 107194
rect 19636 107140 19660 107142
rect 19716 107140 19740 107142
rect 19796 107140 19820 107142
rect 19580 107120 19876 107140
rect 4220 106652 4516 106672
rect 4276 106650 4300 106652
rect 4356 106650 4380 106652
rect 4436 106650 4460 106652
rect 4298 106598 4300 106650
rect 4362 106598 4374 106650
rect 4436 106598 4438 106650
rect 4276 106596 4300 106598
rect 4356 106596 4380 106598
rect 4436 106596 4460 106598
rect 4220 106576 4516 106596
rect 19580 106108 19876 106128
rect 19636 106106 19660 106108
rect 19716 106106 19740 106108
rect 19796 106106 19820 106108
rect 19658 106054 19660 106106
rect 19722 106054 19734 106106
rect 19796 106054 19798 106106
rect 19636 106052 19660 106054
rect 19716 106052 19740 106054
rect 19796 106052 19820 106054
rect 19580 106032 19876 106052
rect 4220 105564 4516 105584
rect 4276 105562 4300 105564
rect 4356 105562 4380 105564
rect 4436 105562 4460 105564
rect 4298 105510 4300 105562
rect 4362 105510 4374 105562
rect 4436 105510 4438 105562
rect 4276 105508 4300 105510
rect 4356 105508 4380 105510
rect 4436 105508 4460 105510
rect 4220 105488 4516 105508
rect 19580 105020 19876 105040
rect 19636 105018 19660 105020
rect 19716 105018 19740 105020
rect 19796 105018 19820 105020
rect 19658 104966 19660 105018
rect 19722 104966 19734 105018
rect 19796 104966 19798 105018
rect 19636 104964 19660 104966
rect 19716 104964 19740 104966
rect 19796 104964 19820 104966
rect 19580 104944 19876 104964
rect 4220 104476 4516 104496
rect 4276 104474 4300 104476
rect 4356 104474 4380 104476
rect 4436 104474 4460 104476
rect 4298 104422 4300 104474
rect 4362 104422 4374 104474
rect 4436 104422 4438 104474
rect 4276 104420 4300 104422
rect 4356 104420 4380 104422
rect 4436 104420 4460 104422
rect 4220 104400 4516 104420
rect 19580 103932 19876 103952
rect 19636 103930 19660 103932
rect 19716 103930 19740 103932
rect 19796 103930 19820 103932
rect 19658 103878 19660 103930
rect 19722 103878 19734 103930
rect 19796 103878 19798 103930
rect 19636 103876 19660 103878
rect 19716 103876 19740 103878
rect 19796 103876 19820 103878
rect 19580 103856 19876 103876
rect 4220 103388 4516 103408
rect 4276 103386 4300 103388
rect 4356 103386 4380 103388
rect 4436 103386 4460 103388
rect 4298 103334 4300 103386
rect 4362 103334 4374 103386
rect 4436 103334 4438 103386
rect 4276 103332 4300 103334
rect 4356 103332 4380 103334
rect 4436 103332 4460 103334
rect 4220 103312 4516 103332
rect 19580 102844 19876 102864
rect 19636 102842 19660 102844
rect 19716 102842 19740 102844
rect 19796 102842 19820 102844
rect 19658 102790 19660 102842
rect 19722 102790 19734 102842
rect 19796 102790 19798 102842
rect 19636 102788 19660 102790
rect 19716 102788 19740 102790
rect 19796 102788 19820 102790
rect 19580 102768 19876 102788
rect 4220 102300 4516 102320
rect 4276 102298 4300 102300
rect 4356 102298 4380 102300
rect 4436 102298 4460 102300
rect 4298 102246 4300 102298
rect 4362 102246 4374 102298
rect 4436 102246 4438 102298
rect 4276 102244 4300 102246
rect 4356 102244 4380 102246
rect 4436 102244 4460 102246
rect 4220 102224 4516 102244
rect 19580 101756 19876 101776
rect 19636 101754 19660 101756
rect 19716 101754 19740 101756
rect 19796 101754 19820 101756
rect 19658 101702 19660 101754
rect 19722 101702 19734 101754
rect 19796 101702 19798 101754
rect 19636 101700 19660 101702
rect 19716 101700 19740 101702
rect 19796 101700 19820 101702
rect 19580 101680 19876 101700
rect 4220 101212 4516 101232
rect 4276 101210 4300 101212
rect 4356 101210 4380 101212
rect 4436 101210 4460 101212
rect 4298 101158 4300 101210
rect 4362 101158 4374 101210
rect 4436 101158 4438 101210
rect 4276 101156 4300 101158
rect 4356 101156 4380 101158
rect 4436 101156 4460 101158
rect 4220 101136 4516 101156
rect 19580 100668 19876 100688
rect 19636 100666 19660 100668
rect 19716 100666 19740 100668
rect 19796 100666 19820 100668
rect 19658 100614 19660 100666
rect 19722 100614 19734 100666
rect 19796 100614 19798 100666
rect 19636 100612 19660 100614
rect 19716 100612 19740 100614
rect 19796 100612 19820 100614
rect 19580 100592 19876 100612
rect 4220 100124 4516 100144
rect 4276 100122 4300 100124
rect 4356 100122 4380 100124
rect 4436 100122 4460 100124
rect 4298 100070 4300 100122
rect 4362 100070 4374 100122
rect 4436 100070 4438 100122
rect 4276 100068 4300 100070
rect 4356 100068 4380 100070
rect 4436 100068 4460 100070
rect 4220 100048 4516 100068
rect 19580 99580 19876 99600
rect 19636 99578 19660 99580
rect 19716 99578 19740 99580
rect 19796 99578 19820 99580
rect 19658 99526 19660 99578
rect 19722 99526 19734 99578
rect 19796 99526 19798 99578
rect 19636 99524 19660 99526
rect 19716 99524 19740 99526
rect 19796 99524 19820 99526
rect 19580 99504 19876 99524
rect 4220 99036 4516 99056
rect 4276 99034 4300 99036
rect 4356 99034 4380 99036
rect 4436 99034 4460 99036
rect 4298 98982 4300 99034
rect 4362 98982 4374 99034
rect 4436 98982 4438 99034
rect 4276 98980 4300 98982
rect 4356 98980 4380 98982
rect 4436 98980 4460 98982
rect 4220 98960 4516 98980
rect 19580 98492 19876 98512
rect 19636 98490 19660 98492
rect 19716 98490 19740 98492
rect 19796 98490 19820 98492
rect 19658 98438 19660 98490
rect 19722 98438 19734 98490
rect 19796 98438 19798 98490
rect 19636 98436 19660 98438
rect 19716 98436 19740 98438
rect 19796 98436 19820 98438
rect 19580 98416 19876 98436
rect 4220 97948 4516 97968
rect 4276 97946 4300 97948
rect 4356 97946 4380 97948
rect 4436 97946 4460 97948
rect 4298 97894 4300 97946
rect 4362 97894 4374 97946
rect 4436 97894 4438 97946
rect 4276 97892 4300 97894
rect 4356 97892 4380 97894
rect 4436 97892 4460 97894
rect 4220 97872 4516 97892
rect 19580 97404 19876 97424
rect 19636 97402 19660 97404
rect 19716 97402 19740 97404
rect 19796 97402 19820 97404
rect 19658 97350 19660 97402
rect 19722 97350 19734 97402
rect 19796 97350 19798 97402
rect 19636 97348 19660 97350
rect 19716 97348 19740 97350
rect 19796 97348 19820 97350
rect 19580 97328 19876 97348
rect 4220 96860 4516 96880
rect 4276 96858 4300 96860
rect 4356 96858 4380 96860
rect 4436 96858 4460 96860
rect 4298 96806 4300 96858
rect 4362 96806 4374 96858
rect 4436 96806 4438 96858
rect 4276 96804 4300 96806
rect 4356 96804 4380 96806
rect 4436 96804 4460 96806
rect 4220 96784 4516 96804
rect 19580 96316 19876 96336
rect 19636 96314 19660 96316
rect 19716 96314 19740 96316
rect 19796 96314 19820 96316
rect 19658 96262 19660 96314
rect 19722 96262 19734 96314
rect 19796 96262 19798 96314
rect 19636 96260 19660 96262
rect 19716 96260 19740 96262
rect 19796 96260 19820 96262
rect 19580 96240 19876 96260
rect 4220 95772 4516 95792
rect 4276 95770 4300 95772
rect 4356 95770 4380 95772
rect 4436 95770 4460 95772
rect 4298 95718 4300 95770
rect 4362 95718 4374 95770
rect 4436 95718 4438 95770
rect 4276 95716 4300 95718
rect 4356 95716 4380 95718
rect 4436 95716 4460 95718
rect 4220 95696 4516 95716
rect 19580 95228 19876 95248
rect 19636 95226 19660 95228
rect 19716 95226 19740 95228
rect 19796 95226 19820 95228
rect 19658 95174 19660 95226
rect 19722 95174 19734 95226
rect 19796 95174 19798 95226
rect 19636 95172 19660 95174
rect 19716 95172 19740 95174
rect 19796 95172 19820 95174
rect 19580 95152 19876 95172
rect 4220 94684 4516 94704
rect 4276 94682 4300 94684
rect 4356 94682 4380 94684
rect 4436 94682 4460 94684
rect 4298 94630 4300 94682
rect 4362 94630 4374 94682
rect 4436 94630 4438 94682
rect 4276 94628 4300 94630
rect 4356 94628 4380 94630
rect 4436 94628 4460 94630
rect 4220 94608 4516 94628
rect 19580 94140 19876 94160
rect 19636 94138 19660 94140
rect 19716 94138 19740 94140
rect 19796 94138 19820 94140
rect 19658 94086 19660 94138
rect 19722 94086 19734 94138
rect 19796 94086 19798 94138
rect 19636 94084 19660 94086
rect 19716 94084 19740 94086
rect 19796 94084 19820 94086
rect 19580 94064 19876 94084
rect 4220 93596 4516 93616
rect 4276 93594 4300 93596
rect 4356 93594 4380 93596
rect 4436 93594 4460 93596
rect 4298 93542 4300 93594
rect 4362 93542 4374 93594
rect 4436 93542 4438 93594
rect 4276 93540 4300 93542
rect 4356 93540 4380 93542
rect 4436 93540 4460 93542
rect 4220 93520 4516 93540
rect 19580 93052 19876 93072
rect 19636 93050 19660 93052
rect 19716 93050 19740 93052
rect 19796 93050 19820 93052
rect 19658 92998 19660 93050
rect 19722 92998 19734 93050
rect 19796 92998 19798 93050
rect 19636 92996 19660 92998
rect 19716 92996 19740 92998
rect 19796 92996 19820 92998
rect 19580 92976 19876 92996
rect 4220 92508 4516 92528
rect 4276 92506 4300 92508
rect 4356 92506 4380 92508
rect 4436 92506 4460 92508
rect 4298 92454 4300 92506
rect 4362 92454 4374 92506
rect 4436 92454 4438 92506
rect 4276 92452 4300 92454
rect 4356 92452 4380 92454
rect 4436 92452 4460 92454
rect 4220 92432 4516 92452
rect 19580 91964 19876 91984
rect 19636 91962 19660 91964
rect 19716 91962 19740 91964
rect 19796 91962 19820 91964
rect 19658 91910 19660 91962
rect 19722 91910 19734 91962
rect 19796 91910 19798 91962
rect 19636 91908 19660 91910
rect 19716 91908 19740 91910
rect 19796 91908 19820 91910
rect 19580 91888 19876 91908
rect 4220 91420 4516 91440
rect 4276 91418 4300 91420
rect 4356 91418 4380 91420
rect 4436 91418 4460 91420
rect 4298 91366 4300 91418
rect 4362 91366 4374 91418
rect 4436 91366 4438 91418
rect 4276 91364 4300 91366
rect 4356 91364 4380 91366
rect 4436 91364 4460 91366
rect 4220 91344 4516 91364
rect 19580 90876 19876 90896
rect 19636 90874 19660 90876
rect 19716 90874 19740 90876
rect 19796 90874 19820 90876
rect 19658 90822 19660 90874
rect 19722 90822 19734 90874
rect 19796 90822 19798 90874
rect 19636 90820 19660 90822
rect 19716 90820 19740 90822
rect 19796 90820 19820 90822
rect 19580 90800 19876 90820
rect 4220 90332 4516 90352
rect 4276 90330 4300 90332
rect 4356 90330 4380 90332
rect 4436 90330 4460 90332
rect 4298 90278 4300 90330
rect 4362 90278 4374 90330
rect 4436 90278 4438 90330
rect 4276 90276 4300 90278
rect 4356 90276 4380 90278
rect 4436 90276 4460 90278
rect 4220 90256 4516 90276
rect 19580 89788 19876 89808
rect 19636 89786 19660 89788
rect 19716 89786 19740 89788
rect 19796 89786 19820 89788
rect 19658 89734 19660 89786
rect 19722 89734 19734 89786
rect 19796 89734 19798 89786
rect 19636 89732 19660 89734
rect 19716 89732 19740 89734
rect 19796 89732 19820 89734
rect 19580 89712 19876 89732
rect 4220 89244 4516 89264
rect 4276 89242 4300 89244
rect 4356 89242 4380 89244
rect 4436 89242 4460 89244
rect 4298 89190 4300 89242
rect 4362 89190 4374 89242
rect 4436 89190 4438 89242
rect 4276 89188 4300 89190
rect 4356 89188 4380 89190
rect 4436 89188 4460 89190
rect 4220 89168 4516 89188
rect 19580 88700 19876 88720
rect 19636 88698 19660 88700
rect 19716 88698 19740 88700
rect 19796 88698 19820 88700
rect 19658 88646 19660 88698
rect 19722 88646 19734 88698
rect 19796 88646 19798 88698
rect 19636 88644 19660 88646
rect 19716 88644 19740 88646
rect 19796 88644 19820 88646
rect 19580 88624 19876 88644
rect 4220 88156 4516 88176
rect 4276 88154 4300 88156
rect 4356 88154 4380 88156
rect 4436 88154 4460 88156
rect 4298 88102 4300 88154
rect 4362 88102 4374 88154
rect 4436 88102 4438 88154
rect 4276 88100 4300 88102
rect 4356 88100 4380 88102
rect 4436 88100 4460 88102
rect 4220 88080 4516 88100
rect 19580 87612 19876 87632
rect 19636 87610 19660 87612
rect 19716 87610 19740 87612
rect 19796 87610 19820 87612
rect 19658 87558 19660 87610
rect 19722 87558 19734 87610
rect 19796 87558 19798 87610
rect 19636 87556 19660 87558
rect 19716 87556 19740 87558
rect 19796 87556 19820 87558
rect 19580 87536 19876 87556
rect 4220 87068 4516 87088
rect 4276 87066 4300 87068
rect 4356 87066 4380 87068
rect 4436 87066 4460 87068
rect 4298 87014 4300 87066
rect 4362 87014 4374 87066
rect 4436 87014 4438 87066
rect 4276 87012 4300 87014
rect 4356 87012 4380 87014
rect 4436 87012 4460 87014
rect 4220 86992 4516 87012
rect 19580 86524 19876 86544
rect 19636 86522 19660 86524
rect 19716 86522 19740 86524
rect 19796 86522 19820 86524
rect 19658 86470 19660 86522
rect 19722 86470 19734 86522
rect 19796 86470 19798 86522
rect 19636 86468 19660 86470
rect 19716 86468 19740 86470
rect 19796 86468 19820 86470
rect 19580 86448 19876 86468
rect 4220 85980 4516 86000
rect 4276 85978 4300 85980
rect 4356 85978 4380 85980
rect 4436 85978 4460 85980
rect 4298 85926 4300 85978
rect 4362 85926 4374 85978
rect 4436 85926 4438 85978
rect 4276 85924 4300 85926
rect 4356 85924 4380 85926
rect 4436 85924 4460 85926
rect 4220 85904 4516 85924
rect 19580 85436 19876 85456
rect 19636 85434 19660 85436
rect 19716 85434 19740 85436
rect 19796 85434 19820 85436
rect 19658 85382 19660 85434
rect 19722 85382 19734 85434
rect 19796 85382 19798 85434
rect 19636 85380 19660 85382
rect 19716 85380 19740 85382
rect 19796 85380 19820 85382
rect 19580 85360 19876 85380
rect 4220 84892 4516 84912
rect 4276 84890 4300 84892
rect 4356 84890 4380 84892
rect 4436 84890 4460 84892
rect 4298 84838 4300 84890
rect 4362 84838 4374 84890
rect 4436 84838 4438 84890
rect 4276 84836 4300 84838
rect 4356 84836 4380 84838
rect 4436 84836 4460 84838
rect 4220 84816 4516 84836
rect 19580 84348 19876 84368
rect 19636 84346 19660 84348
rect 19716 84346 19740 84348
rect 19796 84346 19820 84348
rect 19658 84294 19660 84346
rect 19722 84294 19734 84346
rect 19796 84294 19798 84346
rect 19636 84292 19660 84294
rect 19716 84292 19740 84294
rect 19796 84292 19820 84294
rect 19580 84272 19876 84292
rect 4220 83804 4516 83824
rect 4276 83802 4300 83804
rect 4356 83802 4380 83804
rect 4436 83802 4460 83804
rect 4298 83750 4300 83802
rect 4362 83750 4374 83802
rect 4436 83750 4438 83802
rect 4276 83748 4300 83750
rect 4356 83748 4380 83750
rect 4436 83748 4460 83750
rect 4220 83728 4516 83748
rect 19580 83260 19876 83280
rect 19636 83258 19660 83260
rect 19716 83258 19740 83260
rect 19796 83258 19820 83260
rect 19658 83206 19660 83258
rect 19722 83206 19734 83258
rect 19796 83206 19798 83258
rect 19636 83204 19660 83206
rect 19716 83204 19740 83206
rect 19796 83204 19820 83206
rect 19580 83184 19876 83204
rect 4220 82716 4516 82736
rect 4276 82714 4300 82716
rect 4356 82714 4380 82716
rect 4436 82714 4460 82716
rect 4298 82662 4300 82714
rect 4362 82662 4374 82714
rect 4436 82662 4438 82714
rect 4276 82660 4300 82662
rect 4356 82660 4380 82662
rect 4436 82660 4460 82662
rect 4220 82640 4516 82660
rect 19580 82172 19876 82192
rect 19636 82170 19660 82172
rect 19716 82170 19740 82172
rect 19796 82170 19820 82172
rect 19658 82118 19660 82170
rect 19722 82118 19734 82170
rect 19796 82118 19798 82170
rect 19636 82116 19660 82118
rect 19716 82116 19740 82118
rect 19796 82116 19820 82118
rect 19580 82096 19876 82116
rect 4220 81628 4516 81648
rect 4276 81626 4300 81628
rect 4356 81626 4380 81628
rect 4436 81626 4460 81628
rect 4298 81574 4300 81626
rect 4362 81574 4374 81626
rect 4436 81574 4438 81626
rect 4276 81572 4300 81574
rect 4356 81572 4380 81574
rect 4436 81572 4460 81574
rect 4220 81552 4516 81572
rect 19580 81084 19876 81104
rect 19636 81082 19660 81084
rect 19716 81082 19740 81084
rect 19796 81082 19820 81084
rect 19658 81030 19660 81082
rect 19722 81030 19734 81082
rect 19796 81030 19798 81082
rect 19636 81028 19660 81030
rect 19716 81028 19740 81030
rect 19796 81028 19820 81030
rect 19580 81008 19876 81028
rect 4220 80540 4516 80560
rect 4276 80538 4300 80540
rect 4356 80538 4380 80540
rect 4436 80538 4460 80540
rect 4298 80486 4300 80538
rect 4362 80486 4374 80538
rect 4436 80486 4438 80538
rect 4276 80484 4300 80486
rect 4356 80484 4380 80486
rect 4436 80484 4460 80486
rect 4220 80464 4516 80484
rect 19580 79996 19876 80016
rect 19636 79994 19660 79996
rect 19716 79994 19740 79996
rect 19796 79994 19820 79996
rect 19658 79942 19660 79994
rect 19722 79942 19734 79994
rect 19796 79942 19798 79994
rect 19636 79940 19660 79942
rect 19716 79940 19740 79942
rect 19796 79940 19820 79942
rect 19580 79920 19876 79940
rect 4220 79452 4516 79472
rect 4276 79450 4300 79452
rect 4356 79450 4380 79452
rect 4436 79450 4460 79452
rect 4298 79398 4300 79450
rect 4362 79398 4374 79450
rect 4436 79398 4438 79450
rect 4276 79396 4300 79398
rect 4356 79396 4380 79398
rect 4436 79396 4460 79398
rect 4220 79376 4516 79396
rect 19580 78908 19876 78928
rect 19636 78906 19660 78908
rect 19716 78906 19740 78908
rect 19796 78906 19820 78908
rect 19658 78854 19660 78906
rect 19722 78854 19734 78906
rect 19796 78854 19798 78906
rect 19636 78852 19660 78854
rect 19716 78852 19740 78854
rect 19796 78852 19820 78854
rect 19580 78832 19876 78852
rect 4220 78364 4516 78384
rect 4276 78362 4300 78364
rect 4356 78362 4380 78364
rect 4436 78362 4460 78364
rect 4298 78310 4300 78362
rect 4362 78310 4374 78362
rect 4436 78310 4438 78362
rect 4276 78308 4300 78310
rect 4356 78308 4380 78310
rect 4436 78308 4460 78310
rect 4220 78288 4516 78308
rect 19580 77820 19876 77840
rect 19636 77818 19660 77820
rect 19716 77818 19740 77820
rect 19796 77818 19820 77820
rect 19658 77766 19660 77818
rect 19722 77766 19734 77818
rect 19796 77766 19798 77818
rect 19636 77764 19660 77766
rect 19716 77764 19740 77766
rect 19796 77764 19820 77766
rect 19580 77744 19876 77764
rect 4220 77276 4516 77296
rect 4276 77274 4300 77276
rect 4356 77274 4380 77276
rect 4436 77274 4460 77276
rect 4298 77222 4300 77274
rect 4362 77222 4374 77274
rect 4436 77222 4438 77274
rect 4276 77220 4300 77222
rect 4356 77220 4380 77222
rect 4436 77220 4460 77222
rect 4220 77200 4516 77220
rect 19580 76732 19876 76752
rect 19636 76730 19660 76732
rect 19716 76730 19740 76732
rect 19796 76730 19820 76732
rect 19658 76678 19660 76730
rect 19722 76678 19734 76730
rect 19796 76678 19798 76730
rect 19636 76676 19660 76678
rect 19716 76676 19740 76678
rect 19796 76676 19820 76678
rect 19580 76656 19876 76676
rect 4220 76188 4516 76208
rect 4276 76186 4300 76188
rect 4356 76186 4380 76188
rect 4436 76186 4460 76188
rect 4298 76134 4300 76186
rect 4362 76134 4374 76186
rect 4436 76134 4438 76186
rect 4276 76132 4300 76134
rect 4356 76132 4380 76134
rect 4436 76132 4460 76134
rect 4220 76112 4516 76132
rect 19580 75644 19876 75664
rect 19636 75642 19660 75644
rect 19716 75642 19740 75644
rect 19796 75642 19820 75644
rect 19658 75590 19660 75642
rect 19722 75590 19734 75642
rect 19796 75590 19798 75642
rect 19636 75588 19660 75590
rect 19716 75588 19740 75590
rect 19796 75588 19820 75590
rect 19580 75568 19876 75588
rect 4220 75100 4516 75120
rect 4276 75098 4300 75100
rect 4356 75098 4380 75100
rect 4436 75098 4460 75100
rect 4298 75046 4300 75098
rect 4362 75046 4374 75098
rect 4436 75046 4438 75098
rect 4276 75044 4300 75046
rect 4356 75044 4380 75046
rect 4436 75044 4460 75046
rect 4220 75024 4516 75044
rect 19580 74556 19876 74576
rect 19636 74554 19660 74556
rect 19716 74554 19740 74556
rect 19796 74554 19820 74556
rect 19658 74502 19660 74554
rect 19722 74502 19734 74554
rect 19796 74502 19798 74554
rect 19636 74500 19660 74502
rect 19716 74500 19740 74502
rect 19796 74500 19820 74502
rect 19580 74480 19876 74500
rect 4220 74012 4516 74032
rect 4276 74010 4300 74012
rect 4356 74010 4380 74012
rect 4436 74010 4460 74012
rect 4298 73958 4300 74010
rect 4362 73958 4374 74010
rect 4436 73958 4438 74010
rect 4276 73956 4300 73958
rect 4356 73956 4380 73958
rect 4436 73956 4460 73958
rect 4220 73936 4516 73956
rect 19580 73468 19876 73488
rect 19636 73466 19660 73468
rect 19716 73466 19740 73468
rect 19796 73466 19820 73468
rect 19658 73414 19660 73466
rect 19722 73414 19734 73466
rect 19796 73414 19798 73466
rect 19636 73412 19660 73414
rect 19716 73412 19740 73414
rect 19796 73412 19820 73414
rect 19580 73392 19876 73412
rect 4220 72924 4516 72944
rect 4276 72922 4300 72924
rect 4356 72922 4380 72924
rect 4436 72922 4460 72924
rect 4298 72870 4300 72922
rect 4362 72870 4374 72922
rect 4436 72870 4438 72922
rect 4276 72868 4300 72870
rect 4356 72868 4380 72870
rect 4436 72868 4460 72870
rect 4220 72848 4516 72868
rect 19580 72380 19876 72400
rect 19636 72378 19660 72380
rect 19716 72378 19740 72380
rect 19796 72378 19820 72380
rect 19658 72326 19660 72378
rect 19722 72326 19734 72378
rect 19796 72326 19798 72378
rect 19636 72324 19660 72326
rect 19716 72324 19740 72326
rect 19796 72324 19820 72326
rect 19580 72304 19876 72324
rect 4220 71836 4516 71856
rect 4276 71834 4300 71836
rect 4356 71834 4380 71836
rect 4436 71834 4460 71836
rect 4298 71782 4300 71834
rect 4362 71782 4374 71834
rect 4436 71782 4438 71834
rect 4276 71780 4300 71782
rect 4356 71780 4380 71782
rect 4436 71780 4460 71782
rect 4220 71760 4516 71780
rect 19580 71292 19876 71312
rect 19636 71290 19660 71292
rect 19716 71290 19740 71292
rect 19796 71290 19820 71292
rect 19658 71238 19660 71290
rect 19722 71238 19734 71290
rect 19796 71238 19798 71290
rect 19636 71236 19660 71238
rect 19716 71236 19740 71238
rect 19796 71236 19820 71238
rect 19580 71216 19876 71236
rect 4220 70748 4516 70768
rect 4276 70746 4300 70748
rect 4356 70746 4380 70748
rect 4436 70746 4460 70748
rect 4298 70694 4300 70746
rect 4362 70694 4374 70746
rect 4436 70694 4438 70746
rect 4276 70692 4300 70694
rect 4356 70692 4380 70694
rect 4436 70692 4460 70694
rect 4220 70672 4516 70692
rect 19580 70204 19876 70224
rect 19636 70202 19660 70204
rect 19716 70202 19740 70204
rect 19796 70202 19820 70204
rect 19658 70150 19660 70202
rect 19722 70150 19734 70202
rect 19796 70150 19798 70202
rect 19636 70148 19660 70150
rect 19716 70148 19740 70150
rect 19796 70148 19820 70150
rect 19580 70128 19876 70148
rect 4220 69660 4516 69680
rect 4276 69658 4300 69660
rect 4356 69658 4380 69660
rect 4436 69658 4460 69660
rect 4298 69606 4300 69658
rect 4362 69606 4374 69658
rect 4436 69606 4438 69658
rect 4276 69604 4300 69606
rect 4356 69604 4380 69606
rect 4436 69604 4460 69606
rect 4220 69584 4516 69604
rect 19580 69116 19876 69136
rect 19636 69114 19660 69116
rect 19716 69114 19740 69116
rect 19796 69114 19820 69116
rect 19658 69062 19660 69114
rect 19722 69062 19734 69114
rect 19796 69062 19798 69114
rect 19636 69060 19660 69062
rect 19716 69060 19740 69062
rect 19796 69060 19820 69062
rect 19580 69040 19876 69060
rect 4220 68572 4516 68592
rect 4276 68570 4300 68572
rect 4356 68570 4380 68572
rect 4436 68570 4460 68572
rect 4298 68518 4300 68570
rect 4362 68518 4374 68570
rect 4436 68518 4438 68570
rect 4276 68516 4300 68518
rect 4356 68516 4380 68518
rect 4436 68516 4460 68518
rect 4220 68496 4516 68516
rect 19580 68028 19876 68048
rect 19636 68026 19660 68028
rect 19716 68026 19740 68028
rect 19796 68026 19820 68028
rect 19658 67974 19660 68026
rect 19722 67974 19734 68026
rect 19796 67974 19798 68026
rect 19636 67972 19660 67974
rect 19716 67972 19740 67974
rect 19796 67972 19820 67974
rect 19580 67952 19876 67972
rect 4220 67484 4516 67504
rect 4276 67482 4300 67484
rect 4356 67482 4380 67484
rect 4436 67482 4460 67484
rect 4298 67430 4300 67482
rect 4362 67430 4374 67482
rect 4436 67430 4438 67482
rect 4276 67428 4300 67430
rect 4356 67428 4380 67430
rect 4436 67428 4460 67430
rect 4220 67408 4516 67428
rect 19580 66940 19876 66960
rect 19636 66938 19660 66940
rect 19716 66938 19740 66940
rect 19796 66938 19820 66940
rect 19658 66886 19660 66938
rect 19722 66886 19734 66938
rect 19796 66886 19798 66938
rect 19636 66884 19660 66886
rect 19716 66884 19740 66886
rect 19796 66884 19820 66886
rect 19580 66864 19876 66884
rect 4220 66396 4516 66416
rect 4276 66394 4300 66396
rect 4356 66394 4380 66396
rect 4436 66394 4460 66396
rect 4298 66342 4300 66394
rect 4362 66342 4374 66394
rect 4436 66342 4438 66394
rect 4276 66340 4300 66342
rect 4356 66340 4380 66342
rect 4436 66340 4460 66342
rect 4220 66320 4516 66340
rect 19580 65852 19876 65872
rect 19636 65850 19660 65852
rect 19716 65850 19740 65852
rect 19796 65850 19820 65852
rect 19658 65798 19660 65850
rect 19722 65798 19734 65850
rect 19796 65798 19798 65850
rect 19636 65796 19660 65798
rect 19716 65796 19740 65798
rect 19796 65796 19820 65798
rect 19580 65776 19876 65796
rect 4220 65308 4516 65328
rect 4276 65306 4300 65308
rect 4356 65306 4380 65308
rect 4436 65306 4460 65308
rect 4298 65254 4300 65306
rect 4362 65254 4374 65306
rect 4436 65254 4438 65306
rect 4276 65252 4300 65254
rect 4356 65252 4380 65254
rect 4436 65252 4460 65254
rect 4220 65232 4516 65252
rect 19580 64764 19876 64784
rect 19636 64762 19660 64764
rect 19716 64762 19740 64764
rect 19796 64762 19820 64764
rect 19658 64710 19660 64762
rect 19722 64710 19734 64762
rect 19796 64710 19798 64762
rect 19636 64708 19660 64710
rect 19716 64708 19740 64710
rect 19796 64708 19820 64710
rect 19580 64688 19876 64708
rect 4220 64220 4516 64240
rect 4276 64218 4300 64220
rect 4356 64218 4380 64220
rect 4436 64218 4460 64220
rect 4298 64166 4300 64218
rect 4362 64166 4374 64218
rect 4436 64166 4438 64218
rect 4276 64164 4300 64166
rect 4356 64164 4380 64166
rect 4436 64164 4460 64166
rect 4220 64144 4516 64164
rect 19580 63676 19876 63696
rect 19636 63674 19660 63676
rect 19716 63674 19740 63676
rect 19796 63674 19820 63676
rect 19658 63622 19660 63674
rect 19722 63622 19734 63674
rect 19796 63622 19798 63674
rect 19636 63620 19660 63622
rect 19716 63620 19740 63622
rect 19796 63620 19820 63622
rect 19580 63600 19876 63620
rect 4220 63132 4516 63152
rect 4276 63130 4300 63132
rect 4356 63130 4380 63132
rect 4436 63130 4460 63132
rect 4298 63078 4300 63130
rect 4362 63078 4374 63130
rect 4436 63078 4438 63130
rect 4276 63076 4300 63078
rect 4356 63076 4380 63078
rect 4436 63076 4460 63078
rect 4220 63056 4516 63076
rect 19580 62588 19876 62608
rect 19636 62586 19660 62588
rect 19716 62586 19740 62588
rect 19796 62586 19820 62588
rect 19658 62534 19660 62586
rect 19722 62534 19734 62586
rect 19796 62534 19798 62586
rect 19636 62532 19660 62534
rect 19716 62532 19740 62534
rect 19796 62532 19820 62534
rect 19580 62512 19876 62532
rect 4220 62044 4516 62064
rect 4276 62042 4300 62044
rect 4356 62042 4380 62044
rect 4436 62042 4460 62044
rect 4298 61990 4300 62042
rect 4362 61990 4374 62042
rect 4436 61990 4438 62042
rect 4276 61988 4300 61990
rect 4356 61988 4380 61990
rect 4436 61988 4460 61990
rect 4220 61968 4516 61988
rect 19580 61500 19876 61520
rect 19636 61498 19660 61500
rect 19716 61498 19740 61500
rect 19796 61498 19820 61500
rect 19658 61446 19660 61498
rect 19722 61446 19734 61498
rect 19796 61446 19798 61498
rect 19636 61444 19660 61446
rect 19716 61444 19740 61446
rect 19796 61444 19820 61446
rect 19580 61424 19876 61444
rect 4220 60956 4516 60976
rect 4276 60954 4300 60956
rect 4356 60954 4380 60956
rect 4436 60954 4460 60956
rect 4298 60902 4300 60954
rect 4362 60902 4374 60954
rect 4436 60902 4438 60954
rect 4276 60900 4300 60902
rect 4356 60900 4380 60902
rect 4436 60900 4460 60902
rect 4220 60880 4516 60900
rect 19580 60412 19876 60432
rect 19636 60410 19660 60412
rect 19716 60410 19740 60412
rect 19796 60410 19820 60412
rect 19658 60358 19660 60410
rect 19722 60358 19734 60410
rect 19796 60358 19798 60410
rect 19636 60356 19660 60358
rect 19716 60356 19740 60358
rect 19796 60356 19820 60358
rect 19580 60336 19876 60356
rect 3056 60172 3108 60178
rect 3056 60114 3108 60120
rect 2042 60072 2098 60081
rect 2042 60007 2044 60016
rect 2096 60007 2098 60016
rect 2044 59978 2096 59984
rect 3068 59770 3096 60114
rect 4220 59868 4516 59888
rect 4276 59866 4300 59868
rect 4356 59866 4380 59868
rect 4436 59866 4460 59868
rect 4298 59814 4300 59866
rect 4362 59814 4374 59866
rect 4436 59814 4438 59866
rect 4276 59812 4300 59814
rect 4356 59812 4380 59814
rect 4436 59812 4460 59814
rect 4220 59792 4516 59812
rect 3056 59764 3108 59770
rect 3056 59706 3108 59712
rect 19580 59324 19876 59344
rect 19636 59322 19660 59324
rect 19716 59322 19740 59324
rect 19796 59322 19820 59324
rect 19658 59270 19660 59322
rect 19722 59270 19734 59322
rect 19796 59270 19798 59322
rect 19636 59268 19660 59270
rect 19716 59268 19740 59270
rect 19796 59268 19820 59270
rect 19580 59248 19876 59268
rect 4220 58780 4516 58800
rect 4276 58778 4300 58780
rect 4356 58778 4380 58780
rect 4436 58778 4460 58780
rect 4298 58726 4300 58778
rect 4362 58726 4374 58778
rect 4436 58726 4438 58778
rect 4276 58724 4300 58726
rect 4356 58724 4380 58726
rect 4436 58724 4460 58726
rect 4220 58704 4516 58724
rect 19580 58236 19876 58256
rect 19636 58234 19660 58236
rect 19716 58234 19740 58236
rect 19796 58234 19820 58236
rect 19658 58182 19660 58234
rect 19722 58182 19734 58234
rect 19796 58182 19798 58234
rect 19636 58180 19660 58182
rect 19716 58180 19740 58182
rect 19796 58180 19820 58182
rect 19580 58160 19876 58180
rect 4220 57692 4516 57712
rect 4276 57690 4300 57692
rect 4356 57690 4380 57692
rect 4436 57690 4460 57692
rect 4298 57638 4300 57690
rect 4362 57638 4374 57690
rect 4436 57638 4438 57690
rect 4276 57636 4300 57638
rect 4356 57636 4380 57638
rect 4436 57636 4460 57638
rect 4220 57616 4516 57636
rect 19580 57148 19876 57168
rect 19636 57146 19660 57148
rect 19716 57146 19740 57148
rect 19796 57146 19820 57148
rect 19658 57094 19660 57146
rect 19722 57094 19734 57146
rect 19796 57094 19798 57146
rect 19636 57092 19660 57094
rect 19716 57092 19740 57094
rect 19796 57092 19820 57094
rect 19580 57072 19876 57092
rect 4220 56604 4516 56624
rect 4276 56602 4300 56604
rect 4356 56602 4380 56604
rect 4436 56602 4460 56604
rect 4298 56550 4300 56602
rect 4362 56550 4374 56602
rect 4436 56550 4438 56602
rect 4276 56548 4300 56550
rect 4356 56548 4380 56550
rect 4436 56548 4460 56550
rect 4220 56528 4516 56548
rect 19580 56060 19876 56080
rect 19636 56058 19660 56060
rect 19716 56058 19740 56060
rect 19796 56058 19820 56060
rect 19658 56006 19660 56058
rect 19722 56006 19734 56058
rect 19796 56006 19798 56058
rect 19636 56004 19660 56006
rect 19716 56004 19740 56006
rect 19796 56004 19820 56006
rect 19580 55984 19876 56004
rect 4220 55516 4516 55536
rect 4276 55514 4300 55516
rect 4356 55514 4380 55516
rect 4436 55514 4460 55516
rect 4298 55462 4300 55514
rect 4362 55462 4374 55514
rect 4436 55462 4438 55514
rect 4276 55460 4300 55462
rect 4356 55460 4380 55462
rect 4436 55460 4460 55462
rect 4220 55440 4516 55460
rect 19580 54972 19876 54992
rect 19636 54970 19660 54972
rect 19716 54970 19740 54972
rect 19796 54970 19820 54972
rect 19658 54918 19660 54970
rect 19722 54918 19734 54970
rect 19796 54918 19798 54970
rect 19636 54916 19660 54918
rect 19716 54916 19740 54918
rect 19796 54916 19820 54918
rect 19580 54896 19876 54916
rect 4220 54428 4516 54448
rect 4276 54426 4300 54428
rect 4356 54426 4380 54428
rect 4436 54426 4460 54428
rect 4298 54374 4300 54426
rect 4362 54374 4374 54426
rect 4436 54374 4438 54426
rect 4276 54372 4300 54374
rect 4356 54372 4380 54374
rect 4436 54372 4460 54374
rect 4220 54352 4516 54372
rect 19580 53884 19876 53904
rect 19636 53882 19660 53884
rect 19716 53882 19740 53884
rect 19796 53882 19820 53884
rect 19658 53830 19660 53882
rect 19722 53830 19734 53882
rect 19796 53830 19798 53882
rect 19636 53828 19660 53830
rect 19716 53828 19740 53830
rect 19796 53828 19820 53830
rect 19580 53808 19876 53828
rect 4220 53340 4516 53360
rect 4276 53338 4300 53340
rect 4356 53338 4380 53340
rect 4436 53338 4460 53340
rect 4298 53286 4300 53338
rect 4362 53286 4374 53338
rect 4436 53286 4438 53338
rect 4276 53284 4300 53286
rect 4356 53284 4380 53286
rect 4436 53284 4460 53286
rect 4220 53264 4516 53284
rect 19580 52796 19876 52816
rect 19636 52794 19660 52796
rect 19716 52794 19740 52796
rect 19796 52794 19820 52796
rect 19658 52742 19660 52794
rect 19722 52742 19734 52794
rect 19796 52742 19798 52794
rect 19636 52740 19660 52742
rect 19716 52740 19740 52742
rect 19796 52740 19820 52742
rect 19580 52720 19876 52740
rect 4220 52252 4516 52272
rect 4276 52250 4300 52252
rect 4356 52250 4380 52252
rect 4436 52250 4460 52252
rect 4298 52198 4300 52250
rect 4362 52198 4374 52250
rect 4436 52198 4438 52250
rect 4276 52196 4300 52198
rect 4356 52196 4380 52198
rect 4436 52196 4460 52198
rect 4220 52176 4516 52196
rect 19580 51708 19876 51728
rect 19636 51706 19660 51708
rect 19716 51706 19740 51708
rect 19796 51706 19820 51708
rect 19658 51654 19660 51706
rect 19722 51654 19734 51706
rect 19796 51654 19798 51706
rect 19636 51652 19660 51654
rect 19716 51652 19740 51654
rect 19796 51652 19820 51654
rect 19580 51632 19876 51652
rect 4220 51164 4516 51184
rect 4276 51162 4300 51164
rect 4356 51162 4380 51164
rect 4436 51162 4460 51164
rect 4298 51110 4300 51162
rect 4362 51110 4374 51162
rect 4436 51110 4438 51162
rect 4276 51108 4300 51110
rect 4356 51108 4380 51110
rect 4436 51108 4460 51110
rect 4220 51088 4516 51108
rect 19580 50620 19876 50640
rect 19636 50618 19660 50620
rect 19716 50618 19740 50620
rect 19796 50618 19820 50620
rect 19658 50566 19660 50618
rect 19722 50566 19734 50618
rect 19796 50566 19798 50618
rect 19636 50564 19660 50566
rect 19716 50564 19740 50566
rect 19796 50564 19820 50566
rect 19580 50544 19876 50564
rect 4220 50076 4516 50096
rect 4276 50074 4300 50076
rect 4356 50074 4380 50076
rect 4436 50074 4460 50076
rect 4298 50022 4300 50074
rect 4362 50022 4374 50074
rect 4436 50022 4438 50074
rect 4276 50020 4300 50022
rect 4356 50020 4380 50022
rect 4436 50020 4460 50022
rect 4220 50000 4516 50020
rect 19580 49532 19876 49552
rect 19636 49530 19660 49532
rect 19716 49530 19740 49532
rect 19796 49530 19820 49532
rect 19658 49478 19660 49530
rect 19722 49478 19734 49530
rect 19796 49478 19798 49530
rect 19636 49476 19660 49478
rect 19716 49476 19740 49478
rect 19796 49476 19820 49478
rect 19580 49456 19876 49476
rect 4220 48988 4516 49008
rect 4276 48986 4300 48988
rect 4356 48986 4380 48988
rect 4436 48986 4460 48988
rect 4298 48934 4300 48986
rect 4362 48934 4374 48986
rect 4436 48934 4438 48986
rect 4276 48932 4300 48934
rect 4356 48932 4380 48934
rect 4436 48932 4460 48934
rect 4220 48912 4516 48932
rect 19580 48444 19876 48464
rect 19636 48442 19660 48444
rect 19716 48442 19740 48444
rect 19796 48442 19820 48444
rect 19658 48390 19660 48442
rect 19722 48390 19734 48442
rect 19796 48390 19798 48442
rect 19636 48388 19660 48390
rect 19716 48388 19740 48390
rect 19796 48388 19820 48390
rect 19580 48368 19876 48388
rect 4220 47900 4516 47920
rect 4276 47898 4300 47900
rect 4356 47898 4380 47900
rect 4436 47898 4460 47900
rect 4298 47846 4300 47898
rect 4362 47846 4374 47898
rect 4436 47846 4438 47898
rect 4276 47844 4300 47846
rect 4356 47844 4380 47846
rect 4436 47844 4460 47846
rect 4220 47824 4516 47844
rect 19580 47356 19876 47376
rect 19636 47354 19660 47356
rect 19716 47354 19740 47356
rect 19796 47354 19820 47356
rect 19658 47302 19660 47354
rect 19722 47302 19734 47354
rect 19796 47302 19798 47354
rect 19636 47300 19660 47302
rect 19716 47300 19740 47302
rect 19796 47300 19820 47302
rect 19580 47280 19876 47300
rect 4220 46812 4516 46832
rect 4276 46810 4300 46812
rect 4356 46810 4380 46812
rect 4436 46810 4460 46812
rect 4298 46758 4300 46810
rect 4362 46758 4374 46810
rect 4436 46758 4438 46810
rect 4276 46756 4300 46758
rect 4356 46756 4380 46758
rect 4436 46756 4460 46758
rect 4220 46736 4516 46756
rect 19580 46268 19876 46288
rect 19636 46266 19660 46268
rect 19716 46266 19740 46268
rect 19796 46266 19820 46268
rect 19658 46214 19660 46266
rect 19722 46214 19734 46266
rect 19796 46214 19798 46266
rect 19636 46212 19660 46214
rect 19716 46212 19740 46214
rect 19796 46212 19820 46214
rect 19580 46192 19876 46212
rect 4220 45724 4516 45744
rect 4276 45722 4300 45724
rect 4356 45722 4380 45724
rect 4436 45722 4460 45724
rect 4298 45670 4300 45722
rect 4362 45670 4374 45722
rect 4436 45670 4438 45722
rect 4276 45668 4300 45670
rect 4356 45668 4380 45670
rect 4436 45668 4460 45670
rect 4220 45648 4516 45668
rect 19580 45180 19876 45200
rect 19636 45178 19660 45180
rect 19716 45178 19740 45180
rect 19796 45178 19820 45180
rect 19658 45126 19660 45178
rect 19722 45126 19734 45178
rect 19796 45126 19798 45178
rect 19636 45124 19660 45126
rect 19716 45124 19740 45126
rect 19796 45124 19820 45126
rect 19580 45104 19876 45124
rect 4220 44636 4516 44656
rect 4276 44634 4300 44636
rect 4356 44634 4380 44636
rect 4436 44634 4460 44636
rect 4298 44582 4300 44634
rect 4362 44582 4374 44634
rect 4436 44582 4438 44634
rect 4276 44580 4300 44582
rect 4356 44580 4380 44582
rect 4436 44580 4460 44582
rect 4220 44560 4516 44580
rect 19580 44092 19876 44112
rect 19636 44090 19660 44092
rect 19716 44090 19740 44092
rect 19796 44090 19820 44092
rect 19658 44038 19660 44090
rect 19722 44038 19734 44090
rect 19796 44038 19798 44090
rect 19636 44036 19660 44038
rect 19716 44036 19740 44038
rect 19796 44036 19820 44038
rect 19580 44016 19876 44036
rect 4220 43548 4516 43568
rect 4276 43546 4300 43548
rect 4356 43546 4380 43548
rect 4436 43546 4460 43548
rect 4298 43494 4300 43546
rect 4362 43494 4374 43546
rect 4436 43494 4438 43546
rect 4276 43492 4300 43494
rect 4356 43492 4380 43494
rect 4436 43492 4460 43494
rect 4220 43472 4516 43492
rect 19580 43004 19876 43024
rect 19636 43002 19660 43004
rect 19716 43002 19740 43004
rect 19796 43002 19820 43004
rect 19658 42950 19660 43002
rect 19722 42950 19734 43002
rect 19796 42950 19798 43002
rect 19636 42948 19660 42950
rect 19716 42948 19740 42950
rect 19796 42948 19820 42950
rect 19580 42928 19876 42948
rect 4220 42460 4516 42480
rect 4276 42458 4300 42460
rect 4356 42458 4380 42460
rect 4436 42458 4460 42460
rect 4298 42406 4300 42458
rect 4362 42406 4374 42458
rect 4436 42406 4438 42458
rect 4276 42404 4300 42406
rect 4356 42404 4380 42406
rect 4436 42404 4460 42406
rect 4220 42384 4516 42404
rect 19580 41916 19876 41936
rect 19636 41914 19660 41916
rect 19716 41914 19740 41916
rect 19796 41914 19820 41916
rect 19658 41862 19660 41914
rect 19722 41862 19734 41914
rect 19796 41862 19798 41914
rect 19636 41860 19660 41862
rect 19716 41860 19740 41862
rect 19796 41860 19820 41862
rect 19580 41840 19876 41860
rect 4220 41372 4516 41392
rect 4276 41370 4300 41372
rect 4356 41370 4380 41372
rect 4436 41370 4460 41372
rect 4298 41318 4300 41370
rect 4362 41318 4374 41370
rect 4436 41318 4438 41370
rect 4276 41316 4300 41318
rect 4356 41316 4380 41318
rect 4436 41316 4460 41318
rect 4220 41296 4516 41316
rect 19580 40828 19876 40848
rect 19636 40826 19660 40828
rect 19716 40826 19740 40828
rect 19796 40826 19820 40828
rect 19658 40774 19660 40826
rect 19722 40774 19734 40826
rect 19796 40774 19798 40826
rect 19636 40772 19660 40774
rect 19716 40772 19740 40774
rect 19796 40772 19820 40774
rect 19580 40752 19876 40772
rect 4220 40284 4516 40304
rect 4276 40282 4300 40284
rect 4356 40282 4380 40284
rect 4436 40282 4460 40284
rect 4298 40230 4300 40282
rect 4362 40230 4374 40282
rect 4436 40230 4438 40282
rect 4276 40228 4300 40230
rect 4356 40228 4380 40230
rect 4436 40228 4460 40230
rect 4220 40208 4516 40228
rect 19580 39740 19876 39760
rect 19636 39738 19660 39740
rect 19716 39738 19740 39740
rect 19796 39738 19820 39740
rect 19658 39686 19660 39738
rect 19722 39686 19734 39738
rect 19796 39686 19798 39738
rect 19636 39684 19660 39686
rect 19716 39684 19740 39686
rect 19796 39684 19820 39686
rect 19580 39664 19876 39684
rect 4220 39196 4516 39216
rect 4276 39194 4300 39196
rect 4356 39194 4380 39196
rect 4436 39194 4460 39196
rect 4298 39142 4300 39194
rect 4362 39142 4374 39194
rect 4436 39142 4438 39194
rect 4276 39140 4300 39142
rect 4356 39140 4380 39142
rect 4436 39140 4460 39142
rect 4220 39120 4516 39140
rect 19580 38652 19876 38672
rect 19636 38650 19660 38652
rect 19716 38650 19740 38652
rect 19796 38650 19820 38652
rect 19658 38598 19660 38650
rect 19722 38598 19734 38650
rect 19796 38598 19798 38650
rect 19636 38596 19660 38598
rect 19716 38596 19740 38598
rect 19796 38596 19820 38598
rect 19580 38576 19876 38596
rect 4220 38108 4516 38128
rect 4276 38106 4300 38108
rect 4356 38106 4380 38108
rect 4436 38106 4460 38108
rect 4298 38054 4300 38106
rect 4362 38054 4374 38106
rect 4436 38054 4438 38106
rect 4276 38052 4300 38054
rect 4356 38052 4380 38054
rect 4436 38052 4460 38054
rect 4220 38032 4516 38052
rect 19580 37564 19876 37584
rect 19636 37562 19660 37564
rect 19716 37562 19740 37564
rect 19796 37562 19820 37564
rect 19658 37510 19660 37562
rect 19722 37510 19734 37562
rect 19796 37510 19798 37562
rect 19636 37508 19660 37510
rect 19716 37508 19740 37510
rect 19796 37508 19820 37510
rect 19580 37488 19876 37508
rect 4220 37020 4516 37040
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4298 36966 4300 37018
rect 4362 36966 4374 37018
rect 4436 36966 4438 37018
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4220 36944 4516 36964
rect 19580 36476 19876 36496
rect 19636 36474 19660 36476
rect 19716 36474 19740 36476
rect 19796 36474 19820 36476
rect 19658 36422 19660 36474
rect 19722 36422 19734 36474
rect 19796 36422 19798 36474
rect 19636 36420 19660 36422
rect 19716 36420 19740 36422
rect 19796 36420 19820 36422
rect 19580 36400 19876 36420
rect 4220 35932 4516 35952
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4298 35878 4300 35930
rect 4362 35878 4374 35930
rect 4436 35878 4438 35930
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4220 35856 4516 35876
rect 19580 35388 19876 35408
rect 19636 35386 19660 35388
rect 19716 35386 19740 35388
rect 19796 35386 19820 35388
rect 19658 35334 19660 35386
rect 19722 35334 19734 35386
rect 19796 35334 19798 35386
rect 19636 35332 19660 35334
rect 19716 35332 19740 35334
rect 19796 35332 19820 35334
rect 19580 35312 19876 35332
rect 4220 34844 4516 34864
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4298 34790 4300 34842
rect 4362 34790 4374 34842
rect 4436 34790 4438 34842
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4220 34768 4516 34788
rect 19580 34300 19876 34320
rect 19636 34298 19660 34300
rect 19716 34298 19740 34300
rect 19796 34298 19820 34300
rect 19658 34246 19660 34298
rect 19722 34246 19734 34298
rect 19796 34246 19798 34298
rect 19636 34244 19660 34246
rect 19716 34244 19740 34246
rect 19796 34244 19820 34246
rect 19580 34224 19876 34244
rect 4220 33756 4516 33776
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4298 33702 4300 33754
rect 4362 33702 4374 33754
rect 4436 33702 4438 33754
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4220 33680 4516 33700
rect 19580 33212 19876 33232
rect 19636 33210 19660 33212
rect 19716 33210 19740 33212
rect 19796 33210 19820 33212
rect 19658 33158 19660 33210
rect 19722 33158 19734 33210
rect 19796 33158 19798 33210
rect 19636 33156 19660 33158
rect 19716 33156 19740 33158
rect 19796 33156 19820 33158
rect 19580 33136 19876 33156
rect 4220 32668 4516 32688
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4298 32614 4300 32666
rect 4362 32614 4374 32666
rect 4436 32614 4438 32666
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4220 32592 4516 32612
rect 19580 32124 19876 32144
rect 19636 32122 19660 32124
rect 19716 32122 19740 32124
rect 19796 32122 19820 32124
rect 19658 32070 19660 32122
rect 19722 32070 19734 32122
rect 19796 32070 19798 32122
rect 19636 32068 19660 32070
rect 19716 32068 19740 32070
rect 19796 32068 19820 32070
rect 19580 32048 19876 32068
rect 4220 31580 4516 31600
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4298 31526 4300 31578
rect 4362 31526 4374 31578
rect 4436 31526 4438 31578
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4220 31504 4516 31524
rect 19580 31036 19876 31056
rect 19636 31034 19660 31036
rect 19716 31034 19740 31036
rect 19796 31034 19820 31036
rect 19658 30982 19660 31034
rect 19722 30982 19734 31034
rect 19796 30982 19798 31034
rect 19636 30980 19660 30982
rect 19716 30980 19740 30982
rect 19796 30980 19820 30982
rect 19580 30960 19876 30980
rect 4220 30492 4516 30512
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4298 30438 4300 30490
rect 4362 30438 4374 30490
rect 4436 30438 4438 30490
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4220 30416 4516 30436
rect 19580 29948 19876 29968
rect 19636 29946 19660 29948
rect 19716 29946 19740 29948
rect 19796 29946 19820 29948
rect 19658 29894 19660 29946
rect 19722 29894 19734 29946
rect 19796 29894 19798 29946
rect 19636 29892 19660 29894
rect 19716 29892 19740 29894
rect 19796 29892 19820 29894
rect 19580 29872 19876 29892
rect 4220 29404 4516 29424
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4298 29350 4300 29402
rect 4362 29350 4374 29402
rect 4436 29350 4438 29402
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4220 29328 4516 29348
rect 19580 28860 19876 28880
rect 19636 28858 19660 28860
rect 19716 28858 19740 28860
rect 19796 28858 19820 28860
rect 19658 28806 19660 28858
rect 19722 28806 19734 28858
rect 19796 28806 19798 28858
rect 19636 28804 19660 28806
rect 19716 28804 19740 28806
rect 19796 28804 19820 28806
rect 19580 28784 19876 28804
rect 4220 28316 4516 28336
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4298 28262 4300 28314
rect 4362 28262 4374 28314
rect 4436 28262 4438 28314
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4220 28240 4516 28260
rect 19580 27772 19876 27792
rect 19636 27770 19660 27772
rect 19716 27770 19740 27772
rect 19796 27770 19820 27772
rect 19658 27718 19660 27770
rect 19722 27718 19734 27770
rect 19796 27718 19798 27770
rect 19636 27716 19660 27718
rect 19716 27716 19740 27718
rect 19796 27716 19820 27718
rect 19580 27696 19876 27716
rect 4220 27228 4516 27248
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4298 27174 4300 27226
rect 4362 27174 4374 27226
rect 4436 27174 4438 27226
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4220 27152 4516 27172
rect 19580 26684 19876 26704
rect 19636 26682 19660 26684
rect 19716 26682 19740 26684
rect 19796 26682 19820 26684
rect 19658 26630 19660 26682
rect 19722 26630 19734 26682
rect 19796 26630 19798 26682
rect 19636 26628 19660 26630
rect 19716 26628 19740 26630
rect 19796 26628 19820 26630
rect 19580 26608 19876 26628
rect 4220 26140 4516 26160
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4298 26086 4300 26138
rect 4362 26086 4374 26138
rect 4436 26086 4438 26138
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4220 26064 4516 26084
rect 19580 25596 19876 25616
rect 19636 25594 19660 25596
rect 19716 25594 19740 25596
rect 19796 25594 19820 25596
rect 19658 25542 19660 25594
rect 19722 25542 19734 25594
rect 19796 25542 19798 25594
rect 19636 25540 19660 25542
rect 19716 25540 19740 25542
rect 19796 25540 19820 25542
rect 19580 25520 19876 25540
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 19580 24508 19876 24528
rect 19636 24506 19660 24508
rect 19716 24506 19740 24508
rect 19796 24506 19820 24508
rect 19658 24454 19660 24506
rect 19722 24454 19734 24506
rect 19796 24454 19798 24506
rect 19636 24452 19660 24454
rect 19716 24452 19740 24454
rect 19796 24452 19820 24454
rect 19580 24432 19876 24452
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 19580 23420 19876 23440
rect 19636 23418 19660 23420
rect 19716 23418 19740 23420
rect 19796 23418 19820 23420
rect 19658 23366 19660 23418
rect 19722 23366 19734 23418
rect 19796 23366 19798 23418
rect 19636 23364 19660 23366
rect 19716 23364 19740 23366
rect 19796 23364 19820 23366
rect 19580 23344 19876 23364
rect 26436 23186 26464 116690
rect 26528 116346 26556 117098
rect 29276 116884 29328 116890
rect 29276 116826 29328 116832
rect 29092 116816 29144 116822
rect 29092 116758 29144 116764
rect 26608 116612 26660 116618
rect 26608 116554 26660 116560
rect 26516 116340 26568 116346
rect 26516 116282 26568 116288
rect 26620 23186 26648 116554
rect 26424 23180 26476 23186
rect 26424 23122 26476 23128
rect 26608 23180 26660 23186
rect 26608 23122 26660 23128
rect 28264 23180 28316 23186
rect 28264 23122 28316 23128
rect 28172 23112 28224 23118
rect 28172 23054 28224 23060
rect 27988 22976 28040 22982
rect 27988 22918 28040 22924
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 19580 22332 19876 22352
rect 19636 22330 19660 22332
rect 19716 22330 19740 22332
rect 19796 22330 19820 22332
rect 19658 22278 19660 22330
rect 19722 22278 19734 22330
rect 19796 22278 19798 22330
rect 19636 22276 19660 22278
rect 19716 22276 19740 22278
rect 19796 22276 19820 22278
rect 19580 22256 19876 22276
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 28000 21486 28028 22918
rect 27988 21480 28040 21486
rect 27988 21422 28040 21428
rect 19580 21244 19876 21264
rect 19636 21242 19660 21244
rect 19716 21242 19740 21244
rect 19796 21242 19820 21244
rect 19658 21190 19660 21242
rect 19722 21190 19734 21242
rect 19796 21190 19798 21242
rect 19636 21188 19660 21190
rect 19716 21188 19740 21190
rect 19796 21188 19820 21190
rect 19580 21168 19876 21188
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 28000 20398 28028 21422
rect 28184 20466 28212 23054
rect 28172 20460 28224 20466
rect 28172 20402 28224 20408
rect 28276 20398 28304 23122
rect 29104 22166 29132 116758
rect 29288 26234 29316 116826
rect 30852 116346 30880 117098
rect 31024 116680 31076 116686
rect 31024 116622 31076 116628
rect 30840 116340 30892 116346
rect 30840 116282 30892 116288
rect 29196 26206 29316 26234
rect 29092 22160 29144 22166
rect 29092 22102 29144 22108
rect 29104 21078 29132 22102
rect 29196 21894 29224 26206
rect 31036 24274 31064 116622
rect 31760 116136 31812 116142
rect 31760 116078 31812 116084
rect 31024 24268 31076 24274
rect 31024 24210 31076 24216
rect 31392 24268 31444 24274
rect 31392 24210 31444 24216
rect 30380 22500 30432 22506
rect 30380 22442 30432 22448
rect 29276 22160 29328 22166
rect 29276 22102 29328 22108
rect 29184 21888 29236 21894
rect 29184 21830 29236 21836
rect 29092 21072 29144 21078
rect 29092 21014 29144 21020
rect 29196 21010 29224 21830
rect 29288 21350 29316 22102
rect 30392 21962 30420 22442
rect 30380 21956 30432 21962
rect 30380 21898 30432 21904
rect 29276 21344 29328 21350
rect 29276 21286 29328 21292
rect 29288 21010 29316 21286
rect 29184 21004 29236 21010
rect 29184 20946 29236 20952
rect 29276 21004 29328 21010
rect 29276 20946 29328 20952
rect 27988 20392 28040 20398
rect 27988 20334 28040 20340
rect 28264 20392 28316 20398
rect 28264 20334 28316 20340
rect 29092 20392 29144 20398
rect 29092 20334 29144 20340
rect 29000 20256 29052 20262
rect 29000 20198 29052 20204
rect 19580 20156 19876 20176
rect 19636 20154 19660 20156
rect 19716 20154 19740 20156
rect 19796 20154 19820 20156
rect 19658 20102 19660 20154
rect 19722 20102 19734 20154
rect 19796 20102 19798 20154
rect 19636 20100 19660 20102
rect 19716 20100 19740 20102
rect 19796 20100 19820 20102
rect 19580 20080 19876 20100
rect 28908 19712 28960 19718
rect 28908 19654 28960 19660
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 19580 19068 19876 19088
rect 19636 19066 19660 19068
rect 19716 19066 19740 19068
rect 19796 19066 19820 19068
rect 19658 19014 19660 19066
rect 19722 19014 19734 19066
rect 19796 19014 19798 19066
rect 19636 19012 19660 19014
rect 19716 19012 19740 19014
rect 19796 19012 19820 19014
rect 19580 18992 19876 19012
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 19580 17980 19876 18000
rect 19636 17978 19660 17980
rect 19716 17978 19740 17980
rect 19796 17978 19820 17980
rect 19658 17926 19660 17978
rect 19722 17926 19734 17978
rect 19796 17926 19798 17978
rect 19636 17924 19660 17926
rect 19716 17924 19740 17926
rect 19796 17924 19820 17926
rect 19580 17904 19876 17924
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 19580 16892 19876 16912
rect 19636 16890 19660 16892
rect 19716 16890 19740 16892
rect 19796 16890 19820 16892
rect 19658 16838 19660 16890
rect 19722 16838 19734 16890
rect 19796 16838 19798 16890
rect 19636 16836 19660 16838
rect 19716 16836 19740 16838
rect 19796 16836 19820 16838
rect 19580 16816 19876 16836
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 19580 15804 19876 15824
rect 19636 15802 19660 15804
rect 19716 15802 19740 15804
rect 19796 15802 19820 15804
rect 19658 15750 19660 15802
rect 19722 15750 19734 15802
rect 19796 15750 19798 15802
rect 19636 15748 19660 15750
rect 19716 15748 19740 15750
rect 19796 15748 19820 15750
rect 19580 15728 19876 15748
rect 28816 15360 28868 15366
rect 28816 15302 28868 15308
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 19580 14716 19876 14736
rect 19636 14714 19660 14716
rect 19716 14714 19740 14716
rect 19796 14714 19820 14716
rect 19658 14662 19660 14714
rect 19722 14662 19734 14714
rect 19796 14662 19798 14714
rect 19636 14660 19660 14662
rect 19716 14660 19740 14662
rect 19796 14660 19820 14662
rect 19580 14640 19876 14660
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 19580 13628 19876 13648
rect 19636 13626 19660 13628
rect 19716 13626 19740 13628
rect 19796 13626 19820 13628
rect 19658 13574 19660 13626
rect 19722 13574 19734 13626
rect 19796 13574 19798 13626
rect 19636 13572 19660 13574
rect 19716 13572 19740 13574
rect 19796 13572 19820 13574
rect 19580 13552 19876 13572
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 19580 12540 19876 12560
rect 19636 12538 19660 12540
rect 19716 12538 19740 12540
rect 19796 12538 19820 12540
rect 19658 12486 19660 12538
rect 19722 12486 19734 12538
rect 19796 12486 19798 12538
rect 19636 12484 19660 12486
rect 19716 12484 19740 12486
rect 19796 12484 19820 12486
rect 19580 12464 19876 12484
rect 28828 12434 28856 15302
rect 28920 15026 28948 19654
rect 29012 15706 29040 20198
rect 29000 15700 29052 15706
rect 29000 15642 29052 15648
rect 29104 15570 29132 20334
rect 29196 19922 29224 20946
rect 29288 20058 29316 20946
rect 29276 20052 29328 20058
rect 29276 19994 29328 20000
rect 30392 19922 30420 21898
rect 30656 20800 30708 20806
rect 30656 20742 30708 20748
rect 29184 19916 29236 19922
rect 29184 19858 29236 19864
rect 30380 19916 30432 19922
rect 30380 19858 30432 19864
rect 30668 18222 30696 20742
rect 31404 19922 31432 24210
rect 31208 19916 31260 19922
rect 31208 19858 31260 19864
rect 31392 19916 31444 19922
rect 31392 19858 31444 19864
rect 31024 19848 31076 19854
rect 31024 19790 31076 19796
rect 30656 18216 30708 18222
rect 30656 18158 30708 18164
rect 29092 15564 29144 15570
rect 29092 15506 29144 15512
rect 30012 15564 30064 15570
rect 30012 15506 30064 15512
rect 28908 15020 28960 15026
rect 28908 14962 28960 14968
rect 30024 14074 30052 15506
rect 31036 14822 31064 19790
rect 31220 18426 31248 19858
rect 31300 19712 31352 19718
rect 31300 19654 31352 19660
rect 31208 18420 31260 18426
rect 31208 18362 31260 18368
rect 31220 18222 31248 18362
rect 31312 18222 31340 19654
rect 31208 18216 31260 18222
rect 31208 18158 31260 18164
rect 31300 18216 31352 18222
rect 31300 18158 31352 18164
rect 31312 17746 31340 18158
rect 31300 17740 31352 17746
rect 31300 17682 31352 17688
rect 31208 15496 31260 15502
rect 31208 15438 31260 15444
rect 31220 15026 31248 15438
rect 31484 15360 31536 15366
rect 31484 15302 31536 15308
rect 31208 15020 31260 15026
rect 31208 14962 31260 14968
rect 31024 14816 31076 14822
rect 31024 14758 31076 14764
rect 31116 14476 31168 14482
rect 31116 14418 31168 14424
rect 30012 14068 30064 14074
rect 30012 14010 30064 14016
rect 30024 13954 30052 14010
rect 29932 13926 30052 13954
rect 30840 13932 30892 13938
rect 28828 12406 28948 12434
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 19580 11452 19876 11472
rect 19636 11450 19660 11452
rect 19716 11450 19740 11452
rect 19796 11450 19820 11452
rect 19658 11398 19660 11450
rect 19722 11398 19734 11450
rect 19796 11398 19798 11450
rect 19636 11396 19660 11398
rect 19716 11396 19740 11398
rect 19796 11396 19820 11398
rect 19580 11376 19876 11396
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 19580 10364 19876 10384
rect 19636 10362 19660 10364
rect 19716 10362 19740 10364
rect 19796 10362 19820 10364
rect 19658 10310 19660 10362
rect 19722 10310 19734 10362
rect 19796 10310 19798 10362
rect 19636 10308 19660 10310
rect 19716 10308 19740 10310
rect 19796 10308 19820 10310
rect 19580 10288 19876 10308
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 28920 9674 28948 12406
rect 28644 9646 28948 9674
rect 19580 9276 19876 9296
rect 19636 9274 19660 9276
rect 19716 9274 19740 9276
rect 19796 9274 19820 9276
rect 19658 9222 19660 9274
rect 19722 9222 19734 9274
rect 19796 9222 19798 9274
rect 19636 9220 19660 9222
rect 19716 9220 19740 9222
rect 19796 9220 19820 9222
rect 19580 9200 19876 9220
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 27804 8288 27856 8294
rect 27804 8230 27856 8236
rect 19580 8188 19876 8208
rect 19636 8186 19660 8188
rect 19716 8186 19740 8188
rect 19796 8186 19820 8188
rect 19658 8134 19660 8186
rect 19722 8134 19734 8186
rect 19796 8134 19798 8186
rect 19636 8132 19660 8134
rect 19716 8132 19740 8134
rect 19796 8132 19820 8134
rect 19580 8112 19876 8132
rect 27816 8022 27844 8230
rect 20996 8016 21048 8022
rect 20994 7984 20996 7993
rect 21272 8016 21324 8022
rect 21048 7984 21050 7993
rect 21272 7958 21324 7964
rect 24216 8016 24268 8022
rect 24216 7958 24268 7964
rect 27804 8016 27856 8022
rect 28172 8016 28224 8022
rect 27804 7958 27856 7964
rect 28170 7984 28172 7993
rect 28224 7984 28226 7993
rect 20994 7919 21050 7928
rect 21180 7948 21232 7954
rect 21180 7890 21232 7896
rect 20996 7880 21048 7886
rect 20996 7822 21048 7828
rect 20812 7744 20864 7750
rect 20812 7686 20864 7692
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 18604 7336 18656 7342
rect 18604 7278 18656 7284
rect 18972 7336 19024 7342
rect 18972 7278 19024 7284
rect 20168 7336 20220 7342
rect 20168 7278 20220 7284
rect 18052 7268 18104 7274
rect 18052 7210 18104 7216
rect 17960 7200 18012 7206
rect 17960 7142 18012 7148
rect 17972 6866 18000 7142
rect 17960 6860 18012 6866
rect 17960 6802 18012 6808
rect 18064 6746 18092 7210
rect 18616 6934 18644 7278
rect 18604 6928 18656 6934
rect 18604 6870 18656 6876
rect 18984 6866 19012 7278
rect 19580 7100 19876 7120
rect 19636 7098 19660 7100
rect 19716 7098 19740 7100
rect 19796 7098 19820 7100
rect 19658 7046 19660 7098
rect 19722 7046 19734 7098
rect 19796 7046 19798 7098
rect 19636 7044 19660 7046
rect 19716 7044 19740 7046
rect 19796 7044 19820 7046
rect 19580 7024 19876 7044
rect 20180 6866 20208 7278
rect 20444 7268 20496 7274
rect 20444 7210 20496 7216
rect 18696 6860 18748 6866
rect 18696 6802 18748 6808
rect 18972 6860 19024 6866
rect 18972 6802 19024 6808
rect 20168 6860 20220 6866
rect 20168 6802 20220 6808
rect 17408 6724 17460 6730
rect 17408 6666 17460 6672
rect 17972 6718 18092 6746
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 17316 6656 17368 6662
rect 17316 6598 17368 6604
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 17328 6254 17356 6598
rect 17316 6248 17368 6254
rect 17316 6190 17368 6196
rect 16580 6112 16632 6118
rect 16580 6054 16632 6060
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 1952 5364 2004 5370
rect 1952 5306 2004 5312
rect 1124 4072 1176 4078
rect 1124 4014 1176 4020
rect 1860 4072 1912 4078
rect 1860 4014 1912 4020
rect 756 3460 808 3466
rect 756 3402 808 3408
rect 388 2984 440 2990
rect 388 2926 440 2932
rect 112 2508 164 2514
rect 112 2450 164 2456
rect 124 800 152 2450
rect 400 800 428 2926
rect 768 800 796 3402
rect 1136 800 1164 4014
rect 1492 3528 1544 3534
rect 1492 3470 1544 3476
rect 1504 800 1532 3470
rect 1674 3088 1730 3097
rect 1674 3023 1676 3032
rect 1728 3023 1730 3032
rect 1676 2994 1728 3000
rect 1674 2544 1730 2553
rect 1674 2479 1676 2488
rect 1728 2479 1730 2488
rect 1676 2450 1728 2456
rect 1872 800 1900 4014
rect 1964 3670 1992 5306
rect 11796 4684 11848 4690
rect 11796 4626 11848 4632
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 5816 4276 5868 4282
rect 5816 4218 5868 4224
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 3160 3738 3188 4082
rect 3148 3732 3200 3738
rect 3148 3674 3200 3680
rect 1952 3664 2004 3670
rect 1952 3606 2004 3612
rect 3332 3596 3384 3602
rect 3332 3538 3384 3544
rect 4804 3596 4856 3602
rect 4804 3538 4856 3544
rect 2688 3392 2740 3398
rect 2688 3334 2740 3340
rect 2700 3194 2728 3334
rect 2688 3188 2740 3194
rect 2688 3130 2740 3136
rect 2228 2984 2280 2990
rect 2228 2926 2280 2932
rect 2240 800 2268 2926
rect 2964 2848 3016 2854
rect 2964 2790 3016 2796
rect 2596 2508 2648 2514
rect 2596 2450 2648 2456
rect 2608 800 2636 2450
rect 2780 2304 2832 2310
rect 2780 2246 2832 2252
rect 2792 1970 2820 2246
rect 2780 1964 2832 1970
rect 2780 1906 2832 1912
rect 2976 800 3004 2790
rect 3344 800 3372 3538
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 3700 2984 3752 2990
rect 3700 2926 3752 2932
rect 3712 800 3740 2926
rect 4620 2848 4672 2854
rect 4620 2790 4672 2796
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 4080 800 4108 2450
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 4632 1442 4660 2790
rect 4448 1414 4660 1442
rect 4448 800 4476 1414
rect 4816 800 4844 3538
rect 5172 2984 5224 2990
rect 5172 2926 5224 2932
rect 5184 800 5212 2926
rect 5828 2582 5856 4218
rect 10968 4072 11020 4078
rect 10968 4014 11020 4020
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 9968 3670 9996 3878
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 6276 3596 6328 3602
rect 6276 3538 6328 3544
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 5816 2576 5868 2582
rect 5816 2518 5868 2524
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 5552 800 5580 2450
rect 5908 2440 5960 2446
rect 5908 2382 5960 2388
rect 5920 800 5948 2382
rect 6288 800 6316 3538
rect 6644 2984 6696 2990
rect 6644 2926 6696 2932
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 9220 2984 9272 2990
rect 9220 2926 9272 2932
rect 6656 800 6684 2926
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 7024 800 7052 2450
rect 7196 2304 7248 2310
rect 7196 2246 7248 2252
rect 7208 1902 7236 2246
rect 7196 1896 7248 1902
rect 7196 1838 7248 1844
rect 7392 800 7420 2586
rect 7760 800 7788 2926
rect 8116 2508 8168 2514
rect 8116 2450 8168 2456
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 8128 800 8156 2450
rect 8496 800 8524 2450
rect 8576 2304 8628 2310
rect 8576 2246 8628 2252
rect 8852 2304 8904 2310
rect 8852 2246 8904 2252
rect 8588 2106 8616 2246
rect 8576 2100 8628 2106
rect 8576 2042 8628 2048
rect 8864 800 8892 2246
rect 9232 800 9260 2926
rect 9600 800 9628 3538
rect 9956 3120 10008 3126
rect 9956 3062 10008 3068
rect 9968 2938 9996 3062
rect 9876 2910 9996 2938
rect 10060 2922 10088 3878
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10140 3528 10192 3534
rect 10138 3496 10140 3505
rect 10192 3496 10194 3505
rect 10138 3431 10194 3440
rect 10048 2916 10100 2922
rect 9876 2854 9904 2910
rect 10048 2858 10100 2864
rect 9864 2848 9916 2854
rect 9864 2790 9916 2796
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 9692 2038 9720 2450
rect 9680 2032 9732 2038
rect 9680 1974 9732 1980
rect 9968 800 9996 2790
rect 10336 800 10364 3538
rect 10704 800 10732 3538
rect 10980 2922 11008 4014
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 11072 800 11100 2790
rect 11428 2508 11480 2514
rect 11428 2450 11480 2456
rect 11440 800 11468 2450
rect 11808 800 11836 4626
rect 14280 4548 14332 4554
rect 14280 4490 14332 4496
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 12072 4004 12124 4010
rect 12072 3946 12124 3952
rect 12256 4004 12308 4010
rect 12256 3946 12308 3952
rect 11886 3768 11942 3777
rect 11886 3703 11942 3712
rect 11900 3126 11928 3703
rect 11980 3392 12032 3398
rect 11980 3334 12032 3340
rect 11888 3120 11940 3126
rect 11992 3097 12020 3334
rect 11888 3062 11940 3068
rect 11978 3088 12034 3097
rect 11978 3023 12034 3032
rect 12084 2990 12112 3946
rect 12268 3670 12296 3946
rect 12360 3670 12388 4082
rect 12716 4072 12768 4078
rect 12438 4040 12494 4049
rect 12716 4014 12768 4020
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 12438 3975 12440 3984
rect 12492 3975 12494 3984
rect 12440 3946 12492 3952
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12636 3777 12664 3878
rect 12622 3768 12678 3777
rect 12622 3703 12678 3712
rect 12256 3664 12308 3670
rect 12256 3606 12308 3612
rect 12348 3664 12400 3670
rect 12348 3606 12400 3612
rect 12164 3392 12216 3398
rect 12164 3334 12216 3340
rect 12072 2984 12124 2990
rect 12072 2926 12124 2932
rect 12176 800 12204 3334
rect 12532 3120 12584 3126
rect 12530 3088 12532 3097
rect 12584 3088 12586 3097
rect 12530 3023 12586 3032
rect 12728 2774 12756 4014
rect 13360 3596 13412 3602
rect 13360 3538 13412 3544
rect 13084 3392 13136 3398
rect 13084 3334 13136 3340
rect 13096 2922 13124 3334
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 13084 2916 13136 2922
rect 13084 2858 13136 2864
rect 13188 2854 13216 3130
rect 13372 3058 13400 3538
rect 13360 3052 13412 3058
rect 13360 2994 13412 3000
rect 13176 2848 13228 2854
rect 13176 2790 13228 2796
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 12544 2746 12756 2774
rect 12544 800 12572 2746
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 12912 800 12940 2382
rect 13280 800 13308 2790
rect 13648 800 13676 4014
rect 13728 4004 13780 4010
rect 13728 3946 13780 3952
rect 13740 3670 13768 3946
rect 13728 3664 13780 3670
rect 13728 3606 13780 3612
rect 14292 2990 14320 4490
rect 14832 4140 14884 4146
rect 14832 4082 14884 4088
rect 14844 3670 14872 4082
rect 14832 3664 14884 3670
rect 14832 3606 14884 3612
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14372 3392 14424 3398
rect 14372 3334 14424 3340
rect 14004 2984 14056 2990
rect 14004 2926 14056 2932
rect 14280 2984 14332 2990
rect 14280 2926 14332 2932
rect 14016 800 14044 2926
rect 14384 800 14412 3334
rect 14752 800 14780 3470
rect 15200 3052 15252 3058
rect 15200 2994 15252 3000
rect 15212 2961 15240 2994
rect 15198 2952 15254 2961
rect 15198 2887 15254 2896
rect 15304 2774 15332 5850
rect 15660 5024 15712 5030
rect 15660 4966 15712 4972
rect 15672 4078 15700 4966
rect 15660 4072 15712 4078
rect 15660 4014 15712 4020
rect 15844 4072 15896 4078
rect 15844 4014 15896 4020
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 15660 3664 15712 3670
rect 15580 3624 15660 3652
rect 15384 3392 15436 3398
rect 15384 3334 15436 3340
rect 15396 3194 15424 3334
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 15304 2746 15424 2774
rect 15108 2508 15160 2514
rect 15108 2450 15160 2456
rect 15120 800 15148 2450
rect 15292 2304 15344 2310
rect 15292 2246 15344 2252
rect 15304 1086 15332 2246
rect 15396 2038 15424 2746
rect 15384 2032 15436 2038
rect 15384 1974 15436 1980
rect 15292 1080 15344 1086
rect 15292 1022 15344 1028
rect 15488 800 15516 3130
rect 15580 2854 15608 3624
rect 15660 3606 15712 3612
rect 15658 3496 15714 3505
rect 15658 3431 15714 3440
rect 15672 2990 15700 3431
rect 15660 2984 15712 2990
rect 15660 2926 15712 2932
rect 15568 2848 15620 2854
rect 15568 2790 15620 2796
rect 15856 800 15884 4014
rect 16224 2922 16252 4014
rect 16592 3602 16620 6054
rect 17328 5778 17356 6190
rect 17420 5914 17448 6666
rect 17972 6662 18000 6718
rect 17960 6656 18012 6662
rect 17960 6598 18012 6604
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17316 5772 17368 5778
rect 17316 5714 17368 5720
rect 17328 5574 17356 5714
rect 17316 5568 17368 5574
rect 17316 5510 17368 5516
rect 17328 5234 17356 5510
rect 17316 5228 17368 5234
rect 17316 5170 17368 5176
rect 16580 3596 16632 3602
rect 16580 3538 16632 3544
rect 16764 3596 16816 3602
rect 16764 3538 16816 3544
rect 16948 3596 17000 3602
rect 16948 3538 17000 3544
rect 16396 3188 16448 3194
rect 16396 3130 16448 3136
rect 16408 2990 16436 3130
rect 16396 2984 16448 2990
rect 16396 2926 16448 2932
rect 16212 2916 16264 2922
rect 16212 2858 16264 2864
rect 16776 2774 16804 3538
rect 16592 2746 16804 2774
rect 16212 2508 16264 2514
rect 16212 2450 16264 2456
rect 16224 800 16252 2450
rect 16396 2304 16448 2310
rect 16396 2246 16448 2252
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1122 0 1178 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7746 0 7802 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16408 134 16436 2246
rect 16592 800 16620 2746
rect 16960 800 16988 3538
rect 17682 3224 17738 3233
rect 17682 3159 17738 3168
rect 17696 3126 17724 3159
rect 17684 3120 17736 3126
rect 17684 3062 17736 3068
rect 17500 2984 17552 2990
rect 17498 2952 17500 2961
rect 17552 2952 17554 2961
rect 17498 2887 17554 2896
rect 17682 2816 17738 2825
rect 17682 2751 17738 2760
rect 17316 2508 17368 2514
rect 17316 2450 17368 2456
rect 17328 800 17356 2450
rect 17696 800 17724 2751
rect 17972 2446 18000 6598
rect 18064 6254 18092 6598
rect 18052 6248 18104 6254
rect 18052 6190 18104 6196
rect 18616 6118 18644 6734
rect 18512 6112 18564 6118
rect 18512 6054 18564 6060
rect 18604 6112 18656 6118
rect 18604 6054 18656 6060
rect 18524 5574 18552 6054
rect 18512 5568 18564 5574
rect 18512 5510 18564 5516
rect 18052 3596 18104 3602
rect 18052 3538 18104 3544
rect 17960 2440 18012 2446
rect 17960 2382 18012 2388
rect 17776 2304 17828 2310
rect 17776 2246 17828 2252
rect 16396 128 16448 134
rect 16396 70 16448 76
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 17788 202 17816 2246
rect 18064 800 18092 3538
rect 18512 2916 18564 2922
rect 18512 2858 18564 2864
rect 18524 2825 18552 2858
rect 18510 2816 18566 2825
rect 18510 2751 18566 2760
rect 18616 2650 18644 6054
rect 18708 5914 18736 6802
rect 19156 6248 19208 6254
rect 19156 6190 19208 6196
rect 18788 6180 18840 6186
rect 18788 6122 18840 6128
rect 18696 5908 18748 5914
rect 18696 5850 18748 5856
rect 18800 5794 18828 6122
rect 18708 5766 18828 5794
rect 18708 5302 18736 5766
rect 19168 5710 19196 6190
rect 20456 6118 20484 7210
rect 20720 7200 20772 7206
rect 20720 7142 20772 7148
rect 20534 6896 20590 6905
rect 20534 6831 20536 6840
rect 20588 6831 20590 6840
rect 20628 6860 20680 6866
rect 20536 6802 20588 6808
rect 20628 6802 20680 6808
rect 20536 6724 20588 6730
rect 20536 6666 20588 6672
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 20444 6112 20496 6118
rect 20444 6054 20496 6060
rect 19156 5704 19208 5710
rect 19156 5646 19208 5652
rect 18696 5296 18748 5302
rect 18696 5238 18748 5244
rect 18708 3398 18736 5238
rect 19168 5234 19196 5646
rect 19156 5228 19208 5234
rect 19156 5170 19208 5176
rect 19352 4214 19380 6054
rect 19580 6012 19876 6032
rect 19636 6010 19660 6012
rect 19716 6010 19740 6012
rect 19796 6010 19820 6012
rect 19658 5958 19660 6010
rect 19722 5958 19734 6010
rect 19796 5958 19798 6010
rect 19636 5956 19660 5958
rect 19716 5956 19740 5958
rect 19796 5956 19820 5958
rect 19580 5936 19876 5956
rect 20548 5302 20576 6666
rect 20640 6390 20668 6802
rect 20628 6384 20680 6390
rect 20628 6326 20680 6332
rect 20732 6254 20760 7142
rect 20720 6248 20772 6254
rect 20720 6190 20772 6196
rect 20720 5772 20772 5778
rect 20824 5760 20852 7686
rect 20904 7336 20956 7342
rect 20904 7278 20956 7284
rect 20916 6866 20944 7278
rect 20904 6860 20956 6866
rect 20904 6802 20956 6808
rect 21008 6769 21036 7822
rect 21088 6996 21140 7002
rect 21088 6938 21140 6944
rect 20994 6760 21050 6769
rect 20994 6695 21050 6704
rect 21008 6254 21036 6695
rect 20996 6248 21048 6254
rect 20996 6190 21048 6196
rect 20772 5732 20852 5760
rect 20720 5714 20772 5720
rect 20628 5704 20680 5710
rect 20626 5672 20628 5681
rect 20680 5672 20682 5681
rect 20626 5607 20682 5616
rect 20536 5296 20588 5302
rect 20536 5238 20588 5244
rect 20548 5030 20576 5238
rect 21100 5166 21128 6938
rect 21192 6662 21220 7890
rect 21180 6656 21232 6662
rect 21180 6598 21232 6604
rect 21192 6322 21220 6598
rect 21284 6458 21312 7958
rect 23480 7744 23532 7750
rect 23480 7686 23532 7692
rect 22190 7576 22246 7585
rect 22190 7511 22192 7520
rect 22244 7511 22246 7520
rect 22192 7482 22244 7488
rect 23020 7336 23072 7342
rect 23020 7278 23072 7284
rect 22008 7268 22060 7274
rect 22008 7210 22060 7216
rect 21732 6928 21784 6934
rect 21732 6870 21784 6876
rect 21548 6860 21600 6866
rect 21548 6802 21600 6808
rect 21560 6769 21588 6802
rect 21546 6760 21602 6769
rect 21744 6730 21772 6870
rect 21546 6695 21602 6704
rect 21732 6724 21784 6730
rect 21732 6666 21784 6672
rect 21272 6452 21324 6458
rect 21272 6394 21324 6400
rect 21180 6316 21232 6322
rect 21180 6258 21232 6264
rect 21548 6112 21600 6118
rect 21548 6054 21600 6060
rect 21824 6112 21876 6118
rect 21824 6054 21876 6060
rect 21088 5160 21140 5166
rect 21088 5102 21140 5108
rect 21560 5098 21588 6054
rect 21640 5704 21692 5710
rect 21638 5672 21640 5681
rect 21692 5672 21694 5681
rect 21638 5607 21694 5616
rect 21640 5568 21692 5574
rect 21640 5510 21692 5516
rect 21548 5092 21600 5098
rect 21548 5034 21600 5040
rect 20536 5024 20588 5030
rect 20536 4966 20588 4972
rect 19580 4924 19876 4944
rect 19636 4922 19660 4924
rect 19716 4922 19740 4924
rect 19796 4922 19820 4924
rect 19658 4870 19660 4922
rect 19722 4870 19734 4922
rect 19796 4870 19798 4922
rect 19636 4868 19660 4870
rect 19716 4868 19740 4870
rect 19796 4868 19820 4870
rect 19580 4848 19876 4868
rect 20076 4820 20128 4826
rect 20076 4762 20128 4768
rect 19340 4208 19392 4214
rect 19340 4150 19392 4156
rect 20088 4078 20116 4762
rect 21548 4684 21600 4690
rect 21548 4626 21600 4632
rect 20076 4072 20128 4078
rect 20076 4014 20128 4020
rect 20260 4072 20312 4078
rect 20260 4014 20312 4020
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 18880 3936 18932 3942
rect 18880 3878 18932 3884
rect 18800 3482 18828 3878
rect 18892 3670 18920 3878
rect 19580 3836 19876 3856
rect 19636 3834 19660 3836
rect 19716 3834 19740 3836
rect 19796 3834 19820 3836
rect 19658 3782 19660 3834
rect 19722 3782 19734 3834
rect 19796 3782 19798 3834
rect 19636 3780 19660 3782
rect 19716 3780 19740 3782
rect 19796 3780 19820 3782
rect 19580 3760 19876 3780
rect 18880 3664 18932 3670
rect 18880 3606 18932 3612
rect 19156 3596 19208 3602
rect 19156 3538 19208 3544
rect 18800 3454 18920 3482
rect 18696 3392 18748 3398
rect 18696 3334 18748 3340
rect 18788 3392 18840 3398
rect 18788 3334 18840 3340
rect 18604 2644 18656 2650
rect 18604 2586 18656 2592
rect 18420 2440 18472 2446
rect 18420 2382 18472 2388
rect 18432 800 18460 2382
rect 18800 800 18828 3334
rect 18892 2938 18920 3454
rect 19064 3392 19116 3398
rect 19064 3334 19116 3340
rect 19076 3233 19104 3334
rect 19062 3224 19118 3233
rect 19062 3159 19118 3168
rect 18892 2922 19012 2938
rect 18892 2916 19024 2922
rect 18892 2910 18972 2916
rect 18972 2858 19024 2864
rect 19168 800 19196 3538
rect 19892 2984 19944 2990
rect 19892 2926 19944 2932
rect 19580 2748 19876 2768
rect 19636 2746 19660 2748
rect 19716 2746 19740 2748
rect 19796 2746 19820 2748
rect 19658 2694 19660 2746
rect 19722 2694 19734 2746
rect 19796 2694 19798 2746
rect 19636 2692 19660 2694
rect 19716 2692 19740 2694
rect 19796 2692 19820 2694
rect 19580 2672 19876 2692
rect 19524 2440 19576 2446
rect 19524 2382 19576 2388
rect 19536 800 19564 2382
rect 19904 800 19932 2926
rect 20272 800 20300 4014
rect 20902 3632 20958 3641
rect 20902 3567 20958 3576
rect 21272 3596 21324 3602
rect 20916 3398 20944 3567
rect 21272 3538 21324 3544
rect 21364 3596 21416 3602
rect 21364 3538 21416 3544
rect 21284 3505 21312 3538
rect 21270 3496 21326 3505
rect 21270 3431 21326 3440
rect 20904 3392 20956 3398
rect 20904 3334 20956 3340
rect 20996 3392 21048 3398
rect 20996 3334 21048 3340
rect 20628 2984 20680 2990
rect 20628 2926 20680 2932
rect 20904 2984 20956 2990
rect 20904 2926 20956 2932
rect 20536 2440 20588 2446
rect 20536 2382 20588 2388
rect 20548 1698 20576 2382
rect 20536 1692 20588 1698
rect 20536 1634 20588 1640
rect 20640 800 20668 2926
rect 17776 196 17828 202
rect 17776 138 17828 144
rect 18050 0 18106 800
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20258 0 20314 800
rect 20626 0 20682 800
rect 20916 406 20944 2926
rect 21008 800 21036 3334
rect 21086 3224 21142 3233
rect 21086 3159 21142 3168
rect 21272 3188 21324 3194
rect 21100 3126 21128 3159
rect 21272 3130 21324 3136
rect 21088 3120 21140 3126
rect 21088 3062 21140 3068
rect 21284 2854 21312 3130
rect 21272 2848 21324 2854
rect 21272 2790 21324 2796
rect 21376 800 21404 3538
rect 21560 3534 21588 4626
rect 21652 4049 21680 5510
rect 21836 4146 21864 6054
rect 22020 5574 22048 7210
rect 22284 7200 22336 7206
rect 22284 7142 22336 7148
rect 22100 6724 22152 6730
rect 22100 6666 22152 6672
rect 22112 5846 22140 6666
rect 22100 5840 22152 5846
rect 22100 5782 22152 5788
rect 22296 5778 22324 7142
rect 23032 6905 23060 7278
rect 23204 7268 23256 7274
rect 23204 7210 23256 7216
rect 23216 7002 23244 7210
rect 23204 6996 23256 7002
rect 23204 6938 23256 6944
rect 23018 6896 23074 6905
rect 23018 6831 23074 6840
rect 23032 6730 23060 6831
rect 23020 6724 23072 6730
rect 23020 6666 23072 6672
rect 23492 5846 23520 7686
rect 23848 6248 23900 6254
rect 23848 6190 23900 6196
rect 23480 5840 23532 5846
rect 23480 5782 23532 5788
rect 23860 5778 23888 6190
rect 22284 5772 22336 5778
rect 22284 5714 22336 5720
rect 23848 5772 23900 5778
rect 23848 5714 23900 5720
rect 24228 5574 24256 7958
rect 25596 7948 25648 7954
rect 25596 7890 25648 7896
rect 25964 7948 26016 7954
rect 25964 7890 26016 7896
rect 26424 7948 26476 7954
rect 26424 7890 26476 7896
rect 27620 7948 27672 7954
rect 27620 7890 27672 7896
rect 27896 7948 27948 7954
rect 28170 7919 28226 7928
rect 28264 7948 28316 7954
rect 27896 7890 27948 7896
rect 28264 7890 28316 7896
rect 25608 7342 25636 7890
rect 25976 7410 26004 7890
rect 26240 7812 26292 7818
rect 26240 7754 26292 7760
rect 25964 7404 26016 7410
rect 25964 7346 26016 7352
rect 25596 7336 25648 7342
rect 25596 7278 25648 7284
rect 26252 7274 26280 7754
rect 26332 7744 26384 7750
rect 26332 7686 26384 7692
rect 26240 7268 26292 7274
rect 26240 7210 26292 7216
rect 24952 7200 25004 7206
rect 24952 7142 25004 7148
rect 25044 7200 25096 7206
rect 25044 7142 25096 7148
rect 24964 6934 24992 7142
rect 24952 6928 25004 6934
rect 24952 6870 25004 6876
rect 25056 6254 25084 7142
rect 25044 6248 25096 6254
rect 25044 6190 25096 6196
rect 26344 5846 26372 7686
rect 26436 7342 26464 7890
rect 26514 7440 26570 7449
rect 26514 7375 26570 7384
rect 27436 7404 27488 7410
rect 26528 7342 26556 7375
rect 27436 7346 27488 7352
rect 26424 7336 26476 7342
rect 26424 7278 26476 7284
rect 26516 7336 26568 7342
rect 26516 7278 26568 7284
rect 26608 7268 26660 7274
rect 26608 7210 26660 7216
rect 26620 6118 26648 7210
rect 26608 6112 26660 6118
rect 26608 6054 26660 6060
rect 27448 5846 27476 7346
rect 27632 7342 27660 7890
rect 27620 7336 27672 7342
rect 27620 7278 27672 7284
rect 27804 6248 27856 6254
rect 27804 6190 27856 6196
rect 26332 5840 26384 5846
rect 26332 5782 26384 5788
rect 27436 5840 27488 5846
rect 27436 5782 27488 5788
rect 27816 5778 27844 6190
rect 27804 5772 27856 5778
rect 27804 5714 27856 5720
rect 22008 5568 22060 5574
rect 24216 5568 24268 5574
rect 22008 5510 22060 5516
rect 24136 5528 24216 5556
rect 23756 5364 23808 5370
rect 23756 5306 23808 5312
rect 23768 4758 23796 5306
rect 23756 4752 23808 4758
rect 23756 4694 23808 4700
rect 21916 4548 21968 4554
rect 21916 4490 21968 4496
rect 21928 4214 21956 4490
rect 21916 4208 21968 4214
rect 21916 4150 21968 4156
rect 21824 4140 21876 4146
rect 21824 4082 21876 4088
rect 22020 4100 22232 4128
rect 21638 4040 21694 4049
rect 21638 3975 21694 3984
rect 21548 3528 21600 3534
rect 21548 3470 21600 3476
rect 22020 3466 22048 4100
rect 22098 4040 22154 4049
rect 22098 3975 22154 3984
rect 22112 3942 22140 3975
rect 22204 3942 22232 4100
rect 22376 4072 22428 4078
rect 22376 4014 22428 4020
rect 22100 3936 22152 3942
rect 22100 3878 22152 3884
rect 22192 3936 22244 3942
rect 22192 3878 22244 3884
rect 22388 3754 22416 4014
rect 22112 3726 22416 3754
rect 22008 3460 22060 3466
rect 22008 3402 22060 3408
rect 22112 2938 22140 3726
rect 22468 3596 22520 3602
rect 22468 3538 22520 3544
rect 23572 3596 23624 3602
rect 23572 3538 23624 3544
rect 22284 3528 22336 3534
rect 22282 3496 22284 3505
rect 22336 3496 22338 3505
rect 22282 3431 22338 3440
rect 22376 3120 22428 3126
rect 22374 3088 22376 3097
rect 22428 3088 22430 3097
rect 22374 3023 22430 3032
rect 22020 2922 22140 2938
rect 22008 2916 22140 2922
rect 22060 2910 22140 2916
rect 22008 2858 22060 2864
rect 22100 2848 22152 2854
rect 22100 2790 22152 2796
rect 21732 2508 21784 2514
rect 21732 2450 21784 2456
rect 21744 800 21772 2450
rect 21916 2304 21968 2310
rect 21916 2246 21968 2252
rect 20904 400 20956 406
rect 20904 342 20956 348
rect 20994 0 21050 800
rect 21362 0 21418 800
rect 21730 0 21786 800
rect 21928 338 21956 2246
rect 22112 800 22140 2790
rect 22480 800 22508 3538
rect 22652 3392 22704 3398
rect 22652 3334 22704 3340
rect 22664 2990 22692 3334
rect 22652 2984 22704 2990
rect 22652 2926 22704 2932
rect 23204 2848 23256 2854
rect 23204 2790 23256 2796
rect 22836 2508 22888 2514
rect 22836 2450 22888 2456
rect 22848 800 22876 2450
rect 23112 2304 23164 2310
rect 23112 2246 23164 2252
rect 21916 332 21968 338
rect 21916 274 21968 280
rect 22098 0 22154 800
rect 22466 0 22522 800
rect 22834 0 22890 800
rect 23124 474 23152 2246
rect 23216 800 23244 2790
rect 23584 800 23612 3538
rect 24136 3534 24164 5528
rect 24216 5510 24268 5516
rect 26608 5568 26660 5574
rect 26608 5510 26660 5516
rect 27804 5568 27856 5574
rect 27908 5556 27936 7890
rect 28276 7818 28304 7890
rect 28264 7812 28316 7818
rect 28264 7754 28316 7760
rect 28538 7712 28594 7721
rect 28538 7647 28594 7656
rect 28552 7342 28580 7647
rect 28448 7336 28500 7342
rect 28446 7304 28448 7313
rect 28540 7336 28592 7342
rect 28500 7304 28502 7313
rect 28540 7278 28592 7284
rect 28446 7239 28502 7248
rect 28644 7177 28672 9646
rect 29092 9512 29144 9518
rect 29092 9454 29144 9460
rect 28816 7880 28868 7886
rect 28816 7822 28868 7828
rect 28828 7324 28856 7822
rect 28906 7576 28962 7585
rect 29104 7562 29132 9454
rect 29932 8022 29960 13926
rect 30840 13874 30892 13880
rect 30852 13394 30880 13874
rect 30840 13388 30892 13394
rect 30840 13330 30892 13336
rect 30852 12850 30880 13330
rect 30840 12844 30892 12850
rect 30840 12786 30892 12792
rect 30196 9444 30248 9450
rect 30196 9386 30248 9392
rect 29920 8016 29972 8022
rect 29920 7958 29972 7964
rect 29368 7948 29420 7954
rect 29368 7890 29420 7896
rect 29184 7880 29236 7886
rect 29184 7822 29236 7828
rect 28962 7534 29132 7562
rect 28906 7511 28962 7520
rect 28908 7336 28960 7342
rect 28828 7296 28908 7324
rect 28908 7278 28960 7284
rect 29196 7274 29224 7822
rect 29276 7744 29328 7750
rect 29276 7686 29328 7692
rect 28724 7268 28776 7274
rect 28724 7210 28776 7216
rect 29184 7268 29236 7274
rect 29184 7210 29236 7216
rect 28630 7168 28686 7177
rect 28630 7103 28686 7112
rect 28538 6760 28594 6769
rect 28538 6695 28594 6704
rect 28552 6662 28580 6695
rect 28540 6656 28592 6662
rect 28540 6598 28592 6604
rect 28552 6118 28580 6598
rect 28540 6112 28592 6118
rect 28540 6054 28592 6060
rect 28736 5642 28764 7210
rect 29092 7200 29144 7206
rect 28906 7168 28962 7177
rect 28906 7103 28962 7112
rect 29012 7160 29092 7188
rect 28920 6866 28948 7103
rect 28908 6860 28960 6866
rect 28908 6802 28960 6808
rect 28908 6248 28960 6254
rect 28828 6196 28908 6202
rect 28828 6190 28960 6196
rect 28828 6174 28948 6190
rect 29012 6186 29040 7160
rect 29092 7142 29144 7148
rect 29196 6934 29224 7210
rect 29288 7206 29316 7686
rect 29380 7206 29408 7890
rect 29644 7540 29696 7546
rect 29644 7482 29696 7488
rect 29656 7313 29684 7482
rect 29932 7342 29960 7958
rect 29920 7336 29972 7342
rect 29642 7304 29698 7313
rect 29920 7278 29972 7284
rect 29642 7239 29698 7248
rect 29276 7200 29328 7206
rect 29276 7142 29328 7148
rect 29368 7200 29420 7206
rect 29368 7142 29420 7148
rect 29184 6928 29236 6934
rect 29184 6870 29236 6876
rect 29196 6662 29224 6870
rect 29380 6866 29408 7142
rect 29368 6860 29420 6866
rect 29368 6802 29420 6808
rect 29184 6656 29236 6662
rect 29184 6598 29236 6604
rect 30208 6458 30236 9386
rect 30932 8968 30984 8974
rect 30932 8910 30984 8916
rect 30380 8016 30432 8022
rect 30380 7958 30432 7964
rect 30288 6792 30340 6798
rect 30286 6760 30288 6769
rect 30340 6760 30342 6769
rect 30286 6695 30342 6704
rect 30196 6452 30248 6458
rect 30196 6394 30248 6400
rect 30392 6390 30420 7958
rect 30472 7948 30524 7954
rect 30472 7890 30524 7896
rect 30484 7546 30512 7890
rect 30472 7540 30524 7546
rect 30472 7482 30524 7488
rect 30748 7472 30800 7478
rect 30748 7414 30800 7420
rect 30656 7336 30708 7342
rect 30470 7304 30526 7313
rect 30656 7278 30708 7284
rect 30470 7239 30526 7248
rect 30380 6384 30432 6390
rect 30380 6326 30432 6332
rect 29000 6180 29052 6186
rect 28724 5636 28776 5642
rect 28724 5578 28776 5584
rect 27856 5528 27936 5556
rect 27988 5568 28040 5574
rect 27804 5510 27856 5516
rect 27988 5510 28040 5516
rect 24952 5160 25004 5166
rect 24952 5102 25004 5108
rect 25412 5160 25464 5166
rect 25412 5102 25464 5108
rect 24964 4146 24992 5102
rect 24952 4140 25004 4146
rect 24952 4082 25004 4088
rect 24676 3596 24728 3602
rect 24676 3538 24728 3544
rect 24124 3528 24176 3534
rect 24124 3470 24176 3476
rect 24320 3318 24624 3346
rect 24320 3194 24348 3318
rect 24596 3194 24624 3318
rect 24308 3188 24360 3194
rect 24308 3130 24360 3136
rect 24492 3188 24544 3194
rect 24492 3130 24544 3136
rect 24584 3188 24636 3194
rect 24584 3130 24636 3136
rect 24504 3074 24532 3130
rect 24228 3046 24532 3074
rect 24228 2774 24256 3046
rect 24308 2984 24360 2990
rect 24584 2984 24636 2990
rect 24360 2932 24584 2938
rect 24308 2926 24636 2932
rect 24320 2910 24624 2926
rect 24228 2746 24348 2774
rect 23940 2508 23992 2514
rect 23940 2450 23992 2456
rect 23952 800 23980 2450
rect 24124 2304 24176 2310
rect 24124 2246 24176 2252
rect 24136 882 24164 2246
rect 24124 876 24176 882
rect 24124 818 24176 824
rect 24320 800 24348 2746
rect 24688 800 24716 3538
rect 25320 3528 25372 3534
rect 25320 3470 25372 3476
rect 25332 2922 25360 3470
rect 25424 3058 25452 5102
rect 26620 4826 26648 5510
rect 28000 5216 28028 5510
rect 28828 5370 28856 6174
rect 29000 6122 29052 6128
rect 29276 5772 29328 5778
rect 29276 5714 29328 5720
rect 28816 5364 28868 5370
rect 28816 5306 28868 5312
rect 29288 5234 29316 5714
rect 27908 5188 28028 5216
rect 28172 5228 28224 5234
rect 26608 4820 26660 4826
rect 26608 4762 26660 4768
rect 27908 4690 27936 5188
rect 28172 5170 28224 5176
rect 29276 5228 29328 5234
rect 29276 5170 29328 5176
rect 27988 5092 28040 5098
rect 27988 5034 28040 5040
rect 28000 4758 28028 5034
rect 27988 4752 28040 4758
rect 27988 4694 28040 4700
rect 27896 4684 27948 4690
rect 27896 4626 27948 4632
rect 28080 4684 28132 4690
rect 28080 4626 28132 4632
rect 25504 4140 25556 4146
rect 25504 4082 25556 4088
rect 25412 3052 25464 3058
rect 25412 2994 25464 3000
rect 25516 2922 25544 4082
rect 27896 3936 27948 3942
rect 27896 3878 27948 3884
rect 25780 3596 25832 3602
rect 25780 3538 25832 3544
rect 26884 3596 26936 3602
rect 26884 3538 26936 3544
rect 25320 2916 25372 2922
rect 25320 2858 25372 2864
rect 25504 2916 25556 2922
rect 25504 2858 25556 2864
rect 25412 2848 25464 2854
rect 25412 2790 25464 2796
rect 25044 2508 25096 2514
rect 25044 2450 25096 2456
rect 25056 800 25084 2450
rect 25424 800 25452 2790
rect 25792 800 25820 3538
rect 26516 2848 26568 2854
rect 26516 2790 26568 2796
rect 26148 2508 26200 2514
rect 26148 2450 26200 2456
rect 25964 2304 26016 2310
rect 25964 2246 26016 2252
rect 23112 468 23164 474
rect 23112 410 23164 416
rect 23202 0 23258 800
rect 23570 0 23626 800
rect 23938 0 23994 800
rect 24306 0 24362 800
rect 24674 0 24730 800
rect 25042 0 25098 800
rect 25410 0 25466 800
rect 25778 0 25834 800
rect 25976 270 26004 2246
rect 26160 800 26188 2450
rect 26528 800 26556 2790
rect 26608 2372 26660 2378
rect 26608 2314 26660 2320
rect 25964 264 26016 270
rect 25964 206 26016 212
rect 26146 0 26202 800
rect 26514 0 26570 800
rect 26620 746 26648 2314
rect 26896 800 26924 3538
rect 27908 2922 27936 3878
rect 27988 3596 28040 3602
rect 27988 3538 28040 3544
rect 27896 2916 27948 2922
rect 27896 2858 27948 2864
rect 27620 2848 27672 2854
rect 27620 2790 27672 2796
rect 27252 2508 27304 2514
rect 27252 2450 27304 2456
rect 27264 800 27292 2450
rect 27344 2372 27396 2378
rect 27344 2314 27396 2320
rect 27356 950 27384 2314
rect 27344 944 27396 950
rect 27344 886 27396 892
rect 27632 800 27660 2790
rect 28000 800 28028 3538
rect 28092 3126 28120 4626
rect 28184 4622 28212 5170
rect 28356 5024 28408 5030
rect 28356 4966 28408 4972
rect 28368 4826 28396 4966
rect 28356 4820 28408 4826
rect 28356 4762 28408 4768
rect 28908 4684 28960 4690
rect 28908 4626 28960 4632
rect 28172 4616 28224 4622
rect 28172 4558 28224 4564
rect 28816 3664 28868 3670
rect 28920 3641 28948 4626
rect 28816 3606 28868 3612
rect 28906 3632 28962 3641
rect 28172 3596 28224 3602
rect 28172 3538 28224 3544
rect 28184 3233 28212 3538
rect 28170 3224 28226 3233
rect 28170 3159 28226 3168
rect 28080 3120 28132 3126
rect 28172 3120 28224 3126
rect 28080 3062 28132 3068
rect 28170 3088 28172 3097
rect 28224 3088 28226 3097
rect 28170 3023 28226 3032
rect 28828 2922 28856 3606
rect 30392 3602 30420 6326
rect 30484 5030 30512 7239
rect 30564 7200 30616 7206
rect 30564 7142 30616 7148
rect 30576 6866 30604 7142
rect 30564 6860 30616 6866
rect 30564 6802 30616 6808
rect 30576 6186 30604 6802
rect 30564 6180 30616 6186
rect 30564 6122 30616 6128
rect 30668 5574 30696 7278
rect 30656 5568 30708 5574
rect 30656 5510 30708 5516
rect 30564 5364 30616 5370
rect 30564 5306 30616 5312
rect 30576 5030 30604 5306
rect 30760 5148 30788 7414
rect 30840 6656 30892 6662
rect 30840 6598 30892 6604
rect 30668 5120 30788 5148
rect 30472 5024 30524 5030
rect 30472 4966 30524 4972
rect 30564 5024 30616 5030
rect 30564 4966 30616 4972
rect 30484 4622 30512 4966
rect 30472 4616 30524 4622
rect 30472 4558 30524 4564
rect 30576 4049 30604 4966
rect 30562 4040 30618 4049
rect 30562 3975 30618 3984
rect 28906 3567 28962 3576
rect 30380 3596 30432 3602
rect 30380 3538 30432 3544
rect 30668 3126 30696 5120
rect 30748 5024 30800 5030
rect 30748 4966 30800 4972
rect 30760 4554 30788 4966
rect 30748 4548 30800 4554
rect 30748 4490 30800 4496
rect 30656 3120 30708 3126
rect 30656 3062 30708 3068
rect 29092 2984 29144 2990
rect 29092 2926 29144 2932
rect 30196 2984 30248 2990
rect 30196 2926 30248 2932
rect 28816 2916 28868 2922
rect 28816 2858 28868 2864
rect 28724 2848 28776 2854
rect 28724 2790 28776 2796
rect 28356 2508 28408 2514
rect 28356 2450 28408 2456
rect 28368 800 28396 2450
rect 28632 2372 28684 2378
rect 28632 2314 28684 2320
rect 28644 814 28672 2314
rect 28632 808 28684 814
rect 26608 740 26660 746
rect 26608 682 26660 688
rect 26882 0 26938 800
rect 27250 0 27306 800
rect 27618 0 27674 800
rect 27986 0 28042 800
rect 28354 0 28410 800
rect 28736 800 28764 2790
rect 29104 800 29132 2926
rect 29460 2508 29512 2514
rect 29460 2450 29512 2456
rect 29472 800 29500 2450
rect 29736 2372 29788 2378
rect 29736 2314 29788 2320
rect 29828 2372 29880 2378
rect 29828 2314 29880 2320
rect 28632 750 28684 756
rect 28722 0 28778 800
rect 29090 0 29146 800
rect 29458 0 29514 800
rect 29748 678 29776 2314
rect 29840 800 29868 2314
rect 30208 800 30236 2926
rect 30564 2508 30616 2514
rect 30564 2450 30616 2456
rect 30576 800 30604 2450
rect 30852 2310 30880 6598
rect 30944 5370 30972 8910
rect 31024 7948 31076 7954
rect 31024 7890 31076 7896
rect 31036 6934 31064 7890
rect 31128 7274 31156 14418
rect 31220 14414 31248 14962
rect 31208 14408 31260 14414
rect 31208 14350 31260 14356
rect 31392 8900 31444 8906
rect 31392 8842 31444 8848
rect 31404 7954 31432 8842
rect 31392 7948 31444 7954
rect 31392 7890 31444 7896
rect 31300 7336 31352 7342
rect 31298 7304 31300 7313
rect 31352 7304 31354 7313
rect 31116 7268 31168 7274
rect 31298 7239 31354 7248
rect 31116 7210 31168 7216
rect 31496 7154 31524 15302
rect 31772 14550 31800 116078
rect 32140 22574 32168 117098
rect 33416 117088 33468 117094
rect 33416 117030 33468 117036
rect 33140 24064 33192 24070
rect 33140 24006 33192 24012
rect 33152 22642 33180 24006
rect 33140 22636 33192 22642
rect 33140 22578 33192 22584
rect 32128 22568 32180 22574
rect 32128 22510 32180 22516
rect 32140 22094 32168 22510
rect 33428 22438 33456 117030
rect 34940 116444 35236 116464
rect 34996 116442 35020 116444
rect 35076 116442 35100 116444
rect 35156 116442 35180 116444
rect 35018 116390 35020 116442
rect 35082 116390 35094 116442
rect 35156 116390 35158 116442
rect 34996 116388 35020 116390
rect 35076 116388 35100 116390
rect 35156 116388 35180 116390
rect 34940 116368 35236 116388
rect 35268 116346 35296 117166
rect 36820 117156 36872 117162
rect 36820 117098 36872 117104
rect 39764 117156 39816 117162
rect 39764 117098 39816 117104
rect 41696 117156 41748 117162
rect 41696 117098 41748 117104
rect 44364 117156 44416 117162
rect 44364 117098 44416 117104
rect 47032 117156 47084 117162
rect 47032 117098 47084 117104
rect 48964 117156 49016 117162
rect 48964 117098 49016 117104
rect 50896 117156 50948 117162
rect 50896 117098 50948 117104
rect 54024 117156 54076 117162
rect 54024 117098 54076 117104
rect 55588 117156 55640 117162
rect 55588 117098 55640 117104
rect 58256 117156 58308 117162
rect 58256 117098 58308 117104
rect 60372 117156 60424 117162
rect 60372 117098 60424 117104
rect 62948 117156 63000 117162
rect 62948 117098 63000 117104
rect 65524 117156 65576 117162
rect 65524 117098 65576 117104
rect 67640 117156 67692 117162
rect 67640 117098 67692 117104
rect 69664 117156 69716 117162
rect 69664 117098 69716 117104
rect 72424 117156 72476 117162
rect 72424 117098 72476 117104
rect 35256 116340 35308 116346
rect 35256 116282 35308 116288
rect 34940 115356 35236 115376
rect 34996 115354 35020 115356
rect 35076 115354 35100 115356
rect 35156 115354 35180 115356
rect 35018 115302 35020 115354
rect 35082 115302 35094 115354
rect 35156 115302 35158 115354
rect 34996 115300 35020 115302
rect 35076 115300 35100 115302
rect 35156 115300 35180 115302
rect 34940 115280 35236 115300
rect 34940 114268 35236 114288
rect 34996 114266 35020 114268
rect 35076 114266 35100 114268
rect 35156 114266 35180 114268
rect 35018 114214 35020 114266
rect 35082 114214 35094 114266
rect 35156 114214 35158 114266
rect 34996 114212 35020 114214
rect 35076 114212 35100 114214
rect 35156 114212 35180 114214
rect 34940 114192 35236 114212
rect 34940 113180 35236 113200
rect 34996 113178 35020 113180
rect 35076 113178 35100 113180
rect 35156 113178 35180 113180
rect 35018 113126 35020 113178
rect 35082 113126 35094 113178
rect 35156 113126 35158 113178
rect 34996 113124 35020 113126
rect 35076 113124 35100 113126
rect 35156 113124 35180 113126
rect 34940 113104 35236 113124
rect 34940 112092 35236 112112
rect 34996 112090 35020 112092
rect 35076 112090 35100 112092
rect 35156 112090 35180 112092
rect 35018 112038 35020 112090
rect 35082 112038 35094 112090
rect 35156 112038 35158 112090
rect 34996 112036 35020 112038
rect 35076 112036 35100 112038
rect 35156 112036 35180 112038
rect 34940 112016 35236 112036
rect 34940 111004 35236 111024
rect 34996 111002 35020 111004
rect 35076 111002 35100 111004
rect 35156 111002 35180 111004
rect 35018 110950 35020 111002
rect 35082 110950 35094 111002
rect 35156 110950 35158 111002
rect 34996 110948 35020 110950
rect 35076 110948 35100 110950
rect 35156 110948 35180 110950
rect 34940 110928 35236 110948
rect 34940 109916 35236 109936
rect 34996 109914 35020 109916
rect 35076 109914 35100 109916
rect 35156 109914 35180 109916
rect 35018 109862 35020 109914
rect 35082 109862 35094 109914
rect 35156 109862 35158 109914
rect 34996 109860 35020 109862
rect 35076 109860 35100 109862
rect 35156 109860 35180 109862
rect 34940 109840 35236 109860
rect 34940 108828 35236 108848
rect 34996 108826 35020 108828
rect 35076 108826 35100 108828
rect 35156 108826 35180 108828
rect 35018 108774 35020 108826
rect 35082 108774 35094 108826
rect 35156 108774 35158 108826
rect 34996 108772 35020 108774
rect 35076 108772 35100 108774
rect 35156 108772 35180 108774
rect 34940 108752 35236 108772
rect 34940 107740 35236 107760
rect 34996 107738 35020 107740
rect 35076 107738 35100 107740
rect 35156 107738 35180 107740
rect 35018 107686 35020 107738
rect 35082 107686 35094 107738
rect 35156 107686 35158 107738
rect 34996 107684 35020 107686
rect 35076 107684 35100 107686
rect 35156 107684 35180 107686
rect 34940 107664 35236 107684
rect 34940 106652 35236 106672
rect 34996 106650 35020 106652
rect 35076 106650 35100 106652
rect 35156 106650 35180 106652
rect 35018 106598 35020 106650
rect 35082 106598 35094 106650
rect 35156 106598 35158 106650
rect 34996 106596 35020 106598
rect 35076 106596 35100 106598
rect 35156 106596 35180 106598
rect 34940 106576 35236 106596
rect 34940 105564 35236 105584
rect 34996 105562 35020 105564
rect 35076 105562 35100 105564
rect 35156 105562 35180 105564
rect 35018 105510 35020 105562
rect 35082 105510 35094 105562
rect 35156 105510 35158 105562
rect 34996 105508 35020 105510
rect 35076 105508 35100 105510
rect 35156 105508 35180 105510
rect 34940 105488 35236 105508
rect 34940 104476 35236 104496
rect 34996 104474 35020 104476
rect 35076 104474 35100 104476
rect 35156 104474 35180 104476
rect 35018 104422 35020 104474
rect 35082 104422 35094 104474
rect 35156 104422 35158 104474
rect 34996 104420 35020 104422
rect 35076 104420 35100 104422
rect 35156 104420 35180 104422
rect 34940 104400 35236 104420
rect 34940 103388 35236 103408
rect 34996 103386 35020 103388
rect 35076 103386 35100 103388
rect 35156 103386 35180 103388
rect 35018 103334 35020 103386
rect 35082 103334 35094 103386
rect 35156 103334 35158 103386
rect 34996 103332 35020 103334
rect 35076 103332 35100 103334
rect 35156 103332 35180 103334
rect 34940 103312 35236 103332
rect 34940 102300 35236 102320
rect 34996 102298 35020 102300
rect 35076 102298 35100 102300
rect 35156 102298 35180 102300
rect 35018 102246 35020 102298
rect 35082 102246 35094 102298
rect 35156 102246 35158 102298
rect 34996 102244 35020 102246
rect 35076 102244 35100 102246
rect 35156 102244 35180 102246
rect 34940 102224 35236 102244
rect 34940 101212 35236 101232
rect 34996 101210 35020 101212
rect 35076 101210 35100 101212
rect 35156 101210 35180 101212
rect 35018 101158 35020 101210
rect 35082 101158 35094 101210
rect 35156 101158 35158 101210
rect 34996 101156 35020 101158
rect 35076 101156 35100 101158
rect 35156 101156 35180 101158
rect 34940 101136 35236 101156
rect 34940 100124 35236 100144
rect 34996 100122 35020 100124
rect 35076 100122 35100 100124
rect 35156 100122 35180 100124
rect 35018 100070 35020 100122
rect 35082 100070 35094 100122
rect 35156 100070 35158 100122
rect 34996 100068 35020 100070
rect 35076 100068 35100 100070
rect 35156 100068 35180 100070
rect 34940 100048 35236 100068
rect 34940 99036 35236 99056
rect 34996 99034 35020 99036
rect 35076 99034 35100 99036
rect 35156 99034 35180 99036
rect 35018 98982 35020 99034
rect 35082 98982 35094 99034
rect 35156 98982 35158 99034
rect 34996 98980 35020 98982
rect 35076 98980 35100 98982
rect 35156 98980 35180 98982
rect 34940 98960 35236 98980
rect 34940 97948 35236 97968
rect 34996 97946 35020 97948
rect 35076 97946 35100 97948
rect 35156 97946 35180 97948
rect 35018 97894 35020 97946
rect 35082 97894 35094 97946
rect 35156 97894 35158 97946
rect 34996 97892 35020 97894
rect 35076 97892 35100 97894
rect 35156 97892 35180 97894
rect 34940 97872 35236 97892
rect 34940 96860 35236 96880
rect 34996 96858 35020 96860
rect 35076 96858 35100 96860
rect 35156 96858 35180 96860
rect 35018 96806 35020 96858
rect 35082 96806 35094 96858
rect 35156 96806 35158 96858
rect 34996 96804 35020 96806
rect 35076 96804 35100 96806
rect 35156 96804 35180 96806
rect 34940 96784 35236 96804
rect 34940 95772 35236 95792
rect 34996 95770 35020 95772
rect 35076 95770 35100 95772
rect 35156 95770 35180 95772
rect 35018 95718 35020 95770
rect 35082 95718 35094 95770
rect 35156 95718 35158 95770
rect 34996 95716 35020 95718
rect 35076 95716 35100 95718
rect 35156 95716 35180 95718
rect 34940 95696 35236 95716
rect 34940 94684 35236 94704
rect 34996 94682 35020 94684
rect 35076 94682 35100 94684
rect 35156 94682 35180 94684
rect 35018 94630 35020 94682
rect 35082 94630 35094 94682
rect 35156 94630 35158 94682
rect 34996 94628 35020 94630
rect 35076 94628 35100 94630
rect 35156 94628 35180 94630
rect 34940 94608 35236 94628
rect 34940 93596 35236 93616
rect 34996 93594 35020 93596
rect 35076 93594 35100 93596
rect 35156 93594 35180 93596
rect 35018 93542 35020 93594
rect 35082 93542 35094 93594
rect 35156 93542 35158 93594
rect 34996 93540 35020 93542
rect 35076 93540 35100 93542
rect 35156 93540 35180 93542
rect 34940 93520 35236 93540
rect 34940 92508 35236 92528
rect 34996 92506 35020 92508
rect 35076 92506 35100 92508
rect 35156 92506 35180 92508
rect 35018 92454 35020 92506
rect 35082 92454 35094 92506
rect 35156 92454 35158 92506
rect 34996 92452 35020 92454
rect 35076 92452 35100 92454
rect 35156 92452 35180 92454
rect 34940 92432 35236 92452
rect 34940 91420 35236 91440
rect 34996 91418 35020 91420
rect 35076 91418 35100 91420
rect 35156 91418 35180 91420
rect 35018 91366 35020 91418
rect 35082 91366 35094 91418
rect 35156 91366 35158 91418
rect 34996 91364 35020 91366
rect 35076 91364 35100 91366
rect 35156 91364 35180 91366
rect 34940 91344 35236 91364
rect 34940 90332 35236 90352
rect 34996 90330 35020 90332
rect 35076 90330 35100 90332
rect 35156 90330 35180 90332
rect 35018 90278 35020 90330
rect 35082 90278 35094 90330
rect 35156 90278 35158 90330
rect 34996 90276 35020 90278
rect 35076 90276 35100 90278
rect 35156 90276 35180 90278
rect 34940 90256 35236 90276
rect 34940 89244 35236 89264
rect 34996 89242 35020 89244
rect 35076 89242 35100 89244
rect 35156 89242 35180 89244
rect 35018 89190 35020 89242
rect 35082 89190 35094 89242
rect 35156 89190 35158 89242
rect 34996 89188 35020 89190
rect 35076 89188 35100 89190
rect 35156 89188 35180 89190
rect 34940 89168 35236 89188
rect 34940 88156 35236 88176
rect 34996 88154 35020 88156
rect 35076 88154 35100 88156
rect 35156 88154 35180 88156
rect 35018 88102 35020 88154
rect 35082 88102 35094 88154
rect 35156 88102 35158 88154
rect 34996 88100 35020 88102
rect 35076 88100 35100 88102
rect 35156 88100 35180 88102
rect 34940 88080 35236 88100
rect 34940 87068 35236 87088
rect 34996 87066 35020 87068
rect 35076 87066 35100 87068
rect 35156 87066 35180 87068
rect 35018 87014 35020 87066
rect 35082 87014 35094 87066
rect 35156 87014 35158 87066
rect 34996 87012 35020 87014
rect 35076 87012 35100 87014
rect 35156 87012 35180 87014
rect 34940 86992 35236 87012
rect 34940 85980 35236 86000
rect 34996 85978 35020 85980
rect 35076 85978 35100 85980
rect 35156 85978 35180 85980
rect 35018 85926 35020 85978
rect 35082 85926 35094 85978
rect 35156 85926 35158 85978
rect 34996 85924 35020 85926
rect 35076 85924 35100 85926
rect 35156 85924 35180 85926
rect 34940 85904 35236 85924
rect 34940 84892 35236 84912
rect 34996 84890 35020 84892
rect 35076 84890 35100 84892
rect 35156 84890 35180 84892
rect 35018 84838 35020 84890
rect 35082 84838 35094 84890
rect 35156 84838 35158 84890
rect 34996 84836 35020 84838
rect 35076 84836 35100 84838
rect 35156 84836 35180 84838
rect 34940 84816 35236 84836
rect 34940 83804 35236 83824
rect 34996 83802 35020 83804
rect 35076 83802 35100 83804
rect 35156 83802 35180 83804
rect 35018 83750 35020 83802
rect 35082 83750 35094 83802
rect 35156 83750 35158 83802
rect 34996 83748 35020 83750
rect 35076 83748 35100 83750
rect 35156 83748 35180 83750
rect 34940 83728 35236 83748
rect 34940 82716 35236 82736
rect 34996 82714 35020 82716
rect 35076 82714 35100 82716
rect 35156 82714 35180 82716
rect 35018 82662 35020 82714
rect 35082 82662 35094 82714
rect 35156 82662 35158 82714
rect 34996 82660 35020 82662
rect 35076 82660 35100 82662
rect 35156 82660 35180 82662
rect 34940 82640 35236 82660
rect 34940 81628 35236 81648
rect 34996 81626 35020 81628
rect 35076 81626 35100 81628
rect 35156 81626 35180 81628
rect 35018 81574 35020 81626
rect 35082 81574 35094 81626
rect 35156 81574 35158 81626
rect 34996 81572 35020 81574
rect 35076 81572 35100 81574
rect 35156 81572 35180 81574
rect 34940 81552 35236 81572
rect 34940 80540 35236 80560
rect 34996 80538 35020 80540
rect 35076 80538 35100 80540
rect 35156 80538 35180 80540
rect 35018 80486 35020 80538
rect 35082 80486 35094 80538
rect 35156 80486 35158 80538
rect 34996 80484 35020 80486
rect 35076 80484 35100 80486
rect 35156 80484 35180 80486
rect 34940 80464 35236 80484
rect 34940 79452 35236 79472
rect 34996 79450 35020 79452
rect 35076 79450 35100 79452
rect 35156 79450 35180 79452
rect 35018 79398 35020 79450
rect 35082 79398 35094 79450
rect 35156 79398 35158 79450
rect 34996 79396 35020 79398
rect 35076 79396 35100 79398
rect 35156 79396 35180 79398
rect 34940 79376 35236 79396
rect 34940 78364 35236 78384
rect 34996 78362 35020 78364
rect 35076 78362 35100 78364
rect 35156 78362 35180 78364
rect 35018 78310 35020 78362
rect 35082 78310 35094 78362
rect 35156 78310 35158 78362
rect 34996 78308 35020 78310
rect 35076 78308 35100 78310
rect 35156 78308 35180 78310
rect 34940 78288 35236 78308
rect 34940 77276 35236 77296
rect 34996 77274 35020 77276
rect 35076 77274 35100 77276
rect 35156 77274 35180 77276
rect 35018 77222 35020 77274
rect 35082 77222 35094 77274
rect 35156 77222 35158 77274
rect 34996 77220 35020 77222
rect 35076 77220 35100 77222
rect 35156 77220 35180 77222
rect 34940 77200 35236 77220
rect 34940 76188 35236 76208
rect 34996 76186 35020 76188
rect 35076 76186 35100 76188
rect 35156 76186 35180 76188
rect 35018 76134 35020 76186
rect 35082 76134 35094 76186
rect 35156 76134 35158 76186
rect 34996 76132 35020 76134
rect 35076 76132 35100 76134
rect 35156 76132 35180 76134
rect 34940 76112 35236 76132
rect 34940 75100 35236 75120
rect 34996 75098 35020 75100
rect 35076 75098 35100 75100
rect 35156 75098 35180 75100
rect 35018 75046 35020 75098
rect 35082 75046 35094 75098
rect 35156 75046 35158 75098
rect 34996 75044 35020 75046
rect 35076 75044 35100 75046
rect 35156 75044 35180 75046
rect 34940 75024 35236 75044
rect 34940 74012 35236 74032
rect 34996 74010 35020 74012
rect 35076 74010 35100 74012
rect 35156 74010 35180 74012
rect 35018 73958 35020 74010
rect 35082 73958 35094 74010
rect 35156 73958 35158 74010
rect 34996 73956 35020 73958
rect 35076 73956 35100 73958
rect 35156 73956 35180 73958
rect 34940 73936 35236 73956
rect 34940 72924 35236 72944
rect 34996 72922 35020 72924
rect 35076 72922 35100 72924
rect 35156 72922 35180 72924
rect 35018 72870 35020 72922
rect 35082 72870 35094 72922
rect 35156 72870 35158 72922
rect 34996 72868 35020 72870
rect 35076 72868 35100 72870
rect 35156 72868 35180 72870
rect 34940 72848 35236 72868
rect 34940 71836 35236 71856
rect 34996 71834 35020 71836
rect 35076 71834 35100 71836
rect 35156 71834 35180 71836
rect 35018 71782 35020 71834
rect 35082 71782 35094 71834
rect 35156 71782 35158 71834
rect 34996 71780 35020 71782
rect 35076 71780 35100 71782
rect 35156 71780 35180 71782
rect 34940 71760 35236 71780
rect 34940 70748 35236 70768
rect 34996 70746 35020 70748
rect 35076 70746 35100 70748
rect 35156 70746 35180 70748
rect 35018 70694 35020 70746
rect 35082 70694 35094 70746
rect 35156 70694 35158 70746
rect 34996 70692 35020 70694
rect 35076 70692 35100 70694
rect 35156 70692 35180 70694
rect 34940 70672 35236 70692
rect 34940 69660 35236 69680
rect 34996 69658 35020 69660
rect 35076 69658 35100 69660
rect 35156 69658 35180 69660
rect 35018 69606 35020 69658
rect 35082 69606 35094 69658
rect 35156 69606 35158 69658
rect 34996 69604 35020 69606
rect 35076 69604 35100 69606
rect 35156 69604 35180 69606
rect 34940 69584 35236 69604
rect 34940 68572 35236 68592
rect 34996 68570 35020 68572
rect 35076 68570 35100 68572
rect 35156 68570 35180 68572
rect 35018 68518 35020 68570
rect 35082 68518 35094 68570
rect 35156 68518 35158 68570
rect 34996 68516 35020 68518
rect 35076 68516 35100 68518
rect 35156 68516 35180 68518
rect 34940 68496 35236 68516
rect 34940 67484 35236 67504
rect 34996 67482 35020 67484
rect 35076 67482 35100 67484
rect 35156 67482 35180 67484
rect 35018 67430 35020 67482
rect 35082 67430 35094 67482
rect 35156 67430 35158 67482
rect 34996 67428 35020 67430
rect 35076 67428 35100 67430
rect 35156 67428 35180 67430
rect 34940 67408 35236 67428
rect 34940 66396 35236 66416
rect 34996 66394 35020 66396
rect 35076 66394 35100 66396
rect 35156 66394 35180 66396
rect 35018 66342 35020 66394
rect 35082 66342 35094 66394
rect 35156 66342 35158 66394
rect 34996 66340 35020 66342
rect 35076 66340 35100 66342
rect 35156 66340 35180 66342
rect 34940 66320 35236 66340
rect 34940 65308 35236 65328
rect 34996 65306 35020 65308
rect 35076 65306 35100 65308
rect 35156 65306 35180 65308
rect 35018 65254 35020 65306
rect 35082 65254 35094 65306
rect 35156 65254 35158 65306
rect 34996 65252 35020 65254
rect 35076 65252 35100 65254
rect 35156 65252 35180 65254
rect 34940 65232 35236 65252
rect 34940 64220 35236 64240
rect 34996 64218 35020 64220
rect 35076 64218 35100 64220
rect 35156 64218 35180 64220
rect 35018 64166 35020 64218
rect 35082 64166 35094 64218
rect 35156 64166 35158 64218
rect 34996 64164 35020 64166
rect 35076 64164 35100 64166
rect 35156 64164 35180 64166
rect 34940 64144 35236 64164
rect 34940 63132 35236 63152
rect 34996 63130 35020 63132
rect 35076 63130 35100 63132
rect 35156 63130 35180 63132
rect 35018 63078 35020 63130
rect 35082 63078 35094 63130
rect 35156 63078 35158 63130
rect 34996 63076 35020 63078
rect 35076 63076 35100 63078
rect 35156 63076 35180 63078
rect 34940 63056 35236 63076
rect 34940 62044 35236 62064
rect 34996 62042 35020 62044
rect 35076 62042 35100 62044
rect 35156 62042 35180 62044
rect 35018 61990 35020 62042
rect 35082 61990 35094 62042
rect 35156 61990 35158 62042
rect 34996 61988 35020 61990
rect 35076 61988 35100 61990
rect 35156 61988 35180 61990
rect 34940 61968 35236 61988
rect 34940 60956 35236 60976
rect 34996 60954 35020 60956
rect 35076 60954 35100 60956
rect 35156 60954 35180 60956
rect 35018 60902 35020 60954
rect 35082 60902 35094 60954
rect 35156 60902 35158 60954
rect 34996 60900 35020 60902
rect 35076 60900 35100 60902
rect 35156 60900 35180 60902
rect 34940 60880 35236 60900
rect 34940 59868 35236 59888
rect 34996 59866 35020 59868
rect 35076 59866 35100 59868
rect 35156 59866 35180 59868
rect 35018 59814 35020 59866
rect 35082 59814 35094 59866
rect 35156 59814 35158 59866
rect 34996 59812 35020 59814
rect 35076 59812 35100 59814
rect 35156 59812 35180 59814
rect 34940 59792 35236 59812
rect 34940 58780 35236 58800
rect 34996 58778 35020 58780
rect 35076 58778 35100 58780
rect 35156 58778 35180 58780
rect 35018 58726 35020 58778
rect 35082 58726 35094 58778
rect 35156 58726 35158 58778
rect 34996 58724 35020 58726
rect 35076 58724 35100 58726
rect 35156 58724 35180 58726
rect 34940 58704 35236 58724
rect 34940 57692 35236 57712
rect 34996 57690 35020 57692
rect 35076 57690 35100 57692
rect 35156 57690 35180 57692
rect 35018 57638 35020 57690
rect 35082 57638 35094 57690
rect 35156 57638 35158 57690
rect 34996 57636 35020 57638
rect 35076 57636 35100 57638
rect 35156 57636 35180 57638
rect 34940 57616 35236 57636
rect 34940 56604 35236 56624
rect 34996 56602 35020 56604
rect 35076 56602 35100 56604
rect 35156 56602 35180 56604
rect 35018 56550 35020 56602
rect 35082 56550 35094 56602
rect 35156 56550 35158 56602
rect 34996 56548 35020 56550
rect 35076 56548 35100 56550
rect 35156 56548 35180 56550
rect 34940 56528 35236 56548
rect 34940 55516 35236 55536
rect 34996 55514 35020 55516
rect 35076 55514 35100 55516
rect 35156 55514 35180 55516
rect 35018 55462 35020 55514
rect 35082 55462 35094 55514
rect 35156 55462 35158 55514
rect 34996 55460 35020 55462
rect 35076 55460 35100 55462
rect 35156 55460 35180 55462
rect 34940 55440 35236 55460
rect 34940 54428 35236 54448
rect 34996 54426 35020 54428
rect 35076 54426 35100 54428
rect 35156 54426 35180 54428
rect 35018 54374 35020 54426
rect 35082 54374 35094 54426
rect 35156 54374 35158 54426
rect 34996 54372 35020 54374
rect 35076 54372 35100 54374
rect 35156 54372 35180 54374
rect 34940 54352 35236 54372
rect 34940 53340 35236 53360
rect 34996 53338 35020 53340
rect 35076 53338 35100 53340
rect 35156 53338 35180 53340
rect 35018 53286 35020 53338
rect 35082 53286 35094 53338
rect 35156 53286 35158 53338
rect 34996 53284 35020 53286
rect 35076 53284 35100 53286
rect 35156 53284 35180 53286
rect 34940 53264 35236 53284
rect 34940 52252 35236 52272
rect 34996 52250 35020 52252
rect 35076 52250 35100 52252
rect 35156 52250 35180 52252
rect 35018 52198 35020 52250
rect 35082 52198 35094 52250
rect 35156 52198 35158 52250
rect 34996 52196 35020 52198
rect 35076 52196 35100 52198
rect 35156 52196 35180 52198
rect 34940 52176 35236 52196
rect 34940 51164 35236 51184
rect 34996 51162 35020 51164
rect 35076 51162 35100 51164
rect 35156 51162 35180 51164
rect 35018 51110 35020 51162
rect 35082 51110 35094 51162
rect 35156 51110 35158 51162
rect 34996 51108 35020 51110
rect 35076 51108 35100 51110
rect 35156 51108 35180 51110
rect 34940 51088 35236 51108
rect 34940 50076 35236 50096
rect 34996 50074 35020 50076
rect 35076 50074 35100 50076
rect 35156 50074 35180 50076
rect 35018 50022 35020 50074
rect 35082 50022 35094 50074
rect 35156 50022 35158 50074
rect 34996 50020 35020 50022
rect 35076 50020 35100 50022
rect 35156 50020 35180 50022
rect 34940 50000 35236 50020
rect 34940 48988 35236 49008
rect 34996 48986 35020 48988
rect 35076 48986 35100 48988
rect 35156 48986 35180 48988
rect 35018 48934 35020 48986
rect 35082 48934 35094 48986
rect 35156 48934 35158 48986
rect 34996 48932 35020 48934
rect 35076 48932 35100 48934
rect 35156 48932 35180 48934
rect 34940 48912 35236 48932
rect 34940 47900 35236 47920
rect 34996 47898 35020 47900
rect 35076 47898 35100 47900
rect 35156 47898 35180 47900
rect 35018 47846 35020 47898
rect 35082 47846 35094 47898
rect 35156 47846 35158 47898
rect 34996 47844 35020 47846
rect 35076 47844 35100 47846
rect 35156 47844 35180 47846
rect 34940 47824 35236 47844
rect 34940 46812 35236 46832
rect 34996 46810 35020 46812
rect 35076 46810 35100 46812
rect 35156 46810 35180 46812
rect 35018 46758 35020 46810
rect 35082 46758 35094 46810
rect 35156 46758 35158 46810
rect 34996 46756 35020 46758
rect 35076 46756 35100 46758
rect 35156 46756 35180 46758
rect 34940 46736 35236 46756
rect 34940 45724 35236 45744
rect 34996 45722 35020 45724
rect 35076 45722 35100 45724
rect 35156 45722 35180 45724
rect 35018 45670 35020 45722
rect 35082 45670 35094 45722
rect 35156 45670 35158 45722
rect 34996 45668 35020 45670
rect 35076 45668 35100 45670
rect 35156 45668 35180 45670
rect 34940 45648 35236 45668
rect 34940 44636 35236 44656
rect 34996 44634 35020 44636
rect 35076 44634 35100 44636
rect 35156 44634 35180 44636
rect 35018 44582 35020 44634
rect 35082 44582 35094 44634
rect 35156 44582 35158 44634
rect 34996 44580 35020 44582
rect 35076 44580 35100 44582
rect 35156 44580 35180 44582
rect 34940 44560 35236 44580
rect 34940 43548 35236 43568
rect 34996 43546 35020 43548
rect 35076 43546 35100 43548
rect 35156 43546 35180 43548
rect 35018 43494 35020 43546
rect 35082 43494 35094 43546
rect 35156 43494 35158 43546
rect 34996 43492 35020 43494
rect 35076 43492 35100 43494
rect 35156 43492 35180 43494
rect 34940 43472 35236 43492
rect 34940 42460 35236 42480
rect 34996 42458 35020 42460
rect 35076 42458 35100 42460
rect 35156 42458 35180 42460
rect 35018 42406 35020 42458
rect 35082 42406 35094 42458
rect 35156 42406 35158 42458
rect 34996 42404 35020 42406
rect 35076 42404 35100 42406
rect 35156 42404 35180 42406
rect 34940 42384 35236 42404
rect 34940 41372 35236 41392
rect 34996 41370 35020 41372
rect 35076 41370 35100 41372
rect 35156 41370 35180 41372
rect 35018 41318 35020 41370
rect 35082 41318 35094 41370
rect 35156 41318 35158 41370
rect 34996 41316 35020 41318
rect 35076 41316 35100 41318
rect 35156 41316 35180 41318
rect 34940 41296 35236 41316
rect 34940 40284 35236 40304
rect 34996 40282 35020 40284
rect 35076 40282 35100 40284
rect 35156 40282 35180 40284
rect 35018 40230 35020 40282
rect 35082 40230 35094 40282
rect 35156 40230 35158 40282
rect 34996 40228 35020 40230
rect 35076 40228 35100 40230
rect 35156 40228 35180 40230
rect 34940 40208 35236 40228
rect 34940 39196 35236 39216
rect 34996 39194 35020 39196
rect 35076 39194 35100 39196
rect 35156 39194 35180 39196
rect 35018 39142 35020 39194
rect 35082 39142 35094 39194
rect 35156 39142 35158 39194
rect 34996 39140 35020 39142
rect 35076 39140 35100 39142
rect 35156 39140 35180 39142
rect 34940 39120 35236 39140
rect 34940 38108 35236 38128
rect 34996 38106 35020 38108
rect 35076 38106 35100 38108
rect 35156 38106 35180 38108
rect 35018 38054 35020 38106
rect 35082 38054 35094 38106
rect 35156 38054 35158 38106
rect 34996 38052 35020 38054
rect 35076 38052 35100 38054
rect 35156 38052 35180 38054
rect 34940 38032 35236 38052
rect 34940 37020 35236 37040
rect 34996 37018 35020 37020
rect 35076 37018 35100 37020
rect 35156 37018 35180 37020
rect 35018 36966 35020 37018
rect 35082 36966 35094 37018
rect 35156 36966 35158 37018
rect 34996 36964 35020 36966
rect 35076 36964 35100 36966
rect 35156 36964 35180 36966
rect 34940 36944 35236 36964
rect 34940 35932 35236 35952
rect 34996 35930 35020 35932
rect 35076 35930 35100 35932
rect 35156 35930 35180 35932
rect 35018 35878 35020 35930
rect 35082 35878 35094 35930
rect 35156 35878 35158 35930
rect 34996 35876 35020 35878
rect 35076 35876 35100 35878
rect 35156 35876 35180 35878
rect 34940 35856 35236 35876
rect 34940 34844 35236 34864
rect 34996 34842 35020 34844
rect 35076 34842 35100 34844
rect 35156 34842 35180 34844
rect 35018 34790 35020 34842
rect 35082 34790 35094 34842
rect 35156 34790 35158 34842
rect 34996 34788 35020 34790
rect 35076 34788 35100 34790
rect 35156 34788 35180 34790
rect 34940 34768 35236 34788
rect 34940 33756 35236 33776
rect 34996 33754 35020 33756
rect 35076 33754 35100 33756
rect 35156 33754 35180 33756
rect 35018 33702 35020 33754
rect 35082 33702 35094 33754
rect 35156 33702 35158 33754
rect 34996 33700 35020 33702
rect 35076 33700 35100 33702
rect 35156 33700 35180 33702
rect 34940 33680 35236 33700
rect 34940 32668 35236 32688
rect 34996 32666 35020 32668
rect 35076 32666 35100 32668
rect 35156 32666 35180 32668
rect 35018 32614 35020 32666
rect 35082 32614 35094 32666
rect 35156 32614 35158 32666
rect 34996 32612 35020 32614
rect 35076 32612 35100 32614
rect 35156 32612 35180 32614
rect 34940 32592 35236 32612
rect 34940 31580 35236 31600
rect 34996 31578 35020 31580
rect 35076 31578 35100 31580
rect 35156 31578 35180 31580
rect 35018 31526 35020 31578
rect 35082 31526 35094 31578
rect 35156 31526 35158 31578
rect 34996 31524 35020 31526
rect 35076 31524 35100 31526
rect 35156 31524 35180 31526
rect 34940 31504 35236 31524
rect 34940 30492 35236 30512
rect 34996 30490 35020 30492
rect 35076 30490 35100 30492
rect 35156 30490 35180 30492
rect 35018 30438 35020 30490
rect 35082 30438 35094 30490
rect 35156 30438 35158 30490
rect 34996 30436 35020 30438
rect 35076 30436 35100 30438
rect 35156 30436 35180 30438
rect 34940 30416 35236 30436
rect 34940 29404 35236 29424
rect 34996 29402 35020 29404
rect 35076 29402 35100 29404
rect 35156 29402 35180 29404
rect 35018 29350 35020 29402
rect 35082 29350 35094 29402
rect 35156 29350 35158 29402
rect 34996 29348 35020 29350
rect 35076 29348 35100 29350
rect 35156 29348 35180 29350
rect 34940 29328 35236 29348
rect 34940 28316 35236 28336
rect 34996 28314 35020 28316
rect 35076 28314 35100 28316
rect 35156 28314 35180 28316
rect 35018 28262 35020 28314
rect 35082 28262 35094 28314
rect 35156 28262 35158 28314
rect 34996 28260 35020 28262
rect 35076 28260 35100 28262
rect 35156 28260 35180 28262
rect 34940 28240 35236 28260
rect 34940 27228 35236 27248
rect 34996 27226 35020 27228
rect 35076 27226 35100 27228
rect 35156 27226 35180 27228
rect 35018 27174 35020 27226
rect 35082 27174 35094 27226
rect 35156 27174 35158 27226
rect 34996 27172 35020 27174
rect 35076 27172 35100 27174
rect 35156 27172 35180 27174
rect 34940 27152 35236 27172
rect 34940 26140 35236 26160
rect 34996 26138 35020 26140
rect 35076 26138 35100 26140
rect 35156 26138 35180 26140
rect 35018 26086 35020 26138
rect 35082 26086 35094 26138
rect 35156 26086 35158 26138
rect 34996 26084 35020 26086
rect 35076 26084 35100 26086
rect 35156 26084 35180 26086
rect 34940 26064 35236 26084
rect 34940 25052 35236 25072
rect 34996 25050 35020 25052
rect 35076 25050 35100 25052
rect 35156 25050 35180 25052
rect 35018 24998 35020 25050
rect 35082 24998 35094 25050
rect 35156 24998 35158 25050
rect 34996 24996 35020 24998
rect 35076 24996 35100 24998
rect 35156 24996 35180 24998
rect 34940 24976 35236 24996
rect 36832 24274 36860 117098
rect 39776 116346 39804 117098
rect 39764 116340 39816 116346
rect 39764 116282 39816 116288
rect 35900 24268 35952 24274
rect 35900 24210 35952 24216
rect 36820 24268 36872 24274
rect 36820 24210 36872 24216
rect 34940 23964 35236 23984
rect 34996 23962 35020 23964
rect 35076 23962 35100 23964
rect 35156 23962 35180 23964
rect 35018 23910 35020 23962
rect 35082 23910 35094 23962
rect 35156 23910 35158 23962
rect 34996 23908 35020 23910
rect 35076 23908 35100 23910
rect 35156 23908 35180 23910
rect 34940 23888 35236 23908
rect 34940 22876 35236 22896
rect 34996 22874 35020 22876
rect 35076 22874 35100 22876
rect 35156 22874 35180 22876
rect 35018 22822 35020 22874
rect 35082 22822 35094 22874
rect 35156 22822 35158 22874
rect 34996 22820 35020 22822
rect 35076 22820 35100 22822
rect 35156 22820 35180 22822
rect 34940 22800 35236 22820
rect 33416 22432 33468 22438
rect 33416 22374 33468 22380
rect 35256 22432 35308 22438
rect 35256 22374 35308 22380
rect 32140 22066 32260 22094
rect 32036 21072 32088 21078
rect 32036 21014 32088 21020
rect 31944 19916 31996 19922
rect 31944 19858 31996 19864
rect 31956 18222 31984 19858
rect 31944 18216 31996 18222
rect 31944 18158 31996 18164
rect 31852 18148 31904 18154
rect 31852 18090 31904 18096
rect 31864 15706 31892 18090
rect 31944 16176 31996 16182
rect 31944 16118 31996 16124
rect 31852 15700 31904 15706
rect 31852 15642 31904 15648
rect 31760 14544 31812 14550
rect 31760 14486 31812 14492
rect 31956 13938 31984 16118
rect 32048 15638 32076 21014
rect 32128 18692 32180 18698
rect 32128 18634 32180 18640
rect 32140 16794 32168 18634
rect 32128 16788 32180 16794
rect 32128 16730 32180 16736
rect 32140 16046 32168 16730
rect 32232 16658 32260 22066
rect 33232 20460 33284 20466
rect 33232 20402 33284 20408
rect 33048 18284 33100 18290
rect 33048 18226 33100 18232
rect 32404 17536 32456 17542
rect 32404 17478 32456 17484
rect 32416 16658 32444 17478
rect 32220 16652 32272 16658
rect 32220 16594 32272 16600
rect 32404 16652 32456 16658
rect 32404 16594 32456 16600
rect 32128 16040 32180 16046
rect 32128 15982 32180 15988
rect 32036 15632 32088 15638
rect 32036 15574 32088 15580
rect 31944 13932 31996 13938
rect 31944 13874 31996 13880
rect 31668 13864 31720 13870
rect 31668 13806 31720 13812
rect 31680 10198 31708 13806
rect 32048 12986 32076 15574
rect 32036 12980 32088 12986
rect 32036 12922 32088 12928
rect 31668 10192 31720 10198
rect 31668 10134 31720 10140
rect 32048 9518 32076 12922
rect 32036 9512 32088 9518
rect 32036 9454 32088 9460
rect 31668 8492 31720 8498
rect 31668 8434 31720 8440
rect 31576 8084 31628 8090
rect 31576 8026 31628 8032
rect 31588 7478 31616 8026
rect 31680 7954 31708 8434
rect 31852 8424 31904 8430
rect 31852 8366 31904 8372
rect 31864 8022 31892 8366
rect 31944 8356 31996 8362
rect 31944 8298 31996 8304
rect 31852 8016 31904 8022
rect 31852 7958 31904 7964
rect 31668 7948 31720 7954
rect 31668 7890 31720 7896
rect 31576 7472 31628 7478
rect 31576 7414 31628 7420
rect 31128 7126 31524 7154
rect 31024 6928 31076 6934
rect 31024 6870 31076 6876
rect 31024 6792 31076 6798
rect 31024 6734 31076 6740
rect 31036 6254 31064 6734
rect 31024 6248 31076 6254
rect 31024 6190 31076 6196
rect 31128 6202 31156 7126
rect 31298 7032 31354 7041
rect 31298 6967 31354 6976
rect 31208 6928 31260 6934
rect 31208 6870 31260 6876
rect 31220 6390 31248 6870
rect 31312 6730 31340 6967
rect 31484 6928 31536 6934
rect 31404 6888 31484 6916
rect 31300 6724 31352 6730
rect 31300 6666 31352 6672
rect 31404 6662 31432 6888
rect 31760 6928 31812 6934
rect 31484 6870 31536 6876
rect 31680 6888 31760 6916
rect 31392 6656 31444 6662
rect 31392 6598 31444 6604
rect 31208 6384 31260 6390
rect 31208 6326 31260 6332
rect 31128 6186 31248 6202
rect 31128 6180 31260 6186
rect 31128 6174 31208 6180
rect 31208 6122 31260 6128
rect 31680 6089 31708 6888
rect 31760 6870 31812 6876
rect 31758 6760 31814 6769
rect 31758 6695 31814 6704
rect 31772 6458 31800 6695
rect 31760 6452 31812 6458
rect 31760 6394 31812 6400
rect 31666 6080 31722 6089
rect 31666 6015 31722 6024
rect 31576 5908 31628 5914
rect 31576 5850 31628 5856
rect 31588 5710 31616 5850
rect 31576 5704 31628 5710
rect 31576 5646 31628 5652
rect 30932 5364 30984 5370
rect 30932 5306 30984 5312
rect 31576 5296 31628 5302
rect 31680 5284 31708 6015
rect 31956 5914 31984 8298
rect 32140 7546 32168 15982
rect 32232 15978 32260 16594
rect 32416 16250 32444 16594
rect 32404 16244 32456 16250
rect 32404 16186 32456 16192
rect 32220 15972 32272 15978
rect 32220 15914 32272 15920
rect 32416 15910 32444 16186
rect 32404 15904 32456 15910
rect 32404 15846 32456 15852
rect 32496 15088 32548 15094
rect 32496 15030 32548 15036
rect 32220 14816 32272 14822
rect 32220 14758 32272 14764
rect 32232 13530 32260 14758
rect 32220 13524 32272 13530
rect 32220 13466 32272 13472
rect 32232 7834 32260 13466
rect 32508 8129 32536 15030
rect 33060 14618 33088 18226
rect 33140 18216 33192 18222
rect 33140 18158 33192 18164
rect 33048 14612 33100 14618
rect 33048 14554 33100 14560
rect 33152 14482 33180 18158
rect 33140 14476 33192 14482
rect 33140 14418 33192 14424
rect 33140 14272 33192 14278
rect 33140 14214 33192 14220
rect 32956 12776 33008 12782
rect 32956 12718 33008 12724
rect 32680 10260 32732 10266
rect 32680 10202 32732 10208
rect 32588 9036 32640 9042
rect 32588 8978 32640 8984
rect 32600 8430 32628 8978
rect 32588 8424 32640 8430
rect 32588 8366 32640 8372
rect 32494 8120 32550 8129
rect 32494 8055 32550 8064
rect 32508 8022 32536 8055
rect 32496 8016 32548 8022
rect 32496 7958 32548 7964
rect 32588 8016 32640 8022
rect 32588 7958 32640 7964
rect 32232 7806 32352 7834
rect 32128 7540 32180 7546
rect 32128 7482 32180 7488
rect 32324 6458 32352 7806
rect 32312 6452 32364 6458
rect 32312 6394 32364 6400
rect 32126 6352 32182 6361
rect 32126 6287 32182 6296
rect 31944 5908 31996 5914
rect 31944 5850 31996 5856
rect 31852 5704 31904 5710
rect 31850 5672 31852 5681
rect 31904 5672 31906 5681
rect 31850 5607 31906 5616
rect 31628 5256 31708 5284
rect 31576 5238 31628 5244
rect 31760 5024 31812 5030
rect 31760 4966 31812 4972
rect 31852 5024 31904 5030
rect 31852 4966 31904 4972
rect 31772 4865 31800 4966
rect 31758 4856 31814 4865
rect 31758 4791 31814 4800
rect 31668 4616 31720 4622
rect 31668 4558 31720 4564
rect 31680 4457 31708 4558
rect 31864 4457 31892 4966
rect 31666 4448 31722 4457
rect 31666 4383 31722 4392
rect 31850 4448 31906 4457
rect 31850 4383 31906 4392
rect 31956 4078 31984 5850
rect 32036 5840 32088 5846
rect 32036 5782 32088 5788
rect 32048 5574 32076 5782
rect 32036 5568 32088 5574
rect 32036 5510 32088 5516
rect 32048 5234 32076 5510
rect 32036 5228 32088 5234
rect 32036 5170 32088 5176
rect 31944 4072 31996 4078
rect 31944 4014 31996 4020
rect 31300 3596 31352 3602
rect 31300 3538 31352 3544
rect 30932 2848 30984 2854
rect 30932 2790 30984 2796
rect 30840 2304 30892 2310
rect 30840 2246 30892 2252
rect 30944 800 30972 2790
rect 31116 2304 31168 2310
rect 31116 2246 31168 2252
rect 31128 1630 31156 2246
rect 31116 1624 31168 1630
rect 31116 1566 31168 1572
rect 31312 800 31340 3538
rect 31576 3120 31628 3126
rect 31576 3062 31628 3068
rect 29736 672 29788 678
rect 29736 614 29788 620
rect 29826 0 29882 800
rect 30194 0 30250 800
rect 30562 0 30618 800
rect 30930 0 30986 800
rect 31298 0 31354 800
rect 31588 542 31616 3062
rect 32036 2848 32088 2854
rect 32036 2790 32088 2796
rect 31668 2508 31720 2514
rect 31668 2450 31720 2456
rect 31680 800 31708 2450
rect 32048 800 32076 2790
rect 32140 2582 32168 6287
rect 32600 4842 32628 7958
rect 32692 6730 32720 10202
rect 32968 10198 32996 12718
rect 32956 10192 33008 10198
rect 32956 10134 33008 10140
rect 33048 8424 33100 8430
rect 33048 8366 33100 8372
rect 32954 8120 33010 8129
rect 32954 8055 33010 8064
rect 32968 8022 32996 8055
rect 32956 8016 33008 8022
rect 32770 7984 32826 7993
rect 32956 7958 33008 7964
rect 32770 7919 32826 7928
rect 32864 7948 32916 7954
rect 32784 7410 32812 7919
rect 32864 7890 32916 7896
rect 32772 7404 32824 7410
rect 32772 7346 32824 7352
rect 32680 6724 32732 6730
rect 32680 6666 32732 6672
rect 32680 6316 32732 6322
rect 32680 6258 32732 6264
rect 32692 5574 32720 6258
rect 32876 6089 32904 7890
rect 33060 7410 33088 8366
rect 33048 7404 33100 7410
rect 33048 7346 33100 7352
rect 33048 7200 33100 7206
rect 33048 7142 33100 7148
rect 32956 6860 33008 6866
rect 32956 6802 33008 6808
rect 32862 6080 32918 6089
rect 32862 6015 32918 6024
rect 32680 5568 32732 5574
rect 32680 5510 32732 5516
rect 32324 4814 32628 4842
rect 32324 4282 32352 4814
rect 32404 4616 32456 4622
rect 32404 4558 32456 4564
rect 32416 4282 32444 4558
rect 32312 4276 32364 4282
rect 32312 4218 32364 4224
rect 32404 4276 32456 4282
rect 32404 4218 32456 4224
rect 32404 3596 32456 3602
rect 32404 3538 32456 3544
rect 32128 2576 32180 2582
rect 32128 2518 32180 2524
rect 32416 800 32444 3538
rect 32496 2508 32548 2514
rect 32496 2450 32548 2456
rect 32772 2508 32824 2514
rect 32772 2450 32824 2456
rect 32508 1834 32536 2450
rect 32496 1828 32548 1834
rect 32496 1770 32548 1776
rect 32784 800 32812 2450
rect 32968 1222 32996 6802
rect 33060 6712 33088 7142
rect 33152 6866 33180 14214
rect 33244 13394 33272 20402
rect 33428 18834 33456 22374
rect 34940 21788 35236 21808
rect 34996 21786 35020 21788
rect 35076 21786 35100 21788
rect 35156 21786 35180 21788
rect 35018 21734 35020 21786
rect 35082 21734 35094 21786
rect 35156 21734 35158 21786
rect 34996 21732 35020 21734
rect 35076 21732 35100 21734
rect 35156 21732 35180 21734
rect 34940 21712 35236 21732
rect 34940 20700 35236 20720
rect 34996 20698 35020 20700
rect 35076 20698 35100 20700
rect 35156 20698 35180 20700
rect 35018 20646 35020 20698
rect 35082 20646 35094 20698
rect 35156 20646 35158 20698
rect 34996 20644 35020 20646
rect 35076 20644 35100 20646
rect 35156 20644 35180 20646
rect 34940 20624 35236 20644
rect 34940 19612 35236 19632
rect 34996 19610 35020 19612
rect 35076 19610 35100 19612
rect 35156 19610 35180 19612
rect 35018 19558 35020 19610
rect 35082 19558 35094 19610
rect 35156 19558 35158 19610
rect 34996 19556 35020 19558
rect 35076 19556 35100 19558
rect 35156 19556 35180 19558
rect 34940 19536 35236 19556
rect 35268 19310 35296 22374
rect 35256 19304 35308 19310
rect 35256 19246 35308 19252
rect 35808 19304 35860 19310
rect 35808 19246 35860 19252
rect 33416 18828 33468 18834
rect 33416 18770 33468 18776
rect 35348 18828 35400 18834
rect 35348 18770 35400 18776
rect 34940 18524 35236 18544
rect 34996 18522 35020 18524
rect 35076 18522 35100 18524
rect 35156 18522 35180 18524
rect 35018 18470 35020 18522
rect 35082 18470 35094 18522
rect 35156 18470 35158 18522
rect 34996 18468 35020 18470
rect 35076 18468 35100 18470
rect 35156 18468 35180 18470
rect 34940 18448 35236 18468
rect 34940 17436 35236 17456
rect 34996 17434 35020 17436
rect 35076 17434 35100 17436
rect 35156 17434 35180 17436
rect 35018 17382 35020 17434
rect 35082 17382 35094 17434
rect 35156 17382 35158 17434
rect 34996 17380 35020 17382
rect 35076 17380 35100 17382
rect 35156 17380 35180 17382
rect 34940 17360 35236 17380
rect 35256 17128 35308 17134
rect 35256 17070 35308 17076
rect 33692 16788 33744 16794
rect 33692 16730 33744 16736
rect 33704 15570 33732 16730
rect 34940 16348 35236 16368
rect 34996 16346 35020 16348
rect 35076 16346 35100 16348
rect 35156 16346 35180 16348
rect 35018 16294 35020 16346
rect 35082 16294 35094 16346
rect 35156 16294 35158 16346
rect 34996 16292 35020 16294
rect 35076 16292 35100 16294
rect 35156 16292 35180 16294
rect 34940 16272 35236 16292
rect 35268 16250 35296 17070
rect 34520 16244 34572 16250
rect 34520 16186 34572 16192
rect 35256 16244 35308 16250
rect 35256 16186 35308 16192
rect 34532 15570 34560 16186
rect 33692 15564 33744 15570
rect 33692 15506 33744 15512
rect 34520 15564 34572 15570
rect 34520 15506 34572 15512
rect 34796 15360 34848 15366
rect 34796 15302 34848 15308
rect 33508 14952 33560 14958
rect 33508 14894 33560 14900
rect 33784 14952 33836 14958
rect 33784 14894 33836 14900
rect 33232 13388 33284 13394
rect 33232 13330 33284 13336
rect 33232 13252 33284 13258
rect 33232 13194 33284 13200
rect 33244 10810 33272 13194
rect 33520 12850 33548 14894
rect 33508 12844 33560 12850
rect 33508 12786 33560 12792
rect 33324 12776 33376 12782
rect 33324 12718 33376 12724
rect 33232 10804 33284 10810
rect 33232 10746 33284 10752
rect 33336 10198 33364 12718
rect 33796 10810 33824 14894
rect 34612 14476 34664 14482
rect 34612 14418 34664 14424
rect 33968 14408 34020 14414
rect 33968 14350 34020 14356
rect 33980 13870 34008 14350
rect 34244 14340 34296 14346
rect 34244 14282 34296 14288
rect 33968 13864 34020 13870
rect 33968 13806 34020 13812
rect 33980 13394 34008 13806
rect 33968 13388 34020 13394
rect 33968 13330 34020 13336
rect 33784 10804 33836 10810
rect 33784 10746 33836 10752
rect 34256 10606 34284 14282
rect 34520 13320 34572 13326
rect 34520 13262 34572 13268
rect 34532 12374 34560 13262
rect 34624 12986 34652 14418
rect 34612 12980 34664 12986
rect 34612 12922 34664 12928
rect 34624 12866 34652 12922
rect 34624 12838 34744 12866
rect 34520 12368 34572 12374
rect 34520 12310 34572 12316
rect 33600 10600 33652 10606
rect 33600 10542 33652 10548
rect 34244 10600 34296 10606
rect 34244 10542 34296 10548
rect 33612 10266 33640 10542
rect 33784 10532 33836 10538
rect 33784 10474 33836 10480
rect 33600 10260 33652 10266
rect 33600 10202 33652 10208
rect 33324 10192 33376 10198
rect 33324 10134 33376 10140
rect 33612 10130 33640 10202
rect 33600 10124 33652 10130
rect 33600 10066 33652 10072
rect 33232 8832 33284 8838
rect 33232 8774 33284 8780
rect 33416 8832 33468 8838
rect 33416 8774 33468 8780
rect 33140 6860 33192 6866
rect 33140 6802 33192 6808
rect 33140 6724 33192 6730
rect 33060 6684 33140 6712
rect 33140 6666 33192 6672
rect 33048 6452 33100 6458
rect 33048 6394 33100 6400
rect 33060 5137 33088 6394
rect 33152 6254 33180 6666
rect 33140 6248 33192 6254
rect 33138 6216 33140 6225
rect 33192 6216 33194 6225
rect 33138 6151 33194 6160
rect 33046 5128 33102 5137
rect 33244 5114 33272 8774
rect 33428 8430 33456 8774
rect 33600 8628 33652 8634
rect 33600 8570 33652 8576
rect 33416 8424 33468 8430
rect 33416 8366 33468 8372
rect 33612 8090 33640 8570
rect 33692 8560 33744 8566
rect 33692 8502 33744 8508
rect 33600 8084 33652 8090
rect 33600 8026 33652 8032
rect 33324 7880 33376 7886
rect 33324 7822 33376 7828
rect 33336 7206 33364 7822
rect 33508 7336 33560 7342
rect 33508 7278 33560 7284
rect 33324 7200 33376 7206
rect 33324 7142 33376 7148
rect 33520 7002 33548 7278
rect 33600 7268 33652 7274
rect 33600 7210 33652 7216
rect 33324 6996 33376 7002
rect 33324 6938 33376 6944
rect 33508 6996 33560 7002
rect 33508 6938 33560 6944
rect 33336 6905 33364 6938
rect 33322 6896 33378 6905
rect 33508 6860 33560 6866
rect 33322 6831 33378 6840
rect 33428 6820 33508 6848
rect 33324 6180 33376 6186
rect 33324 6122 33376 6128
rect 33152 5098 33272 5114
rect 33046 5063 33102 5072
rect 33140 5092 33272 5098
rect 33192 5086 33272 5092
rect 33140 5034 33192 5040
rect 33140 4548 33192 4554
rect 33140 4490 33192 4496
rect 33152 3738 33180 4490
rect 33140 3732 33192 3738
rect 33140 3674 33192 3680
rect 33232 3732 33284 3738
rect 33232 3674 33284 3680
rect 33244 2990 33272 3674
rect 33232 2984 33284 2990
rect 33232 2926 33284 2932
rect 33140 2848 33192 2854
rect 33140 2790 33192 2796
rect 32956 1216 33008 1222
rect 32956 1158 33008 1164
rect 33152 800 33180 2790
rect 33336 1902 33364 6122
rect 33428 2106 33456 6820
rect 33508 6802 33560 6808
rect 33612 5556 33640 7210
rect 33704 5914 33732 8502
rect 33796 8090 33824 10474
rect 34716 10146 34744 12838
rect 34808 12442 34836 15302
rect 34940 15260 35236 15280
rect 34996 15258 35020 15260
rect 35076 15258 35100 15260
rect 35156 15258 35180 15260
rect 35018 15206 35020 15258
rect 35082 15206 35094 15258
rect 35156 15206 35158 15258
rect 34996 15204 35020 15206
rect 35076 15204 35100 15206
rect 35156 15204 35180 15206
rect 34940 15184 35236 15204
rect 35360 14890 35388 18770
rect 35820 17678 35848 19246
rect 35808 17672 35860 17678
rect 35808 17614 35860 17620
rect 35820 17202 35848 17614
rect 35808 17196 35860 17202
rect 35808 17138 35860 17144
rect 35912 17134 35940 24210
rect 41708 19310 41736 117098
rect 44376 116346 44404 117098
rect 44364 116340 44416 116346
rect 44364 116282 44416 116288
rect 47044 22094 47072 117098
rect 48976 116346 49004 117098
rect 50300 116988 50596 117008
rect 50356 116986 50380 116988
rect 50436 116986 50460 116988
rect 50516 116986 50540 116988
rect 50378 116934 50380 116986
rect 50442 116934 50454 116986
rect 50516 116934 50518 116986
rect 50356 116932 50380 116934
rect 50436 116932 50460 116934
rect 50516 116932 50540 116934
rect 50300 116912 50596 116932
rect 48964 116340 49016 116346
rect 48964 116282 49016 116288
rect 50300 115900 50596 115920
rect 50356 115898 50380 115900
rect 50436 115898 50460 115900
rect 50516 115898 50540 115900
rect 50378 115846 50380 115898
rect 50442 115846 50454 115898
rect 50516 115846 50518 115898
rect 50356 115844 50380 115846
rect 50436 115844 50460 115846
rect 50516 115844 50540 115846
rect 50300 115824 50596 115844
rect 50300 114812 50596 114832
rect 50356 114810 50380 114812
rect 50436 114810 50460 114812
rect 50516 114810 50540 114812
rect 50378 114758 50380 114810
rect 50442 114758 50454 114810
rect 50516 114758 50518 114810
rect 50356 114756 50380 114758
rect 50436 114756 50460 114758
rect 50516 114756 50540 114758
rect 50300 114736 50596 114756
rect 50300 113724 50596 113744
rect 50356 113722 50380 113724
rect 50436 113722 50460 113724
rect 50516 113722 50540 113724
rect 50378 113670 50380 113722
rect 50442 113670 50454 113722
rect 50516 113670 50518 113722
rect 50356 113668 50380 113670
rect 50436 113668 50460 113670
rect 50516 113668 50540 113670
rect 50300 113648 50596 113668
rect 50300 112636 50596 112656
rect 50356 112634 50380 112636
rect 50436 112634 50460 112636
rect 50516 112634 50540 112636
rect 50378 112582 50380 112634
rect 50442 112582 50454 112634
rect 50516 112582 50518 112634
rect 50356 112580 50380 112582
rect 50436 112580 50460 112582
rect 50516 112580 50540 112582
rect 50300 112560 50596 112580
rect 50300 111548 50596 111568
rect 50356 111546 50380 111548
rect 50436 111546 50460 111548
rect 50516 111546 50540 111548
rect 50378 111494 50380 111546
rect 50442 111494 50454 111546
rect 50516 111494 50518 111546
rect 50356 111492 50380 111494
rect 50436 111492 50460 111494
rect 50516 111492 50540 111494
rect 50300 111472 50596 111492
rect 50300 110460 50596 110480
rect 50356 110458 50380 110460
rect 50436 110458 50460 110460
rect 50516 110458 50540 110460
rect 50378 110406 50380 110458
rect 50442 110406 50454 110458
rect 50516 110406 50518 110458
rect 50356 110404 50380 110406
rect 50436 110404 50460 110406
rect 50516 110404 50540 110406
rect 50300 110384 50596 110404
rect 50300 109372 50596 109392
rect 50356 109370 50380 109372
rect 50436 109370 50460 109372
rect 50516 109370 50540 109372
rect 50378 109318 50380 109370
rect 50442 109318 50454 109370
rect 50516 109318 50518 109370
rect 50356 109316 50380 109318
rect 50436 109316 50460 109318
rect 50516 109316 50540 109318
rect 50300 109296 50596 109316
rect 50300 108284 50596 108304
rect 50356 108282 50380 108284
rect 50436 108282 50460 108284
rect 50516 108282 50540 108284
rect 50378 108230 50380 108282
rect 50442 108230 50454 108282
rect 50516 108230 50518 108282
rect 50356 108228 50380 108230
rect 50436 108228 50460 108230
rect 50516 108228 50540 108230
rect 50300 108208 50596 108228
rect 50300 107196 50596 107216
rect 50356 107194 50380 107196
rect 50436 107194 50460 107196
rect 50516 107194 50540 107196
rect 50378 107142 50380 107194
rect 50442 107142 50454 107194
rect 50516 107142 50518 107194
rect 50356 107140 50380 107142
rect 50436 107140 50460 107142
rect 50516 107140 50540 107142
rect 50300 107120 50596 107140
rect 50300 106108 50596 106128
rect 50356 106106 50380 106108
rect 50436 106106 50460 106108
rect 50516 106106 50540 106108
rect 50378 106054 50380 106106
rect 50442 106054 50454 106106
rect 50516 106054 50518 106106
rect 50356 106052 50380 106054
rect 50436 106052 50460 106054
rect 50516 106052 50540 106054
rect 50300 106032 50596 106052
rect 50300 105020 50596 105040
rect 50356 105018 50380 105020
rect 50436 105018 50460 105020
rect 50516 105018 50540 105020
rect 50378 104966 50380 105018
rect 50442 104966 50454 105018
rect 50516 104966 50518 105018
rect 50356 104964 50380 104966
rect 50436 104964 50460 104966
rect 50516 104964 50540 104966
rect 50300 104944 50596 104964
rect 50300 103932 50596 103952
rect 50356 103930 50380 103932
rect 50436 103930 50460 103932
rect 50516 103930 50540 103932
rect 50378 103878 50380 103930
rect 50442 103878 50454 103930
rect 50516 103878 50518 103930
rect 50356 103876 50380 103878
rect 50436 103876 50460 103878
rect 50516 103876 50540 103878
rect 50300 103856 50596 103876
rect 50300 102844 50596 102864
rect 50356 102842 50380 102844
rect 50436 102842 50460 102844
rect 50516 102842 50540 102844
rect 50378 102790 50380 102842
rect 50442 102790 50454 102842
rect 50516 102790 50518 102842
rect 50356 102788 50380 102790
rect 50436 102788 50460 102790
rect 50516 102788 50540 102790
rect 50300 102768 50596 102788
rect 50300 101756 50596 101776
rect 50356 101754 50380 101756
rect 50436 101754 50460 101756
rect 50516 101754 50540 101756
rect 50378 101702 50380 101754
rect 50442 101702 50454 101754
rect 50516 101702 50518 101754
rect 50356 101700 50380 101702
rect 50436 101700 50460 101702
rect 50516 101700 50540 101702
rect 50300 101680 50596 101700
rect 50300 100668 50596 100688
rect 50356 100666 50380 100668
rect 50436 100666 50460 100668
rect 50516 100666 50540 100668
rect 50378 100614 50380 100666
rect 50442 100614 50454 100666
rect 50516 100614 50518 100666
rect 50356 100612 50380 100614
rect 50436 100612 50460 100614
rect 50516 100612 50540 100614
rect 50300 100592 50596 100612
rect 50300 99580 50596 99600
rect 50356 99578 50380 99580
rect 50436 99578 50460 99580
rect 50516 99578 50540 99580
rect 50378 99526 50380 99578
rect 50442 99526 50454 99578
rect 50516 99526 50518 99578
rect 50356 99524 50380 99526
rect 50436 99524 50460 99526
rect 50516 99524 50540 99526
rect 50300 99504 50596 99524
rect 50300 98492 50596 98512
rect 50356 98490 50380 98492
rect 50436 98490 50460 98492
rect 50516 98490 50540 98492
rect 50378 98438 50380 98490
rect 50442 98438 50454 98490
rect 50516 98438 50518 98490
rect 50356 98436 50380 98438
rect 50436 98436 50460 98438
rect 50516 98436 50540 98438
rect 50300 98416 50596 98436
rect 50300 97404 50596 97424
rect 50356 97402 50380 97404
rect 50436 97402 50460 97404
rect 50516 97402 50540 97404
rect 50378 97350 50380 97402
rect 50442 97350 50454 97402
rect 50516 97350 50518 97402
rect 50356 97348 50380 97350
rect 50436 97348 50460 97350
rect 50516 97348 50540 97350
rect 50300 97328 50596 97348
rect 50300 96316 50596 96336
rect 50356 96314 50380 96316
rect 50436 96314 50460 96316
rect 50516 96314 50540 96316
rect 50378 96262 50380 96314
rect 50442 96262 50454 96314
rect 50516 96262 50518 96314
rect 50356 96260 50380 96262
rect 50436 96260 50460 96262
rect 50516 96260 50540 96262
rect 50300 96240 50596 96260
rect 50300 95228 50596 95248
rect 50356 95226 50380 95228
rect 50436 95226 50460 95228
rect 50516 95226 50540 95228
rect 50378 95174 50380 95226
rect 50442 95174 50454 95226
rect 50516 95174 50518 95226
rect 50356 95172 50380 95174
rect 50436 95172 50460 95174
rect 50516 95172 50540 95174
rect 50300 95152 50596 95172
rect 50300 94140 50596 94160
rect 50356 94138 50380 94140
rect 50436 94138 50460 94140
rect 50516 94138 50540 94140
rect 50378 94086 50380 94138
rect 50442 94086 50454 94138
rect 50516 94086 50518 94138
rect 50356 94084 50380 94086
rect 50436 94084 50460 94086
rect 50516 94084 50540 94086
rect 50300 94064 50596 94084
rect 50300 93052 50596 93072
rect 50356 93050 50380 93052
rect 50436 93050 50460 93052
rect 50516 93050 50540 93052
rect 50378 92998 50380 93050
rect 50442 92998 50454 93050
rect 50516 92998 50518 93050
rect 50356 92996 50380 92998
rect 50436 92996 50460 92998
rect 50516 92996 50540 92998
rect 50300 92976 50596 92996
rect 50300 91964 50596 91984
rect 50356 91962 50380 91964
rect 50436 91962 50460 91964
rect 50516 91962 50540 91964
rect 50378 91910 50380 91962
rect 50442 91910 50454 91962
rect 50516 91910 50518 91962
rect 50356 91908 50380 91910
rect 50436 91908 50460 91910
rect 50516 91908 50540 91910
rect 50300 91888 50596 91908
rect 50300 90876 50596 90896
rect 50356 90874 50380 90876
rect 50436 90874 50460 90876
rect 50516 90874 50540 90876
rect 50378 90822 50380 90874
rect 50442 90822 50454 90874
rect 50516 90822 50518 90874
rect 50356 90820 50380 90822
rect 50436 90820 50460 90822
rect 50516 90820 50540 90822
rect 50300 90800 50596 90820
rect 50300 89788 50596 89808
rect 50356 89786 50380 89788
rect 50436 89786 50460 89788
rect 50516 89786 50540 89788
rect 50378 89734 50380 89786
rect 50442 89734 50454 89786
rect 50516 89734 50518 89786
rect 50356 89732 50380 89734
rect 50436 89732 50460 89734
rect 50516 89732 50540 89734
rect 50300 89712 50596 89732
rect 50300 88700 50596 88720
rect 50356 88698 50380 88700
rect 50436 88698 50460 88700
rect 50516 88698 50540 88700
rect 50378 88646 50380 88698
rect 50442 88646 50454 88698
rect 50516 88646 50518 88698
rect 50356 88644 50380 88646
rect 50436 88644 50460 88646
rect 50516 88644 50540 88646
rect 50300 88624 50596 88644
rect 50300 87612 50596 87632
rect 50356 87610 50380 87612
rect 50436 87610 50460 87612
rect 50516 87610 50540 87612
rect 50378 87558 50380 87610
rect 50442 87558 50454 87610
rect 50516 87558 50518 87610
rect 50356 87556 50380 87558
rect 50436 87556 50460 87558
rect 50516 87556 50540 87558
rect 50300 87536 50596 87556
rect 50300 86524 50596 86544
rect 50356 86522 50380 86524
rect 50436 86522 50460 86524
rect 50516 86522 50540 86524
rect 50378 86470 50380 86522
rect 50442 86470 50454 86522
rect 50516 86470 50518 86522
rect 50356 86468 50380 86470
rect 50436 86468 50460 86470
rect 50516 86468 50540 86470
rect 50300 86448 50596 86468
rect 50300 85436 50596 85456
rect 50356 85434 50380 85436
rect 50436 85434 50460 85436
rect 50516 85434 50540 85436
rect 50378 85382 50380 85434
rect 50442 85382 50454 85434
rect 50516 85382 50518 85434
rect 50356 85380 50380 85382
rect 50436 85380 50460 85382
rect 50516 85380 50540 85382
rect 50300 85360 50596 85380
rect 50300 84348 50596 84368
rect 50356 84346 50380 84348
rect 50436 84346 50460 84348
rect 50516 84346 50540 84348
rect 50378 84294 50380 84346
rect 50442 84294 50454 84346
rect 50516 84294 50518 84346
rect 50356 84292 50380 84294
rect 50436 84292 50460 84294
rect 50516 84292 50540 84294
rect 50300 84272 50596 84292
rect 50300 83260 50596 83280
rect 50356 83258 50380 83260
rect 50436 83258 50460 83260
rect 50516 83258 50540 83260
rect 50378 83206 50380 83258
rect 50442 83206 50454 83258
rect 50516 83206 50518 83258
rect 50356 83204 50380 83206
rect 50436 83204 50460 83206
rect 50516 83204 50540 83206
rect 50300 83184 50596 83204
rect 50300 82172 50596 82192
rect 50356 82170 50380 82172
rect 50436 82170 50460 82172
rect 50516 82170 50540 82172
rect 50378 82118 50380 82170
rect 50442 82118 50454 82170
rect 50516 82118 50518 82170
rect 50356 82116 50380 82118
rect 50436 82116 50460 82118
rect 50516 82116 50540 82118
rect 50300 82096 50596 82116
rect 50300 81084 50596 81104
rect 50356 81082 50380 81084
rect 50436 81082 50460 81084
rect 50516 81082 50540 81084
rect 50378 81030 50380 81082
rect 50442 81030 50454 81082
rect 50516 81030 50518 81082
rect 50356 81028 50380 81030
rect 50436 81028 50460 81030
rect 50516 81028 50540 81030
rect 50300 81008 50596 81028
rect 50300 79996 50596 80016
rect 50356 79994 50380 79996
rect 50436 79994 50460 79996
rect 50516 79994 50540 79996
rect 50378 79942 50380 79994
rect 50442 79942 50454 79994
rect 50516 79942 50518 79994
rect 50356 79940 50380 79942
rect 50436 79940 50460 79942
rect 50516 79940 50540 79942
rect 50300 79920 50596 79940
rect 50300 78908 50596 78928
rect 50356 78906 50380 78908
rect 50436 78906 50460 78908
rect 50516 78906 50540 78908
rect 50378 78854 50380 78906
rect 50442 78854 50454 78906
rect 50516 78854 50518 78906
rect 50356 78852 50380 78854
rect 50436 78852 50460 78854
rect 50516 78852 50540 78854
rect 50300 78832 50596 78852
rect 50300 77820 50596 77840
rect 50356 77818 50380 77820
rect 50436 77818 50460 77820
rect 50516 77818 50540 77820
rect 50378 77766 50380 77818
rect 50442 77766 50454 77818
rect 50516 77766 50518 77818
rect 50356 77764 50380 77766
rect 50436 77764 50460 77766
rect 50516 77764 50540 77766
rect 50300 77744 50596 77764
rect 50300 76732 50596 76752
rect 50356 76730 50380 76732
rect 50436 76730 50460 76732
rect 50516 76730 50540 76732
rect 50378 76678 50380 76730
rect 50442 76678 50454 76730
rect 50516 76678 50518 76730
rect 50356 76676 50380 76678
rect 50436 76676 50460 76678
rect 50516 76676 50540 76678
rect 50300 76656 50596 76676
rect 50300 75644 50596 75664
rect 50356 75642 50380 75644
rect 50436 75642 50460 75644
rect 50516 75642 50540 75644
rect 50378 75590 50380 75642
rect 50442 75590 50454 75642
rect 50516 75590 50518 75642
rect 50356 75588 50380 75590
rect 50436 75588 50460 75590
rect 50516 75588 50540 75590
rect 50300 75568 50596 75588
rect 50300 74556 50596 74576
rect 50356 74554 50380 74556
rect 50436 74554 50460 74556
rect 50516 74554 50540 74556
rect 50378 74502 50380 74554
rect 50442 74502 50454 74554
rect 50516 74502 50518 74554
rect 50356 74500 50380 74502
rect 50436 74500 50460 74502
rect 50516 74500 50540 74502
rect 50300 74480 50596 74500
rect 50300 73468 50596 73488
rect 50356 73466 50380 73468
rect 50436 73466 50460 73468
rect 50516 73466 50540 73468
rect 50378 73414 50380 73466
rect 50442 73414 50454 73466
rect 50516 73414 50518 73466
rect 50356 73412 50380 73414
rect 50436 73412 50460 73414
rect 50516 73412 50540 73414
rect 50300 73392 50596 73412
rect 50300 72380 50596 72400
rect 50356 72378 50380 72380
rect 50436 72378 50460 72380
rect 50516 72378 50540 72380
rect 50378 72326 50380 72378
rect 50442 72326 50454 72378
rect 50516 72326 50518 72378
rect 50356 72324 50380 72326
rect 50436 72324 50460 72326
rect 50516 72324 50540 72326
rect 50300 72304 50596 72324
rect 50300 71292 50596 71312
rect 50356 71290 50380 71292
rect 50436 71290 50460 71292
rect 50516 71290 50540 71292
rect 50378 71238 50380 71290
rect 50442 71238 50454 71290
rect 50516 71238 50518 71290
rect 50356 71236 50380 71238
rect 50436 71236 50460 71238
rect 50516 71236 50540 71238
rect 50300 71216 50596 71236
rect 50300 70204 50596 70224
rect 50356 70202 50380 70204
rect 50436 70202 50460 70204
rect 50516 70202 50540 70204
rect 50378 70150 50380 70202
rect 50442 70150 50454 70202
rect 50516 70150 50518 70202
rect 50356 70148 50380 70150
rect 50436 70148 50460 70150
rect 50516 70148 50540 70150
rect 50300 70128 50596 70148
rect 50300 69116 50596 69136
rect 50356 69114 50380 69116
rect 50436 69114 50460 69116
rect 50516 69114 50540 69116
rect 50378 69062 50380 69114
rect 50442 69062 50454 69114
rect 50516 69062 50518 69114
rect 50356 69060 50380 69062
rect 50436 69060 50460 69062
rect 50516 69060 50540 69062
rect 50300 69040 50596 69060
rect 50300 68028 50596 68048
rect 50356 68026 50380 68028
rect 50436 68026 50460 68028
rect 50516 68026 50540 68028
rect 50378 67974 50380 68026
rect 50442 67974 50454 68026
rect 50516 67974 50518 68026
rect 50356 67972 50380 67974
rect 50436 67972 50460 67974
rect 50516 67972 50540 67974
rect 50300 67952 50596 67972
rect 50300 66940 50596 66960
rect 50356 66938 50380 66940
rect 50436 66938 50460 66940
rect 50516 66938 50540 66940
rect 50378 66886 50380 66938
rect 50442 66886 50454 66938
rect 50516 66886 50518 66938
rect 50356 66884 50380 66886
rect 50436 66884 50460 66886
rect 50516 66884 50540 66886
rect 50300 66864 50596 66884
rect 50300 65852 50596 65872
rect 50356 65850 50380 65852
rect 50436 65850 50460 65852
rect 50516 65850 50540 65852
rect 50378 65798 50380 65850
rect 50442 65798 50454 65850
rect 50516 65798 50518 65850
rect 50356 65796 50380 65798
rect 50436 65796 50460 65798
rect 50516 65796 50540 65798
rect 50300 65776 50596 65796
rect 50300 64764 50596 64784
rect 50356 64762 50380 64764
rect 50436 64762 50460 64764
rect 50516 64762 50540 64764
rect 50378 64710 50380 64762
rect 50442 64710 50454 64762
rect 50516 64710 50518 64762
rect 50356 64708 50380 64710
rect 50436 64708 50460 64710
rect 50516 64708 50540 64710
rect 50300 64688 50596 64708
rect 50300 63676 50596 63696
rect 50356 63674 50380 63676
rect 50436 63674 50460 63676
rect 50516 63674 50540 63676
rect 50378 63622 50380 63674
rect 50442 63622 50454 63674
rect 50516 63622 50518 63674
rect 50356 63620 50380 63622
rect 50436 63620 50460 63622
rect 50516 63620 50540 63622
rect 50300 63600 50596 63620
rect 50300 62588 50596 62608
rect 50356 62586 50380 62588
rect 50436 62586 50460 62588
rect 50516 62586 50540 62588
rect 50378 62534 50380 62586
rect 50442 62534 50454 62586
rect 50516 62534 50518 62586
rect 50356 62532 50380 62534
rect 50436 62532 50460 62534
rect 50516 62532 50540 62534
rect 50300 62512 50596 62532
rect 50300 61500 50596 61520
rect 50356 61498 50380 61500
rect 50436 61498 50460 61500
rect 50516 61498 50540 61500
rect 50378 61446 50380 61498
rect 50442 61446 50454 61498
rect 50516 61446 50518 61498
rect 50356 61444 50380 61446
rect 50436 61444 50460 61446
rect 50516 61444 50540 61446
rect 50300 61424 50596 61444
rect 50300 60412 50596 60432
rect 50356 60410 50380 60412
rect 50436 60410 50460 60412
rect 50516 60410 50540 60412
rect 50378 60358 50380 60410
rect 50442 60358 50454 60410
rect 50516 60358 50518 60410
rect 50356 60356 50380 60358
rect 50436 60356 50460 60358
rect 50516 60356 50540 60358
rect 50300 60336 50596 60356
rect 50300 59324 50596 59344
rect 50356 59322 50380 59324
rect 50436 59322 50460 59324
rect 50516 59322 50540 59324
rect 50378 59270 50380 59322
rect 50442 59270 50454 59322
rect 50516 59270 50518 59322
rect 50356 59268 50380 59270
rect 50436 59268 50460 59270
rect 50516 59268 50540 59270
rect 50300 59248 50596 59268
rect 50300 58236 50596 58256
rect 50356 58234 50380 58236
rect 50436 58234 50460 58236
rect 50516 58234 50540 58236
rect 50378 58182 50380 58234
rect 50442 58182 50454 58234
rect 50516 58182 50518 58234
rect 50356 58180 50380 58182
rect 50436 58180 50460 58182
rect 50516 58180 50540 58182
rect 50300 58160 50596 58180
rect 50300 57148 50596 57168
rect 50356 57146 50380 57148
rect 50436 57146 50460 57148
rect 50516 57146 50540 57148
rect 50378 57094 50380 57146
rect 50442 57094 50454 57146
rect 50516 57094 50518 57146
rect 50356 57092 50380 57094
rect 50436 57092 50460 57094
rect 50516 57092 50540 57094
rect 50300 57072 50596 57092
rect 50300 56060 50596 56080
rect 50356 56058 50380 56060
rect 50436 56058 50460 56060
rect 50516 56058 50540 56060
rect 50378 56006 50380 56058
rect 50442 56006 50454 56058
rect 50516 56006 50518 56058
rect 50356 56004 50380 56006
rect 50436 56004 50460 56006
rect 50516 56004 50540 56006
rect 50300 55984 50596 56004
rect 50300 54972 50596 54992
rect 50356 54970 50380 54972
rect 50436 54970 50460 54972
rect 50516 54970 50540 54972
rect 50378 54918 50380 54970
rect 50442 54918 50454 54970
rect 50516 54918 50518 54970
rect 50356 54916 50380 54918
rect 50436 54916 50460 54918
rect 50516 54916 50540 54918
rect 50300 54896 50596 54916
rect 50300 53884 50596 53904
rect 50356 53882 50380 53884
rect 50436 53882 50460 53884
rect 50516 53882 50540 53884
rect 50378 53830 50380 53882
rect 50442 53830 50454 53882
rect 50516 53830 50518 53882
rect 50356 53828 50380 53830
rect 50436 53828 50460 53830
rect 50516 53828 50540 53830
rect 50300 53808 50596 53828
rect 50300 52796 50596 52816
rect 50356 52794 50380 52796
rect 50436 52794 50460 52796
rect 50516 52794 50540 52796
rect 50378 52742 50380 52794
rect 50442 52742 50454 52794
rect 50516 52742 50518 52794
rect 50356 52740 50380 52742
rect 50436 52740 50460 52742
rect 50516 52740 50540 52742
rect 50300 52720 50596 52740
rect 50300 51708 50596 51728
rect 50356 51706 50380 51708
rect 50436 51706 50460 51708
rect 50516 51706 50540 51708
rect 50378 51654 50380 51706
rect 50442 51654 50454 51706
rect 50516 51654 50518 51706
rect 50356 51652 50380 51654
rect 50436 51652 50460 51654
rect 50516 51652 50540 51654
rect 50300 51632 50596 51652
rect 50300 50620 50596 50640
rect 50356 50618 50380 50620
rect 50436 50618 50460 50620
rect 50516 50618 50540 50620
rect 50378 50566 50380 50618
rect 50442 50566 50454 50618
rect 50516 50566 50518 50618
rect 50356 50564 50380 50566
rect 50436 50564 50460 50566
rect 50516 50564 50540 50566
rect 50300 50544 50596 50564
rect 50300 49532 50596 49552
rect 50356 49530 50380 49532
rect 50436 49530 50460 49532
rect 50516 49530 50540 49532
rect 50378 49478 50380 49530
rect 50442 49478 50454 49530
rect 50516 49478 50518 49530
rect 50356 49476 50380 49478
rect 50436 49476 50460 49478
rect 50516 49476 50540 49478
rect 50300 49456 50596 49476
rect 50300 48444 50596 48464
rect 50356 48442 50380 48444
rect 50436 48442 50460 48444
rect 50516 48442 50540 48444
rect 50378 48390 50380 48442
rect 50442 48390 50454 48442
rect 50516 48390 50518 48442
rect 50356 48388 50380 48390
rect 50436 48388 50460 48390
rect 50516 48388 50540 48390
rect 50300 48368 50596 48388
rect 50300 47356 50596 47376
rect 50356 47354 50380 47356
rect 50436 47354 50460 47356
rect 50516 47354 50540 47356
rect 50378 47302 50380 47354
rect 50442 47302 50454 47354
rect 50516 47302 50518 47354
rect 50356 47300 50380 47302
rect 50436 47300 50460 47302
rect 50516 47300 50540 47302
rect 50300 47280 50596 47300
rect 50300 46268 50596 46288
rect 50356 46266 50380 46268
rect 50436 46266 50460 46268
rect 50516 46266 50540 46268
rect 50378 46214 50380 46266
rect 50442 46214 50454 46266
rect 50516 46214 50518 46266
rect 50356 46212 50380 46214
rect 50436 46212 50460 46214
rect 50516 46212 50540 46214
rect 50300 46192 50596 46212
rect 50300 45180 50596 45200
rect 50356 45178 50380 45180
rect 50436 45178 50460 45180
rect 50516 45178 50540 45180
rect 50378 45126 50380 45178
rect 50442 45126 50454 45178
rect 50516 45126 50518 45178
rect 50356 45124 50380 45126
rect 50436 45124 50460 45126
rect 50516 45124 50540 45126
rect 50300 45104 50596 45124
rect 50300 44092 50596 44112
rect 50356 44090 50380 44092
rect 50436 44090 50460 44092
rect 50516 44090 50540 44092
rect 50378 44038 50380 44090
rect 50442 44038 50454 44090
rect 50516 44038 50518 44090
rect 50356 44036 50380 44038
rect 50436 44036 50460 44038
rect 50516 44036 50540 44038
rect 50300 44016 50596 44036
rect 50300 43004 50596 43024
rect 50356 43002 50380 43004
rect 50436 43002 50460 43004
rect 50516 43002 50540 43004
rect 50378 42950 50380 43002
rect 50442 42950 50454 43002
rect 50516 42950 50518 43002
rect 50356 42948 50380 42950
rect 50436 42948 50460 42950
rect 50516 42948 50540 42950
rect 50300 42928 50596 42948
rect 50300 41916 50596 41936
rect 50356 41914 50380 41916
rect 50436 41914 50460 41916
rect 50516 41914 50540 41916
rect 50378 41862 50380 41914
rect 50442 41862 50454 41914
rect 50516 41862 50518 41914
rect 50356 41860 50380 41862
rect 50436 41860 50460 41862
rect 50516 41860 50540 41862
rect 50300 41840 50596 41860
rect 50300 40828 50596 40848
rect 50356 40826 50380 40828
rect 50436 40826 50460 40828
rect 50516 40826 50540 40828
rect 50378 40774 50380 40826
rect 50442 40774 50454 40826
rect 50516 40774 50518 40826
rect 50356 40772 50380 40774
rect 50436 40772 50460 40774
rect 50516 40772 50540 40774
rect 50300 40752 50596 40772
rect 50300 39740 50596 39760
rect 50356 39738 50380 39740
rect 50436 39738 50460 39740
rect 50516 39738 50540 39740
rect 50378 39686 50380 39738
rect 50442 39686 50454 39738
rect 50516 39686 50518 39738
rect 50356 39684 50380 39686
rect 50436 39684 50460 39686
rect 50516 39684 50540 39686
rect 50300 39664 50596 39684
rect 50300 38652 50596 38672
rect 50356 38650 50380 38652
rect 50436 38650 50460 38652
rect 50516 38650 50540 38652
rect 50378 38598 50380 38650
rect 50442 38598 50454 38650
rect 50516 38598 50518 38650
rect 50356 38596 50380 38598
rect 50436 38596 50460 38598
rect 50516 38596 50540 38598
rect 50300 38576 50596 38596
rect 50300 37564 50596 37584
rect 50356 37562 50380 37564
rect 50436 37562 50460 37564
rect 50516 37562 50540 37564
rect 50378 37510 50380 37562
rect 50442 37510 50454 37562
rect 50516 37510 50518 37562
rect 50356 37508 50380 37510
rect 50436 37508 50460 37510
rect 50516 37508 50540 37510
rect 50300 37488 50596 37508
rect 50300 36476 50596 36496
rect 50356 36474 50380 36476
rect 50436 36474 50460 36476
rect 50516 36474 50540 36476
rect 50378 36422 50380 36474
rect 50442 36422 50454 36474
rect 50516 36422 50518 36474
rect 50356 36420 50380 36422
rect 50436 36420 50460 36422
rect 50516 36420 50540 36422
rect 50300 36400 50596 36420
rect 50300 35388 50596 35408
rect 50356 35386 50380 35388
rect 50436 35386 50460 35388
rect 50516 35386 50540 35388
rect 50378 35334 50380 35386
rect 50442 35334 50454 35386
rect 50516 35334 50518 35386
rect 50356 35332 50380 35334
rect 50436 35332 50460 35334
rect 50516 35332 50540 35334
rect 50300 35312 50596 35332
rect 50300 34300 50596 34320
rect 50356 34298 50380 34300
rect 50436 34298 50460 34300
rect 50516 34298 50540 34300
rect 50378 34246 50380 34298
rect 50442 34246 50454 34298
rect 50516 34246 50518 34298
rect 50356 34244 50380 34246
rect 50436 34244 50460 34246
rect 50516 34244 50540 34246
rect 50300 34224 50596 34244
rect 50300 33212 50596 33232
rect 50356 33210 50380 33212
rect 50436 33210 50460 33212
rect 50516 33210 50540 33212
rect 50378 33158 50380 33210
rect 50442 33158 50454 33210
rect 50516 33158 50518 33210
rect 50356 33156 50380 33158
rect 50436 33156 50460 33158
rect 50516 33156 50540 33158
rect 50300 33136 50596 33156
rect 50300 32124 50596 32144
rect 50356 32122 50380 32124
rect 50436 32122 50460 32124
rect 50516 32122 50540 32124
rect 50378 32070 50380 32122
rect 50442 32070 50454 32122
rect 50516 32070 50518 32122
rect 50356 32068 50380 32070
rect 50436 32068 50460 32070
rect 50516 32068 50540 32070
rect 50300 32048 50596 32068
rect 50300 31036 50596 31056
rect 50356 31034 50380 31036
rect 50436 31034 50460 31036
rect 50516 31034 50540 31036
rect 50378 30982 50380 31034
rect 50442 30982 50454 31034
rect 50516 30982 50518 31034
rect 50356 30980 50380 30982
rect 50436 30980 50460 30982
rect 50516 30980 50540 30982
rect 50300 30960 50596 30980
rect 50300 29948 50596 29968
rect 50356 29946 50380 29948
rect 50436 29946 50460 29948
rect 50516 29946 50540 29948
rect 50378 29894 50380 29946
rect 50442 29894 50454 29946
rect 50516 29894 50518 29946
rect 50356 29892 50380 29894
rect 50436 29892 50460 29894
rect 50516 29892 50540 29894
rect 50300 29872 50596 29892
rect 50300 28860 50596 28880
rect 50356 28858 50380 28860
rect 50436 28858 50460 28860
rect 50516 28858 50540 28860
rect 50378 28806 50380 28858
rect 50442 28806 50454 28858
rect 50516 28806 50518 28858
rect 50356 28804 50380 28806
rect 50436 28804 50460 28806
rect 50516 28804 50540 28806
rect 50300 28784 50596 28804
rect 50300 27772 50596 27792
rect 50356 27770 50380 27772
rect 50436 27770 50460 27772
rect 50516 27770 50540 27772
rect 50378 27718 50380 27770
rect 50442 27718 50454 27770
rect 50516 27718 50518 27770
rect 50356 27716 50380 27718
rect 50436 27716 50460 27718
rect 50516 27716 50540 27718
rect 50300 27696 50596 27716
rect 50300 26684 50596 26704
rect 50356 26682 50380 26684
rect 50436 26682 50460 26684
rect 50516 26682 50540 26684
rect 50378 26630 50380 26682
rect 50442 26630 50454 26682
rect 50516 26630 50518 26682
rect 50356 26628 50380 26630
rect 50436 26628 50460 26630
rect 50516 26628 50540 26630
rect 50300 26608 50596 26628
rect 50300 25596 50596 25616
rect 50356 25594 50380 25596
rect 50436 25594 50460 25596
rect 50516 25594 50540 25596
rect 50378 25542 50380 25594
rect 50442 25542 50454 25594
rect 50516 25542 50518 25594
rect 50356 25540 50380 25542
rect 50436 25540 50460 25542
rect 50516 25540 50540 25542
rect 50300 25520 50596 25540
rect 50300 24508 50596 24528
rect 50356 24506 50380 24508
rect 50436 24506 50460 24508
rect 50516 24506 50540 24508
rect 50378 24454 50380 24506
rect 50442 24454 50454 24506
rect 50516 24454 50518 24506
rect 50356 24452 50380 24454
rect 50436 24452 50460 24454
rect 50516 24452 50540 24454
rect 50300 24432 50596 24452
rect 50300 23420 50596 23440
rect 50356 23418 50380 23420
rect 50436 23418 50460 23420
rect 50516 23418 50540 23420
rect 50378 23366 50380 23418
rect 50442 23366 50454 23418
rect 50516 23366 50518 23418
rect 50356 23364 50380 23366
rect 50436 23364 50460 23366
rect 50516 23364 50540 23366
rect 50300 23344 50596 23364
rect 50300 22332 50596 22352
rect 50356 22330 50380 22332
rect 50436 22330 50460 22332
rect 50516 22330 50540 22332
rect 50378 22278 50380 22330
rect 50442 22278 50454 22330
rect 50516 22278 50518 22330
rect 50356 22276 50380 22278
rect 50436 22276 50460 22278
rect 50516 22276 50540 22278
rect 50300 22256 50596 22276
rect 47044 22066 47164 22094
rect 37740 19304 37792 19310
rect 37740 19246 37792 19252
rect 41696 19304 41748 19310
rect 41696 19246 41748 19252
rect 37464 19168 37516 19174
rect 37464 19110 37516 19116
rect 37476 18222 37504 19110
rect 37464 18216 37516 18222
rect 37464 18158 37516 18164
rect 37476 17746 37504 18158
rect 37752 17746 37780 19246
rect 42800 19168 42852 19174
rect 42800 19110 42852 19116
rect 43444 19168 43496 19174
rect 43444 19110 43496 19116
rect 42812 18834 42840 19110
rect 42800 18828 42852 18834
rect 42800 18770 42852 18776
rect 42892 18624 42944 18630
rect 42892 18566 42944 18572
rect 41420 18216 41472 18222
rect 41420 18158 41472 18164
rect 41144 18148 41196 18154
rect 41144 18090 41196 18096
rect 37464 17740 37516 17746
rect 37464 17682 37516 17688
rect 37740 17740 37792 17746
rect 37740 17682 37792 17688
rect 38752 17740 38804 17746
rect 38752 17682 38804 17688
rect 35900 17128 35952 17134
rect 35900 17070 35952 17076
rect 35348 14884 35400 14890
rect 35348 14826 35400 14832
rect 34940 14172 35236 14192
rect 34996 14170 35020 14172
rect 35076 14170 35100 14172
rect 35156 14170 35180 14172
rect 35018 14118 35020 14170
rect 35082 14118 35094 14170
rect 35156 14118 35158 14170
rect 34996 14116 35020 14118
rect 35076 14116 35100 14118
rect 35156 14116 35180 14118
rect 34940 14096 35236 14116
rect 35256 14000 35308 14006
rect 35256 13942 35308 13948
rect 34940 13084 35236 13104
rect 34996 13082 35020 13084
rect 35076 13082 35100 13084
rect 35156 13082 35180 13084
rect 35018 13030 35020 13082
rect 35082 13030 35094 13082
rect 35156 13030 35158 13082
rect 34996 13028 35020 13030
rect 35076 13028 35100 13030
rect 35156 13028 35180 13030
rect 34940 13008 35236 13028
rect 34796 12436 34848 12442
rect 34796 12378 34848 12384
rect 34940 11996 35236 12016
rect 34996 11994 35020 11996
rect 35076 11994 35100 11996
rect 35156 11994 35180 11996
rect 35018 11942 35020 11994
rect 35082 11942 35094 11994
rect 35156 11942 35158 11994
rect 34996 11940 35020 11942
rect 35076 11940 35100 11942
rect 35156 11940 35180 11942
rect 34940 11920 35236 11940
rect 34940 10908 35236 10928
rect 34996 10906 35020 10908
rect 35076 10906 35100 10908
rect 35156 10906 35180 10908
rect 35018 10854 35020 10906
rect 35082 10854 35094 10906
rect 35156 10854 35158 10906
rect 34996 10852 35020 10854
rect 35076 10852 35100 10854
rect 35156 10852 35180 10854
rect 34940 10832 35236 10852
rect 34716 10118 34836 10146
rect 34704 10056 34756 10062
rect 34704 9998 34756 10004
rect 34428 9988 34480 9994
rect 34428 9930 34480 9936
rect 33876 9036 33928 9042
rect 33876 8978 33928 8984
rect 33888 8430 33916 8978
rect 33876 8424 33928 8430
rect 33876 8366 33928 8372
rect 33784 8084 33836 8090
rect 33784 8026 33836 8032
rect 33888 7886 33916 8366
rect 33968 8084 34020 8090
rect 33968 8026 34020 8032
rect 33876 7880 33928 7886
rect 33876 7822 33928 7828
rect 33784 7812 33836 7818
rect 33784 7754 33836 7760
rect 33796 7410 33824 7754
rect 33784 7404 33836 7410
rect 33784 7346 33836 7352
rect 33888 7342 33916 7822
rect 33980 7721 34008 8026
rect 34336 8016 34388 8022
rect 34336 7958 34388 7964
rect 33966 7712 34022 7721
rect 33966 7647 34022 7656
rect 33876 7336 33928 7342
rect 33876 7278 33928 7284
rect 34060 7336 34112 7342
rect 34060 7278 34112 7284
rect 34242 7304 34298 7313
rect 33876 7200 33928 7206
rect 33876 7142 33928 7148
rect 33784 6860 33836 6866
rect 33784 6802 33836 6808
rect 33796 6186 33824 6802
rect 33784 6180 33836 6186
rect 33784 6122 33836 6128
rect 33796 6089 33824 6122
rect 33782 6080 33838 6089
rect 33782 6015 33838 6024
rect 33692 5908 33744 5914
rect 33692 5850 33744 5856
rect 33692 5568 33744 5574
rect 33612 5528 33692 5556
rect 33692 5510 33744 5516
rect 33704 4554 33732 5510
rect 33796 4622 33824 6015
rect 33888 5778 33916 7142
rect 34072 6866 34100 7278
rect 34242 7239 34298 7248
rect 34256 7206 34284 7239
rect 34152 7200 34204 7206
rect 34150 7168 34152 7177
rect 34244 7200 34296 7206
rect 34204 7168 34206 7177
rect 34244 7142 34296 7148
rect 34150 7103 34206 7112
rect 34060 6860 34112 6866
rect 34060 6802 34112 6808
rect 33876 5772 33928 5778
rect 33876 5714 33928 5720
rect 34060 5636 34112 5642
rect 34060 5578 34112 5584
rect 33784 4616 33836 4622
rect 33784 4558 33836 4564
rect 33692 4548 33744 4554
rect 33692 4490 33744 4496
rect 34072 4214 34100 5578
rect 34060 4208 34112 4214
rect 34060 4150 34112 4156
rect 34164 4010 34192 7103
rect 34348 5370 34376 7958
rect 34440 6458 34468 9930
rect 34716 7018 34744 9998
rect 34808 7460 34836 10118
rect 34940 9820 35236 9840
rect 34996 9818 35020 9820
rect 35076 9818 35100 9820
rect 35156 9818 35180 9820
rect 35018 9766 35020 9818
rect 35082 9766 35094 9818
rect 35156 9766 35158 9818
rect 34996 9764 35020 9766
rect 35076 9764 35100 9766
rect 35156 9764 35180 9766
rect 34940 9744 35236 9764
rect 34940 8732 35236 8752
rect 34996 8730 35020 8732
rect 35076 8730 35100 8732
rect 35156 8730 35180 8732
rect 35018 8678 35020 8730
rect 35082 8678 35094 8730
rect 35156 8678 35158 8730
rect 34996 8676 35020 8678
rect 35076 8676 35100 8678
rect 35156 8676 35180 8678
rect 34940 8656 35236 8676
rect 34940 7644 35236 7664
rect 34996 7642 35020 7644
rect 35076 7642 35100 7644
rect 35156 7642 35180 7644
rect 35018 7590 35020 7642
rect 35082 7590 35094 7642
rect 35156 7590 35158 7642
rect 34996 7588 35020 7590
rect 35076 7588 35100 7590
rect 35156 7588 35180 7590
rect 34940 7568 35236 7588
rect 34808 7432 35020 7460
rect 34796 7268 34848 7274
rect 34796 7210 34848 7216
rect 34808 7177 34836 7210
rect 34794 7168 34850 7177
rect 34992 7154 35020 7432
rect 35268 7342 35296 13942
rect 35360 13734 35388 14826
rect 35912 13802 35940 17070
rect 36360 16992 36412 16998
rect 36360 16934 36412 16940
rect 36084 15972 36136 15978
rect 36084 15914 36136 15920
rect 35900 13796 35952 13802
rect 35900 13738 35952 13744
rect 35348 13728 35400 13734
rect 35348 13670 35400 13676
rect 35912 13190 35940 13738
rect 35900 13184 35952 13190
rect 35900 13126 35952 13132
rect 35440 12368 35492 12374
rect 35440 12310 35492 12316
rect 35256 7336 35308 7342
rect 35254 7304 35256 7313
rect 35308 7304 35310 7313
rect 35254 7239 35310 7248
rect 34992 7126 35296 7154
rect 34794 7103 34850 7112
rect 34716 6990 34928 7018
rect 34796 6928 34848 6934
rect 34796 6870 34848 6876
rect 34428 6452 34480 6458
rect 34428 6394 34480 6400
rect 34428 6112 34480 6118
rect 34428 6054 34480 6060
rect 34244 5364 34296 5370
rect 34244 5306 34296 5312
rect 34336 5364 34388 5370
rect 34336 5306 34388 5312
rect 34256 4690 34284 5306
rect 34244 4684 34296 4690
rect 34244 4626 34296 4632
rect 34152 4004 34204 4010
rect 34152 3946 34204 3952
rect 33508 3596 33560 3602
rect 33508 3538 33560 3544
rect 33416 2100 33468 2106
rect 33416 2042 33468 2048
rect 33324 1896 33376 1902
rect 33324 1838 33376 1844
rect 33520 800 33548 3538
rect 34348 3482 34376 5306
rect 34256 3454 34376 3482
rect 34256 3398 34284 3454
rect 34244 3392 34296 3398
rect 34244 3334 34296 3340
rect 34336 3392 34388 3398
rect 34336 3334 34388 3340
rect 34348 2990 34376 3334
rect 34336 2984 34388 2990
rect 34336 2926 34388 2932
rect 34244 2848 34296 2854
rect 34244 2790 34296 2796
rect 33876 2508 33928 2514
rect 33876 2450 33928 2456
rect 33784 2440 33836 2446
rect 33784 2382 33836 2388
rect 33796 2038 33824 2382
rect 33784 2032 33836 2038
rect 33784 1974 33836 1980
rect 33888 800 33916 2450
rect 34256 800 34284 2790
rect 34440 1154 34468 6054
rect 34808 5302 34836 6870
rect 34900 6730 34928 6990
rect 34888 6724 34940 6730
rect 34888 6666 34940 6672
rect 34940 6556 35236 6576
rect 34996 6554 35020 6556
rect 35076 6554 35100 6556
rect 35156 6554 35180 6556
rect 35018 6502 35020 6554
rect 35082 6502 35094 6554
rect 35156 6502 35158 6554
rect 34996 6500 35020 6502
rect 35076 6500 35100 6502
rect 35156 6500 35180 6502
rect 34940 6480 35236 6500
rect 35268 5681 35296 7126
rect 35348 6452 35400 6458
rect 35348 6394 35400 6400
rect 35360 6118 35388 6394
rect 35348 6112 35400 6118
rect 35348 6054 35400 6060
rect 35254 5672 35310 5681
rect 35254 5607 35310 5616
rect 34940 5468 35236 5488
rect 34996 5466 35020 5468
rect 35076 5466 35100 5468
rect 35156 5466 35180 5468
rect 35018 5414 35020 5466
rect 35082 5414 35094 5466
rect 35156 5414 35158 5466
rect 34996 5412 35020 5414
rect 35076 5412 35100 5414
rect 35156 5412 35180 5414
rect 34940 5392 35236 5412
rect 34796 5296 34848 5302
rect 34796 5238 34848 5244
rect 34518 5128 34574 5137
rect 34518 5063 34520 5072
rect 34572 5063 34574 5072
rect 34520 5034 34572 5040
rect 34940 4380 35236 4400
rect 34996 4378 35020 4380
rect 35076 4378 35100 4380
rect 35156 4378 35180 4380
rect 35018 4326 35020 4378
rect 35082 4326 35094 4378
rect 35156 4326 35158 4378
rect 34996 4324 35020 4326
rect 35076 4324 35100 4326
rect 35156 4324 35180 4326
rect 34940 4304 35236 4324
rect 34612 3596 34664 3602
rect 34612 3538 34664 3544
rect 34520 2304 34572 2310
rect 34520 2246 34572 2252
rect 34532 1902 34560 2246
rect 34520 1896 34572 1902
rect 34520 1838 34572 1844
rect 34428 1148 34480 1154
rect 34428 1090 34480 1096
rect 34624 800 34652 3538
rect 35360 3466 35388 6054
rect 35452 5778 35480 12310
rect 35532 12096 35584 12102
rect 35532 12038 35584 12044
rect 35544 6322 35572 12038
rect 35808 10532 35860 10538
rect 35808 10474 35860 10480
rect 35624 8560 35676 8566
rect 35624 8502 35676 8508
rect 35636 7206 35664 8502
rect 35820 7546 35848 10474
rect 35912 9024 35940 13126
rect 36096 12986 36124 15914
rect 36372 13938 36400 16934
rect 36636 14000 36688 14006
rect 36636 13942 36688 13948
rect 36360 13932 36412 13938
rect 36360 13874 36412 13880
rect 36544 13796 36596 13802
rect 36544 13738 36596 13744
rect 36176 13320 36228 13326
rect 36176 13262 36228 13268
rect 36084 12980 36136 12986
rect 36084 12922 36136 12928
rect 36096 12306 36124 12922
rect 36188 12850 36216 13262
rect 36176 12844 36228 12850
rect 36176 12786 36228 12792
rect 36084 12300 36136 12306
rect 36084 12242 36136 12248
rect 36096 9450 36124 12242
rect 36556 12238 36584 13738
rect 36544 12232 36596 12238
rect 36544 12174 36596 12180
rect 36268 9512 36320 9518
rect 36268 9454 36320 9460
rect 36084 9444 36136 9450
rect 36084 9386 36136 9392
rect 35912 8996 36124 9024
rect 35900 8492 35952 8498
rect 35900 8434 35952 8440
rect 35912 8362 35940 8434
rect 35900 8356 35952 8362
rect 35900 8298 35952 8304
rect 35808 7540 35860 7546
rect 35808 7482 35860 7488
rect 35624 7200 35676 7206
rect 35624 7142 35676 7148
rect 35912 7041 35940 8298
rect 35992 7948 36044 7954
rect 35992 7890 36044 7896
rect 35898 7032 35954 7041
rect 35898 6967 35954 6976
rect 36004 6866 36032 7890
rect 36096 6905 36124 8996
rect 36176 7540 36228 7546
rect 36176 7482 36228 7488
rect 36188 7449 36216 7482
rect 36174 7440 36230 7449
rect 36174 7375 36230 7384
rect 36082 6896 36138 6905
rect 35992 6860 36044 6866
rect 36082 6831 36138 6840
rect 35992 6802 36044 6808
rect 35900 6656 35952 6662
rect 35900 6598 35952 6604
rect 35532 6316 35584 6322
rect 35532 6258 35584 6264
rect 35624 6248 35676 6254
rect 35624 6190 35676 6196
rect 35440 5772 35492 5778
rect 35440 5714 35492 5720
rect 35452 5574 35480 5714
rect 35440 5568 35492 5574
rect 35440 5510 35492 5516
rect 35348 3460 35400 3466
rect 35348 3402 35400 3408
rect 35440 3460 35492 3466
rect 35440 3402 35492 3408
rect 34940 3292 35236 3312
rect 34996 3290 35020 3292
rect 35076 3290 35100 3292
rect 35156 3290 35180 3292
rect 35018 3238 35020 3290
rect 35082 3238 35094 3290
rect 35156 3238 35158 3290
rect 34996 3236 35020 3238
rect 35076 3236 35100 3238
rect 35156 3236 35180 3238
rect 34940 3216 35236 3236
rect 35452 2990 35480 3402
rect 35440 2984 35492 2990
rect 35440 2926 35492 2932
rect 35348 2848 35400 2854
rect 35348 2790 35400 2796
rect 35256 2508 35308 2514
rect 35256 2450 35308 2456
rect 34940 2204 35236 2224
rect 34996 2202 35020 2204
rect 35076 2202 35100 2204
rect 35156 2202 35180 2204
rect 35018 2150 35020 2202
rect 35082 2150 35094 2202
rect 35156 2150 35158 2202
rect 34996 2148 35020 2150
rect 35076 2148 35100 2150
rect 35156 2148 35180 2150
rect 34940 2128 35236 2148
rect 35268 1306 35296 2450
rect 34992 1278 35296 1306
rect 34992 800 35020 1278
rect 35360 800 35388 2790
rect 35636 1358 35664 6190
rect 35912 4486 35940 6598
rect 36004 6118 36032 6802
rect 35992 6112 36044 6118
rect 35992 6054 36044 6060
rect 36096 5370 36124 6831
rect 36176 6316 36228 6322
rect 36176 6258 36228 6264
rect 36188 6225 36216 6258
rect 36174 6216 36230 6225
rect 36174 6151 36230 6160
rect 36280 5778 36308 9454
rect 36360 8016 36412 8022
rect 36412 7976 36492 8004
rect 36360 7958 36412 7964
rect 36360 7812 36412 7818
rect 36360 7754 36412 7760
rect 36372 7342 36400 7754
rect 36360 7336 36412 7342
rect 36360 7278 36412 7284
rect 36464 7274 36492 7976
rect 36452 7268 36504 7274
rect 36452 7210 36504 7216
rect 36648 6905 36676 13942
rect 38764 13802 38792 17682
rect 38844 17604 38896 17610
rect 38844 17546 38896 17552
rect 38856 13938 38884 17546
rect 41156 16658 41184 18090
rect 41328 18080 41380 18086
rect 41328 18022 41380 18028
rect 40960 16652 41012 16658
rect 40960 16594 41012 16600
rect 41144 16652 41196 16658
rect 41144 16594 41196 16600
rect 39672 14544 39724 14550
rect 39672 14486 39724 14492
rect 39580 14000 39632 14006
rect 39580 13942 39632 13948
rect 38844 13932 38896 13938
rect 38844 13874 38896 13880
rect 38752 13796 38804 13802
rect 38752 13738 38804 13744
rect 38200 13524 38252 13530
rect 38200 13466 38252 13472
rect 37004 12844 37056 12850
rect 37004 12786 37056 12792
rect 37016 12306 37044 12786
rect 37188 12776 37240 12782
rect 37188 12718 37240 12724
rect 37004 12300 37056 12306
rect 37004 12242 37056 12248
rect 37004 12164 37056 12170
rect 37004 12106 37056 12112
rect 36728 7812 36780 7818
rect 36728 7754 36780 7760
rect 36740 7342 36768 7754
rect 36728 7336 36780 7342
rect 36728 7278 36780 7284
rect 36820 7200 36872 7206
rect 36820 7142 36872 7148
rect 36832 6934 36860 7142
rect 36820 6928 36872 6934
rect 36634 6896 36690 6905
rect 36820 6870 36872 6876
rect 36634 6831 36636 6840
rect 36688 6831 36690 6840
rect 36636 6802 36688 6808
rect 36648 6771 36676 6802
rect 36728 6792 36780 6798
rect 36912 6792 36964 6798
rect 36728 6734 36780 6740
rect 36832 6740 36912 6746
rect 36832 6734 36964 6740
rect 36544 6724 36596 6730
rect 36544 6666 36596 6672
rect 36556 6458 36584 6666
rect 36452 6452 36504 6458
rect 36452 6394 36504 6400
rect 36544 6452 36596 6458
rect 36544 6394 36596 6400
rect 36464 6254 36492 6394
rect 36452 6248 36504 6254
rect 36452 6190 36504 6196
rect 36268 5772 36320 5778
rect 36268 5714 36320 5720
rect 36544 5568 36596 5574
rect 36544 5510 36596 5516
rect 35992 5364 36044 5370
rect 35992 5306 36044 5312
rect 36084 5364 36136 5370
rect 36084 5306 36136 5312
rect 36004 4570 36032 5306
rect 36268 5024 36320 5030
rect 36268 4966 36320 4972
rect 36004 4554 36124 4570
rect 36004 4548 36136 4554
rect 36004 4542 36084 4548
rect 35900 4480 35952 4486
rect 35900 4422 35952 4428
rect 36004 4146 36032 4542
rect 36084 4490 36136 4496
rect 36082 4176 36138 4185
rect 35992 4140 36044 4146
rect 36082 4111 36138 4120
rect 35992 4082 36044 4088
rect 36096 4078 36124 4111
rect 36084 4072 36136 4078
rect 36084 4014 36136 4020
rect 35716 3596 35768 3602
rect 35716 3538 35768 3544
rect 35624 1352 35676 1358
rect 35624 1294 35676 1300
rect 35728 800 35756 3538
rect 36280 2922 36308 4966
rect 36452 3528 36504 3534
rect 36452 3470 36504 3476
rect 36464 3126 36492 3470
rect 36452 3120 36504 3126
rect 36452 3062 36504 3068
rect 36268 2916 36320 2922
rect 36268 2858 36320 2864
rect 36452 2848 36504 2854
rect 36452 2790 36504 2796
rect 36084 2508 36136 2514
rect 36084 2450 36136 2456
rect 36096 800 36124 2450
rect 36464 800 36492 2790
rect 36556 2582 36584 5510
rect 36636 4752 36688 4758
rect 36636 4694 36688 4700
rect 36648 4486 36676 4694
rect 36636 4480 36688 4486
rect 36636 4422 36688 4428
rect 36544 2576 36596 2582
rect 36544 2518 36596 2524
rect 36740 1290 36768 6734
rect 36832 6718 36952 6734
rect 36832 6662 36860 6718
rect 36820 6656 36872 6662
rect 36820 6598 36872 6604
rect 36912 6316 36964 6322
rect 36912 6258 36964 6264
rect 36924 4622 36952 6258
rect 37016 4826 37044 12106
rect 37200 9654 37228 12718
rect 37188 9648 37240 9654
rect 37188 9590 37240 9596
rect 37372 9444 37424 9450
rect 37372 9386 37424 9392
rect 37096 7404 37148 7410
rect 37096 7346 37148 7352
rect 37108 5030 37136 7346
rect 37280 7200 37332 7206
rect 37280 7142 37332 7148
rect 37188 6792 37240 6798
rect 37188 6734 37240 6740
rect 37200 6225 37228 6734
rect 37186 6216 37242 6225
rect 37186 6151 37242 6160
rect 37188 5840 37240 5846
rect 37188 5782 37240 5788
rect 37096 5024 37148 5030
rect 37096 4966 37148 4972
rect 37004 4820 37056 4826
rect 37004 4762 37056 4768
rect 36912 4616 36964 4622
rect 36912 4558 36964 4564
rect 37200 4554 37228 5782
rect 37292 5302 37320 7142
rect 37384 6458 37412 9386
rect 37740 9376 37792 9382
rect 37740 9318 37792 9324
rect 37464 7948 37516 7954
rect 37464 7890 37516 7896
rect 37372 6452 37424 6458
rect 37372 6394 37424 6400
rect 37280 5296 37332 5302
rect 37280 5238 37332 5244
rect 37278 4856 37334 4865
rect 37278 4791 37280 4800
rect 37332 4791 37334 4800
rect 37280 4762 37332 4768
rect 37188 4548 37240 4554
rect 37188 4490 37240 4496
rect 37476 3942 37504 7890
rect 37646 6896 37702 6905
rect 37646 6831 37648 6840
rect 37700 6831 37702 6840
rect 37648 6802 37700 6808
rect 37556 6384 37608 6390
rect 37556 6326 37608 6332
rect 37568 5710 37596 6326
rect 37752 5817 37780 9318
rect 37832 6792 37884 6798
rect 37832 6734 37884 6740
rect 37844 6322 37872 6734
rect 37832 6316 37884 6322
rect 37832 6258 37884 6264
rect 37844 6118 37872 6258
rect 38212 6186 38240 13466
rect 38568 13320 38620 13326
rect 38568 13262 38620 13268
rect 38580 9654 38608 13262
rect 38764 12986 38792 13738
rect 38752 12980 38804 12986
rect 38752 12922 38804 12928
rect 39212 12980 39264 12986
rect 39212 12922 39264 12928
rect 38752 12776 38804 12782
rect 38752 12718 38804 12724
rect 38764 10198 38792 12718
rect 38752 10192 38804 10198
rect 38752 10134 38804 10140
rect 38568 9648 38620 9654
rect 38568 9590 38620 9596
rect 38384 9444 38436 9450
rect 38384 9386 38436 9392
rect 38292 8492 38344 8498
rect 38292 8434 38344 8440
rect 38304 8022 38332 8434
rect 38292 8016 38344 8022
rect 38292 7958 38344 7964
rect 38396 6798 38424 9386
rect 38476 8900 38528 8906
rect 38476 8842 38528 8848
rect 38384 6792 38436 6798
rect 38384 6734 38436 6740
rect 38292 6316 38344 6322
rect 38292 6258 38344 6264
rect 38304 6225 38332 6258
rect 38290 6216 38346 6225
rect 38200 6180 38252 6186
rect 38290 6151 38346 6160
rect 38200 6122 38252 6128
rect 37832 6112 37884 6118
rect 37832 6054 37884 6060
rect 37738 5808 37794 5817
rect 37738 5743 37794 5752
rect 38108 5772 38160 5778
rect 38108 5714 38160 5720
rect 37556 5704 37608 5710
rect 38120 5681 38148 5714
rect 37556 5646 37608 5652
rect 38106 5672 38162 5681
rect 38106 5607 38162 5616
rect 38292 5364 38344 5370
rect 38292 5306 38344 5312
rect 38304 5166 38332 5306
rect 38292 5160 38344 5166
rect 38292 5102 38344 5108
rect 38304 4690 38332 5102
rect 38488 5098 38516 8842
rect 38660 8356 38712 8362
rect 38660 8298 38712 8304
rect 38672 8129 38700 8298
rect 39118 8256 39174 8265
rect 39118 8191 39174 8200
rect 38658 8120 38714 8129
rect 38658 8055 38714 8064
rect 38568 8016 38620 8022
rect 38568 7958 38620 7964
rect 38580 6866 38608 7958
rect 38672 7342 38700 8055
rect 39132 7886 39160 8191
rect 39224 7993 39252 12922
rect 39304 8424 39356 8430
rect 39304 8366 39356 8372
rect 39316 8022 39344 8366
rect 39488 8356 39540 8362
rect 39488 8298 39540 8304
rect 39500 8090 39528 8298
rect 39488 8084 39540 8090
rect 39488 8026 39540 8032
rect 39304 8016 39356 8022
rect 39210 7984 39266 7993
rect 39304 7958 39356 7964
rect 39210 7919 39266 7928
rect 39120 7880 39172 7886
rect 39120 7822 39172 7828
rect 39486 7576 39542 7585
rect 39396 7540 39448 7546
rect 39486 7511 39542 7520
rect 39396 7482 39448 7488
rect 39408 7449 39436 7482
rect 39500 7478 39528 7511
rect 39488 7472 39540 7478
rect 39394 7440 39450 7449
rect 39488 7414 39540 7420
rect 39394 7375 39450 7384
rect 38660 7336 38712 7342
rect 38660 7278 38712 7284
rect 38844 7336 38896 7342
rect 38844 7278 38896 7284
rect 38568 6860 38620 6866
rect 38568 6802 38620 6808
rect 38752 6180 38804 6186
rect 38752 6122 38804 6128
rect 38660 5568 38712 5574
rect 38660 5510 38712 5516
rect 38672 5098 38700 5510
rect 38384 5092 38436 5098
rect 38384 5034 38436 5040
rect 38476 5092 38528 5098
rect 38476 5034 38528 5040
rect 38660 5092 38712 5098
rect 38660 5034 38712 5040
rect 38396 4978 38424 5034
rect 38672 4978 38700 5034
rect 38396 4950 38700 4978
rect 38660 4820 38712 4826
rect 38660 4762 38712 4768
rect 38292 4684 38344 4690
rect 38292 4626 38344 4632
rect 38304 4146 38332 4626
rect 38292 4140 38344 4146
rect 38292 4082 38344 4088
rect 38200 4072 38252 4078
rect 38200 4014 38252 4020
rect 37464 3936 37516 3942
rect 37464 3878 37516 3884
rect 37476 3602 37504 3878
rect 38212 3602 38240 4014
rect 38384 4004 38436 4010
rect 38384 3946 38436 3952
rect 37464 3596 37516 3602
rect 37464 3538 37516 3544
rect 37924 3596 37976 3602
rect 37924 3538 37976 3544
rect 38200 3596 38252 3602
rect 38200 3538 38252 3544
rect 36820 2984 36872 2990
rect 36820 2926 36872 2932
rect 36728 1284 36780 1290
rect 36728 1226 36780 1232
rect 36832 800 36860 2926
rect 37556 2848 37608 2854
rect 37556 2790 37608 2796
rect 37280 2644 37332 2650
rect 37280 2586 37332 2592
rect 37188 2508 37240 2514
rect 37292 2496 37320 2586
rect 37292 2468 37412 2496
rect 37188 2450 37240 2456
rect 37200 800 37228 2450
rect 37384 2310 37412 2468
rect 37280 2304 37332 2310
rect 37280 2246 37332 2252
rect 37372 2304 37424 2310
rect 37372 2246 37424 2252
rect 37292 1766 37320 2246
rect 37280 1760 37332 1766
rect 37280 1702 37332 1708
rect 37568 800 37596 2790
rect 37936 800 37964 3538
rect 38396 2922 38424 3946
rect 38672 3194 38700 4762
rect 38660 3188 38712 3194
rect 38660 3130 38712 3136
rect 38384 2916 38436 2922
rect 38384 2858 38436 2864
rect 38660 2848 38712 2854
rect 38660 2790 38712 2796
rect 38292 2508 38344 2514
rect 38292 2450 38344 2456
rect 38304 800 38332 2450
rect 38672 800 38700 2790
rect 38764 1970 38792 6122
rect 38856 2310 38884 7278
rect 39592 7274 39620 13942
rect 39684 13870 39712 14486
rect 40972 13938 41000 16594
rect 41340 16590 41368 18022
rect 41432 16590 41460 18158
rect 42904 16794 42932 18566
rect 43352 17128 43404 17134
rect 43352 17070 43404 17076
rect 42892 16788 42944 16794
rect 42892 16730 42944 16736
rect 43364 16658 43392 17070
rect 43352 16652 43404 16658
rect 43352 16594 43404 16600
rect 41328 16584 41380 16590
rect 41328 16526 41380 16532
rect 41420 16584 41472 16590
rect 41420 16526 41472 16532
rect 41144 14068 41196 14074
rect 41144 14010 41196 14016
rect 40960 13932 41012 13938
rect 40960 13874 41012 13880
rect 39672 13864 39724 13870
rect 39672 13806 39724 13812
rect 39856 13864 39908 13870
rect 39856 13806 39908 13812
rect 39868 12434 39896 13806
rect 40132 13728 40184 13734
rect 40132 13670 40184 13676
rect 39776 12406 39896 12434
rect 39776 10130 39804 12406
rect 39764 10124 39816 10130
rect 39764 10066 39816 10072
rect 39776 9518 39804 10066
rect 39764 9512 39816 9518
rect 39764 9454 39816 9460
rect 39856 8492 39908 8498
rect 39856 8434 39908 8440
rect 39764 7404 39816 7410
rect 39764 7346 39816 7352
rect 39580 7268 39632 7274
rect 39580 7210 39632 7216
rect 39672 7268 39724 7274
rect 39672 7210 39724 7216
rect 39488 7200 39540 7206
rect 39684 7154 39712 7210
rect 39540 7148 39712 7154
rect 39488 7142 39712 7148
rect 39500 7126 39712 7142
rect 39776 6798 39804 7346
rect 39764 6792 39816 6798
rect 39764 6734 39816 6740
rect 39304 6112 39356 6118
rect 39304 6054 39356 6060
rect 39212 5092 39264 5098
rect 39212 5034 39264 5040
rect 39224 4486 39252 5034
rect 39212 4480 39264 4486
rect 39212 4422 39264 4428
rect 39120 3120 39172 3126
rect 39120 3062 39172 3068
rect 39028 3052 39080 3058
rect 39028 2994 39080 3000
rect 38844 2304 38896 2310
rect 38844 2246 38896 2252
rect 38752 1964 38804 1970
rect 38752 1906 38804 1912
rect 39040 800 39068 2994
rect 39132 2922 39160 3062
rect 39120 2916 39172 2922
rect 39120 2858 39172 2864
rect 39120 2304 39172 2310
rect 39120 2246 39172 2252
rect 39132 2106 39160 2246
rect 39120 2100 39172 2106
rect 39120 2042 39172 2048
rect 31576 536 31628 542
rect 31576 478 31628 484
rect 31666 0 31722 800
rect 32034 0 32090 800
rect 32402 0 32458 800
rect 32770 0 32826 800
rect 33138 0 33194 800
rect 33506 0 33562 800
rect 33874 0 33930 800
rect 34242 0 34298 800
rect 34610 0 34666 800
rect 34978 0 35034 800
rect 35346 0 35402 800
rect 35714 0 35770 800
rect 36082 0 36138 800
rect 36450 0 36506 800
rect 36818 0 36874 800
rect 37186 0 37242 800
rect 37554 0 37610 800
rect 37922 0 37978 800
rect 38290 0 38346 800
rect 38658 0 38714 800
rect 39026 0 39082 800
rect 39316 610 39344 6054
rect 39486 5808 39542 5817
rect 39486 5743 39488 5752
rect 39540 5743 39542 5752
rect 39488 5714 39540 5720
rect 39776 4690 39804 6734
rect 39868 5302 39896 8434
rect 39946 8120 40002 8129
rect 39946 8055 40002 8064
rect 39960 7954 39988 8055
rect 40144 7954 40172 13670
rect 40960 13320 41012 13326
rect 40960 13262 41012 13268
rect 40972 12850 41000 13262
rect 40960 12844 41012 12850
rect 40960 12786 41012 12792
rect 40868 12776 40920 12782
rect 40868 12718 40920 12724
rect 40776 10056 40828 10062
rect 40776 9998 40828 10004
rect 40592 9444 40644 9450
rect 40592 9386 40644 9392
rect 39948 7948 40000 7954
rect 39948 7890 40000 7896
rect 40132 7948 40184 7954
rect 40132 7890 40184 7896
rect 40040 7880 40092 7886
rect 39960 7828 40040 7834
rect 39960 7822 40092 7828
rect 39960 7806 40080 7822
rect 39960 7750 39988 7806
rect 39948 7744 40000 7750
rect 39948 7686 40000 7692
rect 40132 7744 40184 7750
rect 40132 7686 40184 7692
rect 40224 7744 40276 7750
rect 40224 7686 40276 7692
rect 39948 7268 40000 7274
rect 39948 7210 40000 7216
rect 39960 7041 39988 7210
rect 40038 7168 40094 7177
rect 40038 7103 40094 7112
rect 39946 7032 40002 7041
rect 39946 6967 40002 6976
rect 39960 6186 39988 6967
rect 40052 6934 40080 7103
rect 40040 6928 40092 6934
rect 40040 6870 40092 6876
rect 39948 6180 40000 6186
rect 39948 6122 40000 6128
rect 39856 5296 39908 5302
rect 39856 5238 39908 5244
rect 39764 4684 39816 4690
rect 39764 4626 39816 4632
rect 39764 4480 39816 4486
rect 39764 4422 39816 4428
rect 39776 4214 39804 4422
rect 39764 4208 39816 4214
rect 39868 4185 39896 5238
rect 39948 5092 40000 5098
rect 39948 5034 40000 5040
rect 39764 4150 39816 4156
rect 39854 4176 39910 4185
rect 39580 4140 39632 4146
rect 39854 4111 39910 4120
rect 39580 4082 39632 4088
rect 39592 3602 39620 4082
rect 39580 3596 39632 3602
rect 39580 3538 39632 3544
rect 39764 3596 39816 3602
rect 39764 3538 39816 3544
rect 39396 2304 39448 2310
rect 39396 2246 39448 2252
rect 39408 800 39436 2246
rect 39776 800 39804 3538
rect 39960 2514 39988 5034
rect 40040 5024 40092 5030
rect 40040 4966 40092 4972
rect 40052 3670 40080 4966
rect 40144 3942 40172 7686
rect 40236 4758 40264 7686
rect 40604 6458 40632 9386
rect 40684 9036 40736 9042
rect 40684 8978 40736 8984
rect 40696 7274 40724 8978
rect 40788 7546 40816 9998
rect 40880 9654 40908 12718
rect 40868 9648 40920 9654
rect 40868 9590 40920 9596
rect 41052 9104 41104 9110
rect 41052 9046 41104 9052
rect 41064 8430 41092 9046
rect 40868 8424 40920 8430
rect 40868 8366 40920 8372
rect 41052 8424 41104 8430
rect 41052 8366 41104 8372
rect 40880 8022 40908 8366
rect 41052 8288 41104 8294
rect 41052 8230 41104 8236
rect 40868 8016 40920 8022
rect 40868 7958 40920 7964
rect 41064 7857 41092 8230
rect 41050 7848 41106 7857
rect 40868 7812 40920 7818
rect 40868 7754 40920 7760
rect 40960 7812 41012 7818
rect 41050 7783 41106 7792
rect 40960 7754 41012 7760
rect 40776 7540 40828 7546
rect 40776 7482 40828 7488
rect 40880 7410 40908 7754
rect 40972 7698 41000 7754
rect 40972 7670 41092 7698
rect 40960 7540 41012 7546
rect 40960 7482 41012 7488
rect 40868 7404 40920 7410
rect 40868 7346 40920 7352
rect 40684 7268 40736 7274
rect 40684 7210 40736 7216
rect 40776 7268 40828 7274
rect 40776 7210 40828 7216
rect 40592 6452 40644 6458
rect 40592 6394 40644 6400
rect 40500 5908 40552 5914
rect 40500 5850 40552 5856
rect 40224 4752 40276 4758
rect 40224 4694 40276 4700
rect 40132 3936 40184 3942
rect 40132 3878 40184 3884
rect 40040 3664 40092 3670
rect 40040 3606 40092 3612
rect 40132 2984 40184 2990
rect 40132 2926 40184 2932
rect 39948 2508 40000 2514
rect 39948 2450 40000 2456
rect 40144 800 40172 2926
rect 40512 2582 40540 5850
rect 40788 4146 40816 7210
rect 40972 7002 41000 7482
rect 40960 6996 41012 7002
rect 40960 6938 41012 6944
rect 40868 6792 40920 6798
rect 40866 6760 40868 6769
rect 40920 6760 40922 6769
rect 40866 6695 40922 6704
rect 40880 6322 40908 6695
rect 40868 6316 40920 6322
rect 40868 6258 40920 6264
rect 40776 4140 40828 4146
rect 40776 4082 40828 4088
rect 40960 4140 41012 4146
rect 40960 4082 41012 4088
rect 40868 3596 40920 3602
rect 40868 3538 40920 3544
rect 40500 2576 40552 2582
rect 40500 2518 40552 2524
rect 40500 2304 40552 2310
rect 40500 2246 40552 2252
rect 40512 800 40540 2246
rect 40880 800 40908 3538
rect 40972 3194 41000 4082
rect 41064 3194 41092 7670
rect 41156 7002 41184 14010
rect 41432 13802 41460 16526
rect 42800 16448 42852 16454
rect 42800 16390 42852 16396
rect 41420 13796 41472 13802
rect 41420 13738 41472 13744
rect 41432 13002 41460 13738
rect 42812 13530 42840 16390
rect 42800 13524 42852 13530
rect 42800 13466 42852 13472
rect 43456 13462 43484 19110
rect 44640 18964 44692 18970
rect 44640 18906 44692 18912
rect 44088 18624 44140 18630
rect 44088 18566 44140 18572
rect 43628 17264 43680 17270
rect 43628 17206 43680 17212
rect 43640 16794 43668 17206
rect 44100 17134 44128 18566
rect 44088 17128 44140 17134
rect 44088 17070 44140 17076
rect 43628 16788 43680 16794
rect 43628 16730 43680 16736
rect 43640 16658 43668 16730
rect 43812 16720 43864 16726
rect 43812 16662 43864 16668
rect 43628 16652 43680 16658
rect 43628 16594 43680 16600
rect 43824 16046 43852 16662
rect 43812 16040 43864 16046
rect 43812 15982 43864 15988
rect 44100 15994 44128 17070
rect 44100 15978 44220 15994
rect 44100 15972 44232 15978
rect 44100 15966 44180 15972
rect 44180 15914 44232 15920
rect 43628 13932 43680 13938
rect 43628 13874 43680 13880
rect 43444 13456 43496 13462
rect 43444 13398 43496 13404
rect 42800 13388 42852 13394
rect 42800 13330 42852 13336
rect 41604 13320 41656 13326
rect 41604 13262 41656 13268
rect 41432 12986 41552 13002
rect 41432 12980 41564 12986
rect 41432 12974 41512 12980
rect 41512 12922 41564 12928
rect 41616 10198 41644 13262
rect 41972 13252 42024 13258
rect 41972 13194 42024 13200
rect 41984 12434 42012 13194
rect 42616 12980 42668 12986
rect 42616 12922 42668 12928
rect 41984 12406 42104 12434
rect 41604 10192 41656 10198
rect 41604 10134 41656 10140
rect 41420 8900 41472 8906
rect 41420 8842 41472 8848
rect 41432 8634 41460 8842
rect 41328 8628 41380 8634
rect 41328 8570 41380 8576
rect 41420 8628 41472 8634
rect 41420 8570 41472 8576
rect 41604 8628 41656 8634
rect 41604 8570 41656 8576
rect 41340 8514 41368 8570
rect 41616 8514 41644 8570
rect 41340 8486 41644 8514
rect 41236 8424 41288 8430
rect 41236 8366 41288 8372
rect 41248 8129 41276 8366
rect 41234 8120 41290 8129
rect 41234 8055 41290 8064
rect 41602 8120 41658 8129
rect 41602 8055 41658 8064
rect 41248 7886 41276 8055
rect 41616 7954 41644 8055
rect 41880 8016 41932 8022
rect 41880 7958 41932 7964
rect 41972 8016 42024 8022
rect 41972 7958 42024 7964
rect 41604 7948 41656 7954
rect 41604 7890 41656 7896
rect 41696 7948 41748 7954
rect 41696 7890 41748 7896
rect 41236 7880 41288 7886
rect 41236 7822 41288 7828
rect 41248 7410 41276 7822
rect 41512 7812 41564 7818
rect 41512 7754 41564 7760
rect 41524 7585 41552 7754
rect 41510 7576 41566 7585
rect 41510 7511 41566 7520
rect 41236 7404 41288 7410
rect 41236 7346 41288 7352
rect 41708 7342 41736 7890
rect 41892 7721 41920 7958
rect 41878 7712 41934 7721
rect 41878 7647 41934 7656
rect 41696 7336 41748 7342
rect 41694 7304 41696 7313
rect 41880 7336 41932 7342
rect 41748 7304 41750 7313
rect 41880 7278 41932 7284
rect 41694 7239 41750 7248
rect 41694 7032 41750 7041
rect 41144 6996 41196 7002
rect 41144 6938 41196 6944
rect 41236 6996 41288 7002
rect 41892 7002 41920 7278
rect 41694 6967 41750 6976
rect 41880 6996 41932 7002
rect 41236 6938 41288 6944
rect 41156 6905 41184 6938
rect 41142 6896 41198 6905
rect 41142 6831 41198 6840
rect 41144 6656 41196 6662
rect 41144 6598 41196 6604
rect 41156 6225 41184 6598
rect 41142 6216 41198 6225
rect 41142 6151 41198 6160
rect 41248 5846 41276 6938
rect 41708 6866 41736 6967
rect 41880 6938 41932 6944
rect 41878 6896 41934 6905
rect 41696 6860 41748 6866
rect 41878 6831 41880 6840
rect 41696 6802 41748 6808
rect 41932 6831 41934 6840
rect 41880 6802 41932 6808
rect 41708 6186 41736 6802
rect 41420 6180 41472 6186
rect 41420 6122 41472 6128
rect 41696 6180 41748 6186
rect 41696 6122 41748 6128
rect 41236 5840 41288 5846
rect 41236 5782 41288 5788
rect 41144 5568 41196 5574
rect 41144 5510 41196 5516
rect 40960 3188 41012 3194
rect 40960 3130 41012 3136
rect 41052 3188 41104 3194
rect 41052 3130 41104 3136
rect 41156 2582 41184 5510
rect 41432 4026 41460 6122
rect 41880 5704 41932 5710
rect 41880 5646 41932 5652
rect 41788 5636 41840 5642
rect 41788 5578 41840 5584
rect 41512 5364 41564 5370
rect 41512 5306 41564 5312
rect 41524 5030 41552 5306
rect 41512 5024 41564 5030
rect 41512 4966 41564 4972
rect 41432 3998 41552 4026
rect 41420 3664 41472 3670
rect 41420 3606 41472 3612
rect 41236 2984 41288 2990
rect 41236 2926 41288 2932
rect 41144 2576 41196 2582
rect 41144 2518 41196 2524
rect 41248 800 41276 2926
rect 41432 1630 41460 3606
rect 41420 1624 41472 1630
rect 41420 1566 41472 1572
rect 41524 1086 41552 3998
rect 41800 2514 41828 5578
rect 41892 5302 41920 5646
rect 41880 5296 41932 5302
rect 41880 5238 41932 5244
rect 41984 4826 42012 7958
rect 42076 6254 42104 12406
rect 42432 12232 42484 12238
rect 42432 12174 42484 12180
rect 42444 9654 42472 12174
rect 42524 10056 42576 10062
rect 42524 9998 42576 10004
rect 42432 9648 42484 9654
rect 42432 9590 42484 9596
rect 42432 9376 42484 9382
rect 42432 9318 42484 9324
rect 42338 7440 42394 7449
rect 42338 7375 42394 7384
rect 42156 7336 42208 7342
rect 42156 7278 42208 7284
rect 42064 6248 42116 6254
rect 42064 6190 42116 6196
rect 42168 5370 42196 7278
rect 42248 7200 42300 7206
rect 42248 7142 42300 7148
rect 42156 5364 42208 5370
rect 42156 5306 42208 5312
rect 41972 4820 42024 4826
rect 41972 4762 42024 4768
rect 42260 4078 42288 7142
rect 42352 6610 42380 7375
rect 42444 6730 42472 9318
rect 42432 6724 42484 6730
rect 42432 6666 42484 6672
rect 42352 6582 42472 6610
rect 42444 6118 42472 6582
rect 42536 6458 42564 9998
rect 42628 7449 42656 12922
rect 42812 7857 42840 13330
rect 43640 13326 43668 13874
rect 44652 13462 44680 18906
rect 46940 18896 46992 18902
rect 46940 18838 46992 18844
rect 46388 18080 46440 18086
rect 46388 18022 46440 18028
rect 46204 17128 46256 17134
rect 46204 17070 46256 17076
rect 46216 16658 46244 17070
rect 46400 16658 46428 18022
rect 46952 17338 46980 18838
rect 47032 18624 47084 18630
rect 47032 18566 47084 18572
rect 47044 18426 47072 18566
rect 47032 18420 47084 18426
rect 47032 18362 47084 18368
rect 47044 18222 47072 18362
rect 47136 18290 47164 22066
rect 50300 21244 50596 21264
rect 50356 21242 50380 21244
rect 50436 21242 50460 21244
rect 50516 21242 50540 21244
rect 50378 21190 50380 21242
rect 50442 21190 50454 21242
rect 50516 21190 50518 21242
rect 50356 21188 50380 21190
rect 50436 21188 50460 21190
rect 50516 21188 50540 21190
rect 50300 21168 50596 21188
rect 50300 20156 50596 20176
rect 50356 20154 50380 20156
rect 50436 20154 50460 20156
rect 50516 20154 50540 20156
rect 50378 20102 50380 20154
rect 50442 20102 50454 20154
rect 50516 20102 50518 20154
rect 50356 20100 50380 20102
rect 50436 20100 50460 20102
rect 50516 20100 50540 20102
rect 50300 20080 50596 20100
rect 50908 19174 50936 117098
rect 54036 116346 54064 117098
rect 54024 116340 54076 116346
rect 54024 116282 54076 116288
rect 54208 116000 54260 116006
rect 54208 115942 54260 115948
rect 50896 19168 50948 19174
rect 50896 19110 50948 19116
rect 50300 19068 50596 19088
rect 50356 19066 50380 19068
rect 50436 19066 50460 19068
rect 50516 19066 50540 19068
rect 50378 19014 50380 19066
rect 50442 19014 50454 19066
rect 50516 19014 50518 19066
rect 50356 19012 50380 19014
rect 50436 19012 50460 19014
rect 50516 19012 50540 19014
rect 50300 18992 50596 19012
rect 47860 18692 47912 18698
rect 47860 18634 47912 18640
rect 47584 18420 47636 18426
rect 47584 18362 47636 18368
rect 47124 18284 47176 18290
rect 47124 18226 47176 18232
rect 47032 18216 47084 18222
rect 47032 18158 47084 18164
rect 46940 17332 46992 17338
rect 46940 17274 46992 17280
rect 46952 16674 46980 17274
rect 46204 16652 46256 16658
rect 46204 16594 46256 16600
rect 46388 16652 46440 16658
rect 46952 16646 47072 16674
rect 46388 16594 46440 16600
rect 44732 16176 44784 16182
rect 44732 16118 44784 16124
rect 45836 16176 45888 16182
rect 45836 16118 45888 16124
rect 44744 13530 44772 16118
rect 44824 13864 44876 13870
rect 44824 13806 44876 13812
rect 44732 13524 44784 13530
rect 44732 13466 44784 13472
rect 44640 13456 44692 13462
rect 44640 13398 44692 13404
rect 43628 13320 43680 13326
rect 43628 13262 43680 13268
rect 44456 13184 44508 13190
rect 44456 13126 44508 13132
rect 43260 8356 43312 8362
rect 43260 8298 43312 8304
rect 42798 7848 42854 7857
rect 42798 7783 42854 7792
rect 42614 7440 42670 7449
rect 42614 7375 42670 7384
rect 42524 6452 42576 6458
rect 42524 6394 42576 6400
rect 42432 6112 42484 6118
rect 42432 6054 42484 6060
rect 42812 5574 42840 7783
rect 43272 5642 43300 8298
rect 43996 8016 44048 8022
rect 43996 7958 44048 7964
rect 44178 7984 44234 7993
rect 44008 7478 44036 7958
rect 44178 7919 44180 7928
rect 44232 7919 44234 7928
rect 44180 7890 44232 7896
rect 43996 7472 44048 7478
rect 43996 7414 44048 7420
rect 44180 7472 44232 7478
rect 44180 7414 44232 7420
rect 43628 7336 43680 7342
rect 43626 7304 43628 7313
rect 43680 7304 43682 7313
rect 43626 7239 43682 7248
rect 43536 6860 43588 6866
rect 43536 6802 43588 6808
rect 43548 5914 43576 6802
rect 43628 6792 43680 6798
rect 43628 6734 43680 6740
rect 44086 6760 44142 6769
rect 43536 5908 43588 5914
rect 43536 5850 43588 5856
rect 43444 5704 43496 5710
rect 43444 5646 43496 5652
rect 43260 5636 43312 5642
rect 43260 5578 43312 5584
rect 42616 5568 42668 5574
rect 42616 5510 42668 5516
rect 42800 5568 42852 5574
rect 42800 5510 42852 5516
rect 42248 4072 42300 4078
rect 42248 4014 42300 4020
rect 41972 3596 42024 3602
rect 41972 3538 42024 3544
rect 41788 2508 41840 2514
rect 41788 2450 41840 2456
rect 41604 2304 41656 2310
rect 41604 2246 41656 2252
rect 41512 1080 41564 1086
rect 41512 1022 41564 1028
rect 41616 800 41644 2246
rect 41984 800 42012 3538
rect 42340 2984 42392 2990
rect 42340 2926 42392 2932
rect 42352 800 42380 2926
rect 42628 1970 42656 5510
rect 43076 3596 43128 3602
rect 43076 3538 43128 3544
rect 42708 2304 42760 2310
rect 42708 2246 42760 2252
rect 42616 1964 42668 1970
rect 42616 1906 42668 1912
rect 42720 800 42748 2246
rect 43088 800 43116 3538
rect 43272 1834 43300 5578
rect 43456 5386 43484 5646
rect 43456 5358 43576 5386
rect 43548 5302 43576 5358
rect 43536 5296 43588 5302
rect 43536 5238 43588 5244
rect 43548 5166 43576 5238
rect 43536 5160 43588 5166
rect 43536 5102 43588 5108
rect 43548 4690 43576 5102
rect 43536 4684 43588 4690
rect 43536 4626 43588 4632
rect 43444 2984 43496 2990
rect 43444 2926 43496 2932
rect 43260 1828 43312 1834
rect 43260 1770 43312 1776
rect 43456 800 43484 2926
rect 43640 1086 43668 6734
rect 44086 6695 44088 6704
rect 44140 6695 44142 6704
rect 44088 6666 44140 6672
rect 44100 6322 44128 6666
rect 43812 6316 43864 6322
rect 44088 6316 44140 6322
rect 43864 6276 43944 6304
rect 43812 6258 43864 6264
rect 43720 6112 43772 6118
rect 43720 6054 43772 6060
rect 43732 5273 43760 6054
rect 43810 5808 43866 5817
rect 43810 5743 43812 5752
rect 43864 5743 43866 5752
rect 43812 5714 43864 5720
rect 43718 5264 43774 5273
rect 43718 5199 43774 5208
rect 43812 2304 43864 2310
rect 43812 2246 43864 2252
rect 43628 1080 43680 1086
rect 43628 1022 43680 1028
rect 43824 800 43852 2246
rect 43916 1018 43944 6276
rect 44088 6258 44140 6264
rect 44192 5166 44220 7414
rect 44468 6866 44496 13126
rect 44652 12986 44680 13398
rect 44836 13326 44864 13806
rect 45468 13388 45520 13394
rect 45468 13330 45520 13336
rect 44824 13320 44876 13326
rect 44824 13262 44876 13268
rect 44640 12980 44692 12986
rect 44640 12922 44692 12928
rect 45480 12850 45508 13330
rect 45652 12980 45704 12986
rect 45652 12922 45704 12928
rect 45468 12844 45520 12850
rect 45468 12786 45520 12792
rect 44548 12776 44600 12782
rect 44548 12718 44600 12724
rect 44560 10198 44588 12718
rect 45480 12306 45508 12786
rect 45664 12434 45692 12922
rect 45848 12850 45876 16118
rect 46216 16046 46244 16594
rect 46204 16040 46256 16046
rect 46204 15982 46256 15988
rect 46400 15978 46428 16594
rect 46940 16584 46992 16590
rect 46940 16526 46992 16532
rect 46952 16114 46980 16526
rect 46940 16108 46992 16114
rect 46940 16050 46992 16056
rect 46388 15972 46440 15978
rect 46388 15914 46440 15920
rect 47044 15910 47072 16646
rect 47216 16652 47268 16658
rect 47216 16594 47268 16600
rect 47032 15904 47084 15910
rect 47032 15846 47084 15852
rect 46940 14272 46992 14278
rect 46940 14214 46992 14220
rect 46480 13320 46532 13326
rect 46480 13262 46532 13268
rect 45836 12844 45888 12850
rect 45836 12786 45888 12792
rect 46112 12640 46164 12646
rect 46112 12582 46164 12588
rect 45572 12406 45692 12434
rect 44916 12300 44968 12306
rect 44916 12242 44968 12248
rect 45468 12300 45520 12306
rect 45468 12242 45520 12248
rect 44548 10192 44600 10198
rect 44548 10134 44600 10140
rect 44732 7744 44784 7750
rect 44732 7686 44784 7692
rect 44638 7032 44694 7041
rect 44638 6967 44694 6976
rect 44652 6866 44680 6967
rect 44456 6860 44508 6866
rect 44456 6802 44508 6808
rect 44640 6860 44692 6866
rect 44640 6802 44692 6808
rect 44364 6792 44416 6798
rect 44364 6734 44416 6740
rect 44270 6216 44326 6225
rect 44270 6151 44326 6160
rect 44180 5160 44232 5166
rect 44180 5102 44232 5108
rect 43996 5024 44048 5030
rect 43996 4966 44048 4972
rect 44008 4146 44036 4966
rect 43996 4140 44048 4146
rect 43996 4082 44048 4088
rect 44180 3596 44232 3602
rect 44180 3538 44232 3544
rect 43904 1012 43956 1018
rect 43904 954 43956 960
rect 44192 800 44220 3538
rect 44284 3058 44312 6151
rect 44272 3052 44324 3058
rect 44272 2994 44324 3000
rect 39304 604 39356 610
rect 39304 546 39356 552
rect 39394 0 39450 800
rect 39762 0 39818 800
rect 40130 0 40186 800
rect 40498 0 40554 800
rect 40866 0 40922 800
rect 41234 0 41290 800
rect 41602 0 41658 800
rect 41970 0 42026 800
rect 42338 0 42394 800
rect 42706 0 42762 800
rect 43074 0 43130 800
rect 43442 0 43498 800
rect 43810 0 43866 800
rect 44178 0 44234 800
rect 44376 134 44404 6734
rect 44468 6662 44496 6802
rect 44456 6656 44508 6662
rect 44456 6598 44508 6604
rect 44640 6248 44692 6254
rect 44640 6190 44692 6196
rect 44456 6112 44508 6118
rect 44456 6054 44508 6060
rect 44468 2514 44496 6054
rect 44548 2984 44600 2990
rect 44548 2926 44600 2932
rect 44456 2508 44508 2514
rect 44456 2450 44508 2456
rect 44560 800 44588 2926
rect 44364 128 44416 134
rect 44364 70 44416 76
rect 44546 0 44602 800
rect 44652 202 44680 6190
rect 44744 1834 44772 7686
rect 44928 7410 44956 12242
rect 45284 9988 45336 9994
rect 45284 9930 45336 9936
rect 45100 7880 45152 7886
rect 45100 7822 45152 7828
rect 44916 7404 44968 7410
rect 44916 7346 44968 7352
rect 44928 6474 44956 7346
rect 45006 7032 45062 7041
rect 45006 6967 45062 6976
rect 44836 6446 44956 6474
rect 45020 6458 45048 6967
rect 45008 6452 45060 6458
rect 44836 5234 44864 6446
rect 45008 6394 45060 6400
rect 44916 6248 44968 6254
rect 45020 6236 45048 6394
rect 44968 6208 45048 6236
rect 44916 6190 44968 6196
rect 45008 5568 45060 5574
rect 45112 5556 45140 7822
rect 45296 6866 45324 9930
rect 45572 8430 45600 12406
rect 45560 8424 45612 8430
rect 45560 8366 45612 8372
rect 46020 8424 46072 8430
rect 46020 8366 46072 8372
rect 45284 6860 45336 6866
rect 45284 6802 45336 6808
rect 45376 6724 45428 6730
rect 45376 6666 45428 6672
rect 45060 5528 45140 5556
rect 45008 5510 45060 5516
rect 44824 5228 44876 5234
rect 44824 5170 44876 5176
rect 45020 3534 45048 5510
rect 45284 5228 45336 5234
rect 45284 5170 45336 5176
rect 45296 4622 45324 5170
rect 45388 5030 45416 6666
rect 45572 6225 45600 8366
rect 45928 8288 45980 8294
rect 46032 8265 46060 8366
rect 45928 8230 45980 8236
rect 46018 8256 46074 8265
rect 45558 6216 45614 6225
rect 45558 6151 45614 6160
rect 45836 5908 45888 5914
rect 45836 5850 45888 5856
rect 45376 5024 45428 5030
rect 45376 4966 45428 4972
rect 45468 5024 45520 5030
rect 45468 4966 45520 4972
rect 45480 4826 45508 4966
rect 45468 4820 45520 4826
rect 45468 4762 45520 4768
rect 45376 4684 45428 4690
rect 45376 4626 45428 4632
rect 45284 4616 45336 4622
rect 45284 4558 45336 4564
rect 45284 3596 45336 3602
rect 45284 3538 45336 3544
rect 45008 3528 45060 3534
rect 45008 3470 45060 3476
rect 45100 3188 45152 3194
rect 45100 3130 45152 3136
rect 45112 2582 45140 3130
rect 45100 2576 45152 2582
rect 45100 2518 45152 2524
rect 45192 2576 45244 2582
rect 45192 2518 45244 2524
rect 44916 2304 44968 2310
rect 44916 2246 44968 2252
rect 44732 1828 44784 1834
rect 44732 1770 44784 1776
rect 44928 800 44956 2246
rect 45204 1970 45232 2518
rect 45192 1964 45244 1970
rect 45192 1906 45244 1912
rect 45296 800 45324 3538
rect 45388 3398 45416 4626
rect 45480 3738 45508 4762
rect 45744 4616 45796 4622
rect 45744 4558 45796 4564
rect 45756 4078 45784 4558
rect 45744 4072 45796 4078
rect 45744 4014 45796 4020
rect 45468 3732 45520 3738
rect 45468 3674 45520 3680
rect 45376 3392 45428 3398
rect 45376 3334 45428 3340
rect 45652 2984 45704 2990
rect 45652 2926 45704 2932
rect 45376 1964 45428 1970
rect 45376 1906 45428 1912
rect 45388 1834 45416 1906
rect 45376 1828 45428 1834
rect 45376 1770 45428 1776
rect 45664 800 45692 2926
rect 45848 1630 45876 5850
rect 45940 5846 45968 8230
rect 46018 8191 46074 8200
rect 46020 8084 46072 8090
rect 46020 8026 46072 8032
rect 46032 7993 46060 8026
rect 46018 7984 46074 7993
rect 46018 7919 46074 7928
rect 46124 6322 46152 12582
rect 46492 10198 46520 13262
rect 46480 10192 46532 10198
rect 46480 10134 46532 10140
rect 46204 10124 46256 10130
rect 46204 10066 46256 10072
rect 46216 6458 46244 10066
rect 46952 10062 46980 14214
rect 47228 13938 47256 16594
rect 47216 13932 47268 13938
rect 47216 13874 47268 13880
rect 47032 13864 47084 13870
rect 47032 13806 47084 13812
rect 47044 12850 47072 13806
rect 47596 13530 47624 18362
rect 47872 16658 47900 18634
rect 48320 18624 48372 18630
rect 48320 18566 48372 18572
rect 48332 18222 48360 18566
rect 54220 18222 54248 115942
rect 55600 18766 55628 117098
rect 58268 116890 58296 117098
rect 58256 116884 58308 116890
rect 58256 116826 58308 116832
rect 58440 116748 58492 116754
rect 58440 116690 58492 116696
rect 57152 116204 57204 116210
rect 57152 116146 57204 116152
rect 57164 19310 57192 116146
rect 58452 116142 58480 116690
rect 60188 116544 60240 116550
rect 60188 116486 60240 116492
rect 59268 116272 59320 116278
rect 59268 116214 59320 116220
rect 58440 116136 58492 116142
rect 58440 116078 58492 116084
rect 59280 19310 59308 116214
rect 60200 19310 60228 116486
rect 57152 19304 57204 19310
rect 57152 19246 57204 19252
rect 58072 19304 58124 19310
rect 58072 19246 58124 19252
rect 59268 19304 59320 19310
rect 60188 19304 60240 19310
rect 59268 19246 59320 19252
rect 60108 19264 60188 19292
rect 55588 18760 55640 18766
rect 55588 18702 55640 18708
rect 48320 18216 48372 18222
rect 48320 18158 48372 18164
rect 49516 18216 49568 18222
rect 49516 18158 49568 18164
rect 52460 18216 52512 18222
rect 52460 18158 52512 18164
rect 53104 18216 53156 18222
rect 53104 18158 53156 18164
rect 54208 18216 54260 18222
rect 54208 18158 54260 18164
rect 48332 17338 48360 18158
rect 48320 17332 48372 17338
rect 48320 17274 48372 17280
rect 48332 16726 48360 17274
rect 49528 17134 49556 18158
rect 49608 18080 49660 18086
rect 49608 18022 49660 18028
rect 49620 17746 49648 18022
rect 50300 17980 50596 18000
rect 50356 17978 50380 17980
rect 50436 17978 50460 17980
rect 50516 17978 50540 17980
rect 50378 17926 50380 17978
rect 50442 17926 50454 17978
rect 50516 17926 50518 17978
rect 50356 17924 50380 17926
rect 50436 17924 50460 17926
rect 50516 17924 50540 17926
rect 50300 17904 50596 17924
rect 52472 17882 52500 18158
rect 52460 17876 52512 17882
rect 52460 17818 52512 17824
rect 49608 17740 49660 17746
rect 49608 17682 49660 17688
rect 49620 17202 49648 17682
rect 49608 17196 49660 17202
rect 49608 17138 49660 17144
rect 49516 17128 49568 17134
rect 49516 17070 49568 17076
rect 49056 16992 49108 16998
rect 49056 16934 49108 16940
rect 48320 16720 48372 16726
rect 48320 16662 48372 16668
rect 47860 16652 47912 16658
rect 47780 16612 47860 16640
rect 47780 13802 47808 16612
rect 47860 16594 47912 16600
rect 48044 14068 48096 14074
rect 48044 14010 48096 14016
rect 47860 14000 47912 14006
rect 47860 13942 47912 13948
rect 47768 13796 47820 13802
rect 47768 13738 47820 13744
rect 47584 13524 47636 13530
rect 47584 13466 47636 13472
rect 47032 12844 47084 12850
rect 47032 12786 47084 12792
rect 47596 12782 47624 13466
rect 47124 12776 47176 12782
rect 47124 12718 47176 12724
rect 47584 12776 47636 12782
rect 47584 12718 47636 12724
rect 47136 12434 47164 12718
rect 47136 12406 47440 12434
rect 47216 12232 47268 12238
rect 47216 12174 47268 12180
rect 47032 10124 47084 10130
rect 47032 10066 47084 10072
rect 46940 10056 46992 10062
rect 46940 9998 46992 10004
rect 46664 9444 46716 9450
rect 46664 9386 46716 9392
rect 46296 8424 46348 8430
rect 46296 8366 46348 8372
rect 46308 8022 46336 8366
rect 46572 8288 46624 8294
rect 46386 8256 46442 8265
rect 46572 8230 46624 8236
rect 46386 8191 46442 8200
rect 46296 8016 46348 8022
rect 46296 7958 46348 7964
rect 46400 7954 46428 8191
rect 46584 7954 46612 8230
rect 46388 7948 46440 7954
rect 46388 7890 46440 7896
rect 46572 7948 46624 7954
rect 46572 7890 46624 7896
rect 46294 7848 46350 7857
rect 46294 7783 46350 7792
rect 46308 7478 46336 7783
rect 46296 7472 46348 7478
rect 46296 7414 46348 7420
rect 46204 6452 46256 6458
rect 46204 6394 46256 6400
rect 46112 6316 46164 6322
rect 46308 6304 46336 7414
rect 46400 6866 46428 7890
rect 46572 7812 46624 7818
rect 46572 7754 46624 7760
rect 46584 7478 46612 7754
rect 46572 7472 46624 7478
rect 46572 7414 46624 7420
rect 46676 7018 46704 9386
rect 46848 8084 46900 8090
rect 46848 8026 46900 8032
rect 46584 6990 46704 7018
rect 46388 6860 46440 6866
rect 46388 6802 46440 6808
rect 46478 6488 46534 6497
rect 46478 6423 46480 6432
rect 46532 6423 46534 6432
rect 46480 6394 46532 6400
rect 46112 6258 46164 6264
rect 46216 6276 46336 6304
rect 46018 5944 46074 5953
rect 46018 5879 46074 5888
rect 45928 5840 45980 5846
rect 45928 5782 45980 5788
rect 46032 5642 46060 5879
rect 46020 5636 46072 5642
rect 46020 5578 46072 5584
rect 46018 5536 46074 5545
rect 46018 5471 46074 5480
rect 46032 4622 46060 5471
rect 46112 4752 46164 4758
rect 46112 4694 46164 4700
rect 46020 4616 46072 4622
rect 46020 4558 46072 4564
rect 46124 4282 46152 4694
rect 46112 4276 46164 4282
rect 46112 4218 46164 4224
rect 46216 3466 46244 6276
rect 46584 6202 46612 6990
rect 46662 6896 46718 6905
rect 46860 6866 46888 8026
rect 46940 7880 46992 7886
rect 46940 7822 46992 7828
rect 46952 7721 46980 7822
rect 46938 7712 46994 7721
rect 46938 7647 46994 7656
rect 46938 7440 46994 7449
rect 46938 7375 46994 7384
rect 46952 7206 46980 7375
rect 46940 7200 46992 7206
rect 46940 7142 46992 7148
rect 46662 6831 46664 6840
rect 46716 6831 46718 6840
rect 46848 6860 46900 6866
rect 46664 6802 46716 6808
rect 46848 6802 46900 6808
rect 47044 6746 47072 10066
rect 47228 9654 47256 12174
rect 47216 9648 47268 9654
rect 47216 9590 47268 9596
rect 47306 8256 47362 8265
rect 47306 8191 47362 8200
rect 47320 7954 47348 8191
rect 47412 8129 47440 12406
rect 47768 10124 47820 10130
rect 47768 10066 47820 10072
rect 47780 9518 47808 10066
rect 47768 9512 47820 9518
rect 47768 9454 47820 9460
rect 47398 8120 47454 8129
rect 47398 8055 47454 8064
rect 47308 7948 47360 7954
rect 47228 7908 47308 7936
rect 47228 7585 47256 7908
rect 47308 7890 47360 7896
rect 47308 7744 47360 7750
rect 47308 7686 47360 7692
rect 47412 7698 47440 8055
rect 47492 7948 47544 7954
rect 47492 7890 47544 7896
rect 47676 7948 47728 7954
rect 47676 7890 47728 7896
rect 47504 7818 47532 7890
rect 47492 7812 47544 7818
rect 47492 7754 47544 7760
rect 47214 7576 47270 7585
rect 47214 7511 47270 7520
rect 47216 6860 47268 6866
rect 47216 6802 47268 6808
rect 46952 6718 47072 6746
rect 47124 6792 47176 6798
rect 47228 6769 47256 6802
rect 47124 6734 47176 6740
rect 47214 6760 47270 6769
rect 46846 6624 46902 6633
rect 46846 6559 46902 6568
rect 46664 6452 46716 6458
rect 46664 6394 46716 6400
rect 46676 6322 46704 6394
rect 46860 6322 46888 6559
rect 46952 6497 46980 6718
rect 46938 6488 46994 6497
rect 46938 6423 46994 6432
rect 46664 6316 46716 6322
rect 46664 6258 46716 6264
rect 46848 6316 46900 6322
rect 46848 6258 46900 6264
rect 46400 6174 46612 6202
rect 46400 5914 46428 6174
rect 46572 6112 46624 6118
rect 46572 6054 46624 6060
rect 46388 5908 46440 5914
rect 46388 5850 46440 5856
rect 46584 5556 46612 6054
rect 46676 5794 46704 6258
rect 46940 6248 46992 6254
rect 46860 6196 46940 6202
rect 46860 6190 46992 6196
rect 46860 6174 46980 6190
rect 46860 6089 46888 6174
rect 46940 6112 46992 6118
rect 46846 6080 46902 6089
rect 46940 6054 46992 6060
rect 46846 6015 46902 6024
rect 46676 5778 46888 5794
rect 46676 5772 46900 5778
rect 46676 5766 46848 5772
rect 46848 5714 46900 5720
rect 46664 5704 46716 5710
rect 46662 5672 46664 5681
rect 46716 5672 46718 5681
rect 46662 5607 46718 5616
rect 46584 5528 46796 5556
rect 46768 5370 46796 5528
rect 46756 5364 46808 5370
rect 46756 5306 46808 5312
rect 46388 5228 46440 5234
rect 46388 5170 46440 5176
rect 46400 5030 46428 5170
rect 46388 5024 46440 5030
rect 46388 4966 46440 4972
rect 46480 5024 46532 5030
rect 46480 4966 46532 4972
rect 46492 4842 46520 4966
rect 46308 4814 46520 4842
rect 46308 4690 46336 4814
rect 46952 4690 46980 6054
rect 47136 5896 47164 6734
rect 47214 6695 47270 6704
rect 47228 6390 47256 6695
rect 47216 6384 47268 6390
rect 47216 6326 47268 6332
rect 47228 5914 47256 6326
rect 47044 5868 47164 5896
rect 47216 5908 47268 5914
rect 47044 5166 47072 5868
rect 47216 5850 47268 5856
rect 47124 5772 47176 5778
rect 47124 5714 47176 5720
rect 47032 5160 47084 5166
rect 47032 5102 47084 5108
rect 47032 5024 47084 5030
rect 47032 4966 47084 4972
rect 47044 4690 47072 4966
rect 46296 4684 46348 4690
rect 46296 4626 46348 4632
rect 46940 4684 46992 4690
rect 46940 4626 46992 4632
rect 47032 4684 47084 4690
rect 47032 4626 47084 4632
rect 46388 3596 46440 3602
rect 46388 3538 46440 3544
rect 46204 3460 46256 3466
rect 46204 3402 46256 3408
rect 46020 2304 46072 2310
rect 46020 2246 46072 2252
rect 45836 1624 45888 1630
rect 45836 1566 45888 1572
rect 46032 800 46060 2246
rect 46400 800 46428 3538
rect 46756 2984 46808 2990
rect 46756 2926 46808 2932
rect 46768 800 46796 2926
rect 47136 2774 47164 5714
rect 47320 5574 47348 7686
rect 47412 7670 47532 7698
rect 47398 6896 47454 6905
rect 47398 6831 47454 6840
rect 47412 6458 47440 6831
rect 47504 6497 47532 7670
rect 47688 7426 47716 7890
rect 47688 7398 47808 7426
rect 47584 7336 47636 7342
rect 47584 7278 47636 7284
rect 47490 6488 47546 6497
rect 47400 6452 47452 6458
rect 47490 6423 47546 6432
rect 47400 6394 47452 6400
rect 47596 6390 47624 7278
rect 47676 7268 47728 7274
rect 47676 7210 47728 7216
rect 47688 7041 47716 7210
rect 47674 7032 47730 7041
rect 47674 6967 47730 6976
rect 47584 6384 47636 6390
rect 47584 6326 47636 6332
rect 47676 6248 47728 6254
rect 47676 6190 47728 6196
rect 47582 6080 47638 6089
rect 47582 6015 47638 6024
rect 47490 5944 47546 5953
rect 47400 5908 47452 5914
rect 47490 5879 47492 5888
rect 47400 5850 47452 5856
rect 47544 5879 47546 5888
rect 47492 5850 47544 5856
rect 47412 5642 47440 5850
rect 47490 5672 47546 5681
rect 47400 5636 47452 5642
rect 47490 5607 47492 5616
rect 47400 5578 47452 5584
rect 47544 5607 47546 5616
rect 47492 5578 47544 5584
rect 47308 5568 47360 5574
rect 47308 5510 47360 5516
rect 47216 5296 47268 5302
rect 47216 5238 47268 5244
rect 47398 5264 47454 5273
rect 47044 2746 47164 2774
rect 47044 2530 47072 2746
rect 47228 2582 47256 5238
rect 47398 5199 47454 5208
rect 47412 5166 47440 5199
rect 47400 5160 47452 5166
rect 47400 5102 47452 5108
rect 47492 3596 47544 3602
rect 47492 3538 47544 3544
rect 46952 2502 47072 2530
rect 47216 2576 47268 2582
rect 47216 2518 47268 2524
rect 46952 2038 46980 2502
rect 47032 2440 47084 2446
rect 47032 2382 47084 2388
rect 47044 2038 47072 2382
rect 47124 2304 47176 2310
rect 47124 2246 47176 2252
rect 46940 2032 46992 2038
rect 46940 1974 46992 1980
rect 47032 2032 47084 2038
rect 47032 1974 47084 1980
rect 47136 800 47164 2246
rect 47504 800 47532 3538
rect 47596 1698 47624 6015
rect 47688 5370 47716 6190
rect 47676 5364 47728 5370
rect 47676 5306 47728 5312
rect 47780 5234 47808 7398
rect 47872 6633 47900 13942
rect 47952 12844 48004 12850
rect 47952 12786 48004 12792
rect 47964 10198 47992 12786
rect 47952 10192 48004 10198
rect 47952 10134 48004 10140
rect 47952 8016 48004 8022
rect 47950 7984 47952 7993
rect 48004 7984 48006 7993
rect 47950 7919 48006 7928
rect 47952 6792 48004 6798
rect 47952 6734 48004 6740
rect 47858 6624 47914 6633
rect 47858 6559 47914 6568
rect 47872 6322 47900 6559
rect 47860 6316 47912 6322
rect 47860 6258 47912 6264
rect 47858 6216 47914 6225
rect 47858 6151 47860 6160
rect 47912 6151 47914 6160
rect 47860 6122 47912 6128
rect 47860 5568 47912 5574
rect 47858 5536 47860 5545
rect 47912 5536 47914 5545
rect 47858 5471 47914 5480
rect 47768 5228 47820 5234
rect 47768 5170 47820 5176
rect 47860 2984 47912 2990
rect 47860 2926 47912 2932
rect 47584 1692 47636 1698
rect 47584 1634 47636 1640
rect 47872 800 47900 2926
rect 47964 1834 47992 6734
rect 48056 5778 48084 14010
rect 49068 13938 49096 16934
rect 49056 13932 49108 13938
rect 49056 13874 49108 13880
rect 49424 13932 49476 13938
rect 49424 13874 49476 13880
rect 48412 13796 48464 13802
rect 48412 13738 48464 13744
rect 48424 12102 48452 13738
rect 48780 13388 48832 13394
rect 48780 13330 48832 13336
rect 48596 13184 48648 13190
rect 48596 13126 48648 13132
rect 48412 12096 48464 12102
rect 48412 12038 48464 12044
rect 48424 9178 48452 12038
rect 48412 9172 48464 9178
rect 48412 9114 48464 9120
rect 48504 8016 48556 8022
rect 48502 7984 48504 7993
rect 48556 7984 48558 7993
rect 48412 7948 48464 7954
rect 48502 7919 48558 7928
rect 48412 7890 48464 7896
rect 48136 7744 48188 7750
rect 48136 7686 48188 7692
rect 48044 5772 48096 5778
rect 48044 5714 48096 5720
rect 48044 5568 48096 5574
rect 48044 5510 48096 5516
rect 48056 3126 48084 5510
rect 48148 4826 48176 7686
rect 48424 7342 48452 7890
rect 48412 7336 48464 7342
rect 48412 7278 48464 7284
rect 48228 7268 48280 7274
rect 48228 7210 48280 7216
rect 48136 4820 48188 4826
rect 48136 4762 48188 4768
rect 48240 3942 48268 7210
rect 48608 6866 48636 13126
rect 48792 12782 48820 13330
rect 49436 13326 49464 13874
rect 49528 13734 49556 17070
rect 50300 16892 50596 16912
rect 50356 16890 50380 16892
rect 50436 16890 50460 16892
rect 50516 16890 50540 16892
rect 50378 16838 50380 16890
rect 50442 16838 50454 16890
rect 50516 16838 50518 16890
rect 50356 16836 50380 16838
rect 50436 16836 50460 16838
rect 50516 16836 50540 16838
rect 50300 16816 50596 16836
rect 52736 16652 52788 16658
rect 52736 16594 52788 16600
rect 50300 15804 50596 15824
rect 50356 15802 50380 15804
rect 50436 15802 50460 15804
rect 50516 15802 50540 15804
rect 50378 15750 50380 15802
rect 50442 15750 50454 15802
rect 50516 15750 50518 15802
rect 50356 15748 50380 15750
rect 50436 15748 50460 15750
rect 50516 15748 50540 15750
rect 50300 15728 50596 15748
rect 50300 14716 50596 14736
rect 50356 14714 50380 14716
rect 50436 14714 50460 14716
rect 50516 14714 50540 14716
rect 50378 14662 50380 14714
rect 50442 14662 50454 14714
rect 50516 14662 50518 14714
rect 50356 14660 50380 14662
rect 50436 14660 50460 14662
rect 50516 14660 50540 14662
rect 50300 14640 50596 14660
rect 49516 13728 49568 13734
rect 49516 13670 49568 13676
rect 50620 13728 50672 13734
rect 50620 13670 50672 13676
rect 50300 13628 50596 13648
rect 50356 13626 50380 13628
rect 50436 13626 50460 13628
rect 50516 13626 50540 13628
rect 50378 13574 50380 13626
rect 50442 13574 50454 13626
rect 50516 13574 50518 13626
rect 50356 13572 50380 13574
rect 50436 13572 50460 13574
rect 50516 13572 50540 13574
rect 50300 13552 50596 13572
rect 49424 13320 49476 13326
rect 49424 13262 49476 13268
rect 48780 12776 48832 12782
rect 48780 12718 48832 12724
rect 50632 12714 50660 13670
rect 52748 13530 52776 16594
rect 53116 16590 53144 18158
rect 54220 16658 54248 18158
rect 54392 18148 54444 18154
rect 54392 18090 54444 18096
rect 54404 16726 54432 18090
rect 56692 17060 56744 17066
rect 56692 17002 56744 17008
rect 56968 17060 57020 17066
rect 56968 17002 57020 17008
rect 54392 16720 54444 16726
rect 54392 16662 54444 16668
rect 56704 16658 56732 17002
rect 53196 16652 53248 16658
rect 53196 16594 53248 16600
rect 54208 16652 54260 16658
rect 54208 16594 54260 16600
rect 56692 16652 56744 16658
rect 56692 16594 56744 16600
rect 56876 16652 56928 16658
rect 56876 16594 56928 16600
rect 53104 16584 53156 16590
rect 53104 16526 53156 16532
rect 52736 13524 52788 13530
rect 52736 13466 52788 13472
rect 53208 13394 53236 16594
rect 56692 16448 56744 16454
rect 56692 16390 56744 16396
rect 56704 16114 56732 16390
rect 56692 16108 56744 16114
rect 56692 16050 56744 16056
rect 56704 15638 56732 16050
rect 56888 15706 56916 16594
rect 56876 15700 56928 15706
rect 56876 15642 56928 15648
rect 56692 15632 56744 15638
rect 56692 15574 56744 15580
rect 56980 15570 57008 17002
rect 57060 15904 57112 15910
rect 57060 15846 57112 15852
rect 56968 15564 57020 15570
rect 56968 15506 57020 15512
rect 55312 15360 55364 15366
rect 55312 15302 55364 15308
rect 55220 14340 55272 14346
rect 55220 14282 55272 14288
rect 55232 13870 55260 14282
rect 55220 13864 55272 13870
rect 55220 13806 55272 13812
rect 55324 13530 55352 15302
rect 56600 14000 56652 14006
rect 56600 13942 56652 13948
rect 55404 13864 55456 13870
rect 55404 13806 55456 13812
rect 55312 13524 55364 13530
rect 55312 13466 55364 13472
rect 52276 13388 52328 13394
rect 52276 13330 52328 13336
rect 53196 13388 53248 13394
rect 53196 13330 53248 13336
rect 55220 13388 55272 13394
rect 55220 13330 55272 13336
rect 50988 12776 51040 12782
rect 50988 12718 51040 12724
rect 50620 12708 50672 12714
rect 50620 12650 50672 12656
rect 50300 12540 50596 12560
rect 50356 12538 50380 12540
rect 50436 12538 50460 12540
rect 50516 12538 50540 12540
rect 50378 12486 50380 12538
rect 50442 12486 50454 12538
rect 50516 12486 50518 12538
rect 50356 12484 50380 12486
rect 50436 12484 50460 12486
rect 50516 12484 50540 12486
rect 50300 12464 50596 12484
rect 50300 11452 50596 11472
rect 50356 11450 50380 11452
rect 50436 11450 50460 11452
rect 50516 11450 50540 11452
rect 50378 11398 50380 11450
rect 50442 11398 50454 11450
rect 50516 11398 50518 11450
rect 50356 11396 50380 11398
rect 50436 11396 50460 11398
rect 50516 11396 50540 11398
rect 50300 11376 50596 11396
rect 50300 10364 50596 10384
rect 50356 10362 50380 10364
rect 50436 10362 50460 10364
rect 50516 10362 50540 10364
rect 50378 10310 50380 10362
rect 50442 10310 50454 10362
rect 50516 10310 50518 10362
rect 50356 10308 50380 10310
rect 50436 10308 50460 10310
rect 50516 10308 50540 10310
rect 50300 10288 50596 10308
rect 50632 9586 50660 12650
rect 51000 9654 51028 12718
rect 52288 12646 52316 13330
rect 54668 13184 54720 13190
rect 54668 13126 54720 13132
rect 54944 13184 54996 13190
rect 54944 13126 54996 13132
rect 52276 12640 52328 12646
rect 52276 12582 52328 12588
rect 50988 9648 51040 9654
rect 50988 9590 51040 9596
rect 49700 9580 49752 9586
rect 49700 9522 49752 9528
rect 50620 9580 50672 9586
rect 50620 9522 50672 9528
rect 49424 9444 49476 9450
rect 49424 9386 49476 9392
rect 48688 8016 48740 8022
rect 48688 7958 48740 7964
rect 48700 7857 48728 7958
rect 49148 7948 49200 7954
rect 49148 7890 49200 7896
rect 48686 7848 48742 7857
rect 48686 7783 48742 7792
rect 48780 7744 48832 7750
rect 48780 7686 48832 7692
rect 49056 7744 49108 7750
rect 49056 7686 49108 7692
rect 48792 7426 48820 7686
rect 48700 7410 48820 7426
rect 49068 7410 49096 7686
rect 48688 7404 48820 7410
rect 48740 7398 48820 7404
rect 49056 7404 49108 7410
rect 48688 7346 48740 7352
rect 49056 7346 49108 7352
rect 49160 7342 49188 7890
rect 49330 7576 49386 7585
rect 49330 7511 49386 7520
rect 49240 7472 49292 7478
rect 49238 7440 49240 7449
rect 49292 7440 49294 7449
rect 49238 7375 49294 7384
rect 49344 7342 49372 7511
rect 48872 7336 48924 7342
rect 48872 7278 48924 7284
rect 49148 7336 49200 7342
rect 49148 7278 49200 7284
rect 49332 7336 49384 7342
rect 49332 7278 49384 7284
rect 48596 6860 48648 6866
rect 48596 6802 48648 6808
rect 48504 6792 48556 6798
rect 48504 6734 48556 6740
rect 48320 4480 48372 4486
rect 48320 4422 48372 4428
rect 48228 3936 48280 3942
rect 48228 3878 48280 3884
rect 48044 3120 48096 3126
rect 48044 3062 48096 3068
rect 48332 2922 48360 4422
rect 48320 2916 48372 2922
rect 48320 2858 48372 2864
rect 48516 2774 48544 6734
rect 48608 6662 48636 6802
rect 48780 6792 48832 6798
rect 48780 6734 48832 6740
rect 48884 6780 48912 7278
rect 49160 7177 49188 7278
rect 49332 7200 49384 7206
rect 49146 7168 49202 7177
rect 49332 7142 49384 7148
rect 49146 7103 49202 7112
rect 48964 6792 49016 6798
rect 48884 6752 48964 6780
rect 48596 6656 48648 6662
rect 48596 6598 48648 6604
rect 48792 6390 48820 6734
rect 48780 6384 48832 6390
rect 48780 6326 48832 6332
rect 48596 6316 48648 6322
rect 48596 6258 48648 6264
rect 48608 4486 48636 6258
rect 48780 6248 48832 6254
rect 48884 6236 48912 6752
rect 48964 6734 49016 6740
rect 48962 6624 49018 6633
rect 48962 6559 49018 6568
rect 48976 6458 49004 6559
rect 48964 6452 49016 6458
rect 48964 6394 49016 6400
rect 49056 6452 49108 6458
rect 49056 6394 49108 6400
rect 48832 6208 48912 6236
rect 48962 6216 49018 6225
rect 48780 6190 48832 6196
rect 48688 6180 48740 6186
rect 48688 6122 48740 6128
rect 48700 6089 48728 6122
rect 48686 6080 48742 6089
rect 48686 6015 48742 6024
rect 48792 5817 48820 6190
rect 48962 6151 48964 6160
rect 49016 6151 49018 6160
rect 48964 6122 49016 6128
rect 48778 5808 48834 5817
rect 49068 5778 49096 6394
rect 49160 6236 49188 7103
rect 49240 6248 49292 6254
rect 49160 6208 49240 6236
rect 49240 6190 49292 6196
rect 48778 5743 48834 5752
rect 49056 5772 49108 5778
rect 49056 5714 49108 5720
rect 48596 4480 48648 4486
rect 48596 4422 48648 4428
rect 49344 4010 49372 7142
rect 49436 6866 49464 9386
rect 49712 8838 49740 9522
rect 50300 9276 50596 9296
rect 50356 9274 50380 9276
rect 50436 9274 50460 9276
rect 50516 9274 50540 9276
rect 50378 9222 50380 9274
rect 50442 9222 50454 9274
rect 50516 9222 50518 9274
rect 50356 9220 50380 9222
rect 50436 9220 50460 9222
rect 50516 9220 50540 9222
rect 50300 9200 50596 9220
rect 52092 9172 52144 9178
rect 52092 9114 52144 9120
rect 49700 8832 49752 8838
rect 49700 8774 49752 8780
rect 50300 8188 50596 8208
rect 50356 8186 50380 8188
rect 50436 8186 50460 8188
rect 50516 8186 50540 8188
rect 50378 8134 50380 8186
rect 50442 8134 50454 8186
rect 50516 8134 50518 8186
rect 50356 8132 50380 8134
rect 50436 8132 50460 8134
rect 50516 8132 50540 8134
rect 50300 8112 50596 8132
rect 49976 7948 50028 7954
rect 49976 7890 50028 7896
rect 49988 7342 50016 7890
rect 50988 7812 51040 7818
rect 50988 7754 51040 7760
rect 51000 7546 51028 7754
rect 50896 7540 50948 7546
rect 50896 7482 50948 7488
rect 50988 7540 51040 7546
rect 50988 7482 51040 7488
rect 50908 7449 50936 7482
rect 50894 7440 50950 7449
rect 50894 7375 50950 7384
rect 51078 7440 51134 7449
rect 51078 7375 51134 7384
rect 49976 7336 50028 7342
rect 49976 7278 50028 7284
rect 50160 7336 50212 7342
rect 50160 7278 50212 7284
rect 49608 7268 49660 7274
rect 49608 7210 49660 7216
rect 49424 6860 49476 6866
rect 49424 6802 49476 6808
rect 49516 6656 49568 6662
rect 49516 6598 49568 6604
rect 49424 6248 49476 6254
rect 49424 6190 49476 6196
rect 49436 5914 49464 6190
rect 49424 5908 49476 5914
rect 49424 5850 49476 5856
rect 49528 5846 49556 6598
rect 49516 5840 49568 5846
rect 49516 5782 49568 5788
rect 49620 4690 49648 7210
rect 50172 7177 50200 7278
rect 50620 7200 50672 7206
rect 50158 7168 50214 7177
rect 50620 7142 50672 7148
rect 50158 7103 50214 7112
rect 49976 6928 50028 6934
rect 49976 6870 50028 6876
rect 49790 6488 49846 6497
rect 49790 6423 49846 6432
rect 49804 6322 49832 6423
rect 49792 6316 49844 6322
rect 49792 6258 49844 6264
rect 49792 6112 49844 6118
rect 49792 6054 49844 6060
rect 49608 4684 49660 4690
rect 49608 4626 49660 4632
rect 49332 4004 49384 4010
rect 49332 3946 49384 3952
rect 48596 3596 48648 3602
rect 48596 3538 48648 3544
rect 49700 3596 49752 3602
rect 49700 3538 49752 3544
rect 48424 2746 48544 2774
rect 48320 2508 48372 2514
rect 48320 2450 48372 2456
rect 48228 2304 48280 2310
rect 48228 2246 48280 2252
rect 47952 1828 48004 1834
rect 47952 1770 48004 1776
rect 48240 800 48268 2246
rect 48332 1970 48360 2450
rect 48320 1964 48372 1970
rect 48320 1906 48372 1912
rect 44640 196 44692 202
rect 44640 138 44692 144
rect 44914 0 44970 800
rect 45282 0 45338 800
rect 45650 0 45706 800
rect 46018 0 46074 800
rect 46386 0 46442 800
rect 46754 0 46810 800
rect 47122 0 47178 800
rect 47490 0 47546 800
rect 47858 0 47914 800
rect 48226 0 48282 800
rect 48424 406 48452 2746
rect 48608 800 48636 3538
rect 48964 2984 49016 2990
rect 48964 2926 49016 2932
rect 48976 800 49004 2926
rect 49332 2304 49384 2310
rect 49332 2246 49384 2252
rect 49344 800 49372 2246
rect 49712 800 49740 3538
rect 49804 2582 49832 6054
rect 49988 5574 50016 6870
rect 50068 6860 50120 6866
rect 50172 6848 50200 7103
rect 50300 7100 50596 7120
rect 50356 7098 50380 7100
rect 50436 7098 50460 7100
rect 50516 7098 50540 7100
rect 50378 7046 50380 7098
rect 50442 7046 50454 7098
rect 50516 7046 50518 7098
rect 50356 7044 50380 7046
rect 50436 7044 50460 7046
rect 50516 7044 50540 7046
rect 50300 7024 50596 7044
rect 50252 6860 50304 6866
rect 50172 6820 50252 6848
rect 50068 6802 50120 6808
rect 50252 6802 50304 6808
rect 50080 6497 50108 6802
rect 50066 6488 50122 6497
rect 50066 6423 50122 6432
rect 50068 6248 50120 6254
rect 50068 6190 50120 6196
rect 50080 6089 50108 6190
rect 50066 6080 50122 6089
rect 50066 6015 50122 6024
rect 50300 6012 50596 6032
rect 50356 6010 50380 6012
rect 50436 6010 50460 6012
rect 50516 6010 50540 6012
rect 50378 5958 50380 6010
rect 50442 5958 50454 6010
rect 50516 5958 50518 6010
rect 50356 5956 50380 5958
rect 50436 5956 50460 5958
rect 50516 5956 50540 5958
rect 50300 5936 50596 5956
rect 49976 5568 50028 5574
rect 49976 5510 50028 5516
rect 50632 5098 50660 7142
rect 51092 6322 51120 7375
rect 51816 6792 51868 6798
rect 51816 6734 51868 6740
rect 51632 6384 51684 6390
rect 51632 6326 51684 6332
rect 51080 6316 51132 6322
rect 51080 6258 51132 6264
rect 50988 6112 51040 6118
rect 50988 6054 51040 6060
rect 50620 5092 50672 5098
rect 50620 5034 50672 5040
rect 49884 5024 49936 5030
rect 49884 4966 49936 4972
rect 49792 2576 49844 2582
rect 49792 2518 49844 2524
rect 49896 2514 49924 4966
rect 50300 4924 50596 4944
rect 50356 4922 50380 4924
rect 50436 4922 50460 4924
rect 50516 4922 50540 4924
rect 50378 4870 50380 4922
rect 50442 4870 50454 4922
rect 50516 4870 50518 4922
rect 50356 4868 50380 4870
rect 50436 4868 50460 4870
rect 50516 4868 50540 4870
rect 50300 4848 50596 4868
rect 50300 3836 50596 3856
rect 50356 3834 50380 3836
rect 50436 3834 50460 3836
rect 50516 3834 50540 3836
rect 50378 3782 50380 3834
rect 50442 3782 50454 3834
rect 50516 3782 50518 3834
rect 50356 3780 50380 3782
rect 50436 3780 50460 3782
rect 50516 3780 50540 3782
rect 50300 3760 50596 3780
rect 50068 2984 50120 2990
rect 50068 2926 50120 2932
rect 50804 2984 50856 2990
rect 50804 2926 50856 2932
rect 49884 2508 49936 2514
rect 49884 2450 49936 2456
rect 50080 800 50108 2926
rect 50300 2748 50596 2768
rect 50356 2746 50380 2748
rect 50436 2746 50460 2748
rect 50516 2746 50540 2748
rect 50378 2694 50380 2746
rect 50442 2694 50454 2746
rect 50516 2694 50518 2746
rect 50356 2692 50380 2694
rect 50436 2692 50460 2694
rect 50516 2692 50540 2694
rect 50300 2672 50596 2692
rect 50436 2304 50488 2310
rect 50436 2246 50488 2252
rect 50448 800 50476 2246
rect 50816 800 50844 2926
rect 51000 2582 51028 6054
rect 51644 4214 51672 6326
rect 51828 4282 51856 6734
rect 52104 5778 52132 9114
rect 52184 6724 52236 6730
rect 52184 6666 52236 6672
rect 52092 5772 52144 5778
rect 52092 5714 52144 5720
rect 52196 5710 52224 6666
rect 52288 6322 52316 12582
rect 54484 9580 54536 9586
rect 54484 9522 54536 9528
rect 53472 9444 53524 9450
rect 53472 9386 53524 9392
rect 53484 6866 53512 9386
rect 54300 8356 54352 8362
rect 54300 8298 54352 8304
rect 52828 6860 52880 6866
rect 52828 6802 52880 6808
rect 53472 6860 53524 6866
rect 53472 6802 53524 6808
rect 52552 6792 52604 6798
rect 52552 6734 52604 6740
rect 52276 6316 52328 6322
rect 52276 6258 52328 6264
rect 52184 5704 52236 5710
rect 52184 5646 52236 5652
rect 52196 4758 52224 5646
rect 52184 4752 52236 4758
rect 52184 4694 52236 4700
rect 51816 4276 51868 4282
rect 51816 4218 51868 4224
rect 51632 4208 51684 4214
rect 51632 4150 51684 4156
rect 51908 2984 51960 2990
rect 51908 2926 51960 2932
rect 52276 2984 52328 2990
rect 52276 2926 52328 2932
rect 50988 2576 51040 2582
rect 50988 2518 51040 2524
rect 51172 2508 51224 2514
rect 51172 2450 51224 2456
rect 51184 800 51212 2450
rect 51540 2304 51592 2310
rect 51540 2246 51592 2252
rect 51552 800 51580 2246
rect 51920 800 51948 2926
rect 52288 800 52316 2926
rect 48412 400 48464 406
rect 48412 342 48464 348
rect 48594 0 48650 800
rect 48962 0 49018 800
rect 49330 0 49386 800
rect 49698 0 49754 800
rect 50066 0 50122 800
rect 50434 0 50490 800
rect 50802 0 50858 800
rect 51170 0 51226 800
rect 51538 0 51594 800
rect 51906 0 51962 800
rect 52274 0 52330 800
rect 52564 338 52592 6734
rect 52840 6390 52868 6802
rect 54024 6792 54076 6798
rect 53944 6752 54024 6780
rect 52828 6384 52880 6390
rect 52828 6326 52880 6332
rect 53840 6180 53892 6186
rect 53840 6122 53892 6128
rect 53104 6112 53156 6118
rect 53104 6054 53156 6060
rect 52828 5568 52880 5574
rect 52828 5510 52880 5516
rect 52920 5568 52972 5574
rect 52920 5510 52972 5516
rect 52840 2582 52868 5510
rect 52828 2576 52880 2582
rect 52828 2518 52880 2524
rect 52644 2304 52696 2310
rect 52644 2246 52696 2252
rect 52656 800 52684 2246
rect 52552 332 52604 338
rect 52552 274 52604 280
rect 52642 0 52698 800
rect 52932 474 52960 5510
rect 53012 2984 53064 2990
rect 53012 2926 53064 2932
rect 53024 800 53052 2926
rect 53116 2514 53144 6054
rect 53194 5808 53250 5817
rect 53194 5743 53196 5752
rect 53248 5743 53250 5752
rect 53196 5714 53248 5720
rect 53852 5710 53880 6122
rect 53840 5704 53892 5710
rect 53840 5646 53892 5652
rect 53944 4758 53972 6752
rect 54024 6734 54076 6740
rect 54206 6488 54262 6497
rect 54206 6423 54262 6432
rect 54220 6118 54248 6423
rect 54024 6112 54076 6118
rect 54024 6054 54076 6060
rect 54208 6112 54260 6118
rect 54208 6054 54260 6060
rect 53932 4752 53984 4758
rect 53932 4694 53984 4700
rect 53380 2984 53432 2990
rect 53380 2926 53432 2932
rect 53104 2508 53156 2514
rect 53104 2450 53156 2456
rect 53288 2440 53340 2446
rect 53288 2382 53340 2388
rect 53300 1834 53328 2382
rect 53288 1828 53340 1834
rect 53288 1770 53340 1776
rect 53392 800 53420 2926
rect 54036 2582 54064 6054
rect 54312 5817 54340 8298
rect 54496 6254 54524 9522
rect 54680 6798 54708 13126
rect 54760 9376 54812 9382
rect 54760 9318 54812 9324
rect 54772 9042 54800 9318
rect 54760 9036 54812 9042
rect 54760 8978 54812 8984
rect 54760 8016 54812 8022
rect 54760 7958 54812 7964
rect 54772 7478 54800 7958
rect 54760 7472 54812 7478
rect 54760 7414 54812 7420
rect 54956 6866 54984 13126
rect 55128 12776 55180 12782
rect 55128 12718 55180 12724
rect 55140 9654 55168 12718
rect 55128 9648 55180 9654
rect 55128 9590 55180 9596
rect 55036 9036 55088 9042
rect 55036 8978 55088 8984
rect 54944 6860 54996 6866
rect 54944 6802 54996 6808
rect 54668 6792 54720 6798
rect 54668 6734 54720 6740
rect 54852 6792 54904 6798
rect 54852 6734 54904 6740
rect 54576 6724 54628 6730
rect 54576 6666 54628 6672
rect 54484 6248 54536 6254
rect 54484 6190 54536 6196
rect 54588 6186 54616 6666
rect 54760 6384 54812 6390
rect 54760 6326 54812 6332
rect 54576 6180 54628 6186
rect 54576 6122 54628 6128
rect 54298 5808 54354 5817
rect 54298 5743 54300 5752
rect 54352 5743 54354 5752
rect 54300 5714 54352 5720
rect 54312 5683 54340 5714
rect 54772 5710 54800 6326
rect 54760 5704 54812 5710
rect 54760 5646 54812 5652
rect 54116 3596 54168 3602
rect 54116 3538 54168 3544
rect 54024 2576 54076 2582
rect 54024 2518 54076 2524
rect 53748 2304 53800 2310
rect 53748 2246 53800 2252
rect 53760 800 53788 2246
rect 54128 800 54156 3538
rect 54484 2984 54536 2990
rect 54484 2926 54536 2932
rect 54496 800 54524 2926
rect 54864 2774 54892 6734
rect 54956 6662 54984 6802
rect 54944 6656 54996 6662
rect 54944 6598 54996 6604
rect 55048 5914 55076 8978
rect 55232 7818 55260 13330
rect 55416 9586 55444 13806
rect 55772 12232 55824 12238
rect 55772 12174 55824 12180
rect 55404 9580 55456 9586
rect 55404 9522 55456 9528
rect 55784 8974 55812 12174
rect 56508 10124 56560 10130
rect 56508 10066 56560 10072
rect 56520 9586 56548 10066
rect 56508 9580 56560 9586
rect 56508 9522 56560 9528
rect 56232 9444 56284 9450
rect 56232 9386 56284 9392
rect 55772 8968 55824 8974
rect 55772 8910 55824 8916
rect 55680 8288 55732 8294
rect 55680 8230 55732 8236
rect 55772 8288 55824 8294
rect 55772 8230 55824 8236
rect 55220 7812 55272 7818
rect 55220 7754 55272 7760
rect 55128 7404 55180 7410
rect 55128 7346 55180 7352
rect 55140 6662 55168 7346
rect 55232 7342 55260 7754
rect 55496 7404 55548 7410
rect 55496 7346 55548 7352
rect 55220 7336 55272 7342
rect 55220 7278 55272 7284
rect 55312 6792 55364 6798
rect 55312 6734 55364 6740
rect 55128 6656 55180 6662
rect 55128 6598 55180 6604
rect 55324 6390 55352 6734
rect 55312 6384 55364 6390
rect 55312 6326 55364 6332
rect 55508 6186 55536 7346
rect 55692 6934 55720 8230
rect 55784 8090 55812 8230
rect 55772 8084 55824 8090
rect 55772 8026 55824 8032
rect 55864 8084 55916 8090
rect 55864 8026 55916 8032
rect 55876 7993 55904 8026
rect 55862 7984 55918 7993
rect 55862 7919 55918 7928
rect 55772 7336 55824 7342
rect 55772 7278 55824 7284
rect 56048 7336 56100 7342
rect 56048 7278 56100 7284
rect 55680 6928 55732 6934
rect 55680 6870 55732 6876
rect 55680 6316 55732 6322
rect 55680 6258 55732 6264
rect 55496 6180 55548 6186
rect 55496 6122 55548 6128
rect 55036 5908 55088 5914
rect 55036 5850 55088 5856
rect 55692 5778 55720 6258
rect 55680 5772 55732 5778
rect 55680 5714 55732 5720
rect 55220 3596 55272 3602
rect 55220 3538 55272 3544
rect 54772 2746 54892 2774
rect 54772 882 54800 2746
rect 54852 2304 54904 2310
rect 54852 2246 54904 2252
rect 54760 876 54812 882
rect 54760 818 54812 824
rect 54864 800 54892 2246
rect 55232 800 55260 3538
rect 55588 2984 55640 2990
rect 55588 2926 55640 2932
rect 55600 800 55628 2926
rect 52920 468 52972 474
rect 52920 410 52972 416
rect 53010 0 53066 800
rect 53378 0 53434 800
rect 53746 0 53802 800
rect 54114 0 54170 800
rect 54482 0 54538 800
rect 54850 0 54906 800
rect 55218 0 55274 800
rect 55586 0 55642 800
rect 55784 270 55812 7278
rect 56060 6730 56088 7278
rect 56244 6866 56272 9386
rect 56612 7410 56640 13942
rect 56692 13728 56744 13734
rect 56692 13670 56744 13676
rect 56704 13258 56732 13670
rect 56692 13252 56744 13258
rect 56692 13194 56744 13200
rect 56704 12850 56732 13194
rect 57072 12850 57100 15846
rect 57164 13394 57192 19246
rect 57244 19168 57296 19174
rect 57244 19110 57296 19116
rect 57256 17270 57284 19110
rect 57244 17264 57296 17270
rect 57244 17206 57296 17212
rect 57256 16658 57284 17206
rect 57244 16652 57296 16658
rect 57244 16594 57296 16600
rect 58084 16046 58112 19246
rect 59360 19168 59412 19174
rect 59360 19110 59412 19116
rect 58348 17604 58400 17610
rect 58348 17546 58400 17552
rect 59176 17604 59228 17610
rect 59176 17546 59228 17552
rect 58360 17134 58388 17546
rect 58348 17128 58400 17134
rect 58348 17070 58400 17076
rect 58256 16652 58308 16658
rect 58256 16594 58308 16600
rect 58716 16652 58768 16658
rect 58716 16594 58768 16600
rect 58072 16040 58124 16046
rect 58072 15982 58124 15988
rect 57244 14068 57296 14074
rect 57244 14010 57296 14016
rect 57152 13388 57204 13394
rect 57152 13330 57204 13336
rect 57164 12986 57192 13330
rect 57152 12980 57204 12986
rect 57152 12922 57204 12928
rect 56692 12844 56744 12850
rect 56692 12786 56744 12792
rect 57060 12844 57112 12850
rect 57060 12786 57112 12792
rect 56704 12306 56732 12786
rect 56968 12640 57020 12646
rect 56968 12582 57020 12588
rect 56692 12300 56744 12306
rect 56692 12242 56744 12248
rect 56876 9920 56928 9926
rect 56876 9862 56928 9868
rect 56888 9518 56916 9862
rect 56876 9512 56928 9518
rect 56876 9454 56928 9460
rect 56888 9042 56916 9454
rect 56876 9036 56928 9042
rect 56876 8978 56928 8984
rect 56980 8362 57008 12582
rect 57060 9444 57112 9450
rect 57060 9386 57112 9392
rect 56968 8356 57020 8362
rect 56968 8298 57020 8304
rect 56692 7880 56744 7886
rect 56692 7822 56744 7828
rect 56600 7404 56652 7410
rect 56600 7346 56652 7352
rect 56704 7342 56732 7822
rect 56876 7812 56928 7818
rect 56876 7754 56928 7760
rect 56692 7336 56744 7342
rect 56692 7278 56744 7284
rect 56600 7268 56652 7274
rect 56600 7210 56652 7216
rect 56612 7002 56640 7210
rect 56600 6996 56652 7002
rect 56600 6938 56652 6944
rect 56888 6866 56916 7754
rect 57072 7546 57100 9386
rect 57060 7540 57112 7546
rect 57060 7482 57112 7488
rect 56232 6860 56284 6866
rect 56232 6802 56284 6808
rect 56876 6860 56928 6866
rect 56876 6802 56928 6808
rect 56048 6724 56100 6730
rect 56048 6666 56100 6672
rect 56060 6390 56088 6666
rect 56048 6384 56100 6390
rect 56048 6326 56100 6332
rect 57256 6322 57284 14010
rect 57520 13388 57572 13394
rect 57520 13330 57572 13336
rect 57980 13388 58032 13394
rect 57980 13330 58032 13336
rect 57532 13190 57560 13330
rect 57612 13320 57664 13326
rect 57612 13262 57664 13268
rect 57520 13184 57572 13190
rect 57520 13126 57572 13132
rect 57624 12850 57652 13262
rect 57888 13252 57940 13258
rect 57888 13194 57940 13200
rect 57900 12850 57928 13194
rect 57612 12844 57664 12850
rect 57612 12786 57664 12792
rect 57888 12844 57940 12850
rect 57888 12786 57940 12792
rect 57900 11762 57928 12786
rect 57888 11756 57940 11762
rect 57888 11698 57940 11704
rect 57992 9654 58020 13330
rect 58084 12646 58112 15982
rect 58268 13530 58296 16594
rect 58256 13524 58308 13530
rect 58256 13466 58308 13472
rect 58728 13190 58756 16594
rect 59188 16590 59216 17546
rect 59372 17202 59400 19110
rect 59544 17740 59596 17746
rect 59544 17682 59596 17688
rect 59556 17626 59584 17682
rect 59464 17598 59584 17626
rect 59360 17196 59412 17202
rect 59360 17138 59412 17144
rect 59464 16658 59492 17598
rect 59544 17536 59596 17542
rect 59544 17478 59596 17484
rect 59452 16652 59504 16658
rect 59452 16594 59504 16600
rect 59176 16584 59228 16590
rect 59004 16546 59176 16574
rect 59004 16454 59032 16546
rect 59176 16526 59228 16532
rect 58992 16448 59044 16454
rect 58992 16390 59044 16396
rect 59004 15978 59032 16390
rect 58992 15972 59044 15978
rect 58992 15914 59044 15920
rect 59556 14958 59584 17478
rect 59728 16992 59780 16998
rect 59728 16934 59780 16940
rect 59740 15570 59768 16934
rect 60108 16794 60136 19264
rect 60188 19246 60240 19252
rect 60188 19168 60240 19174
rect 60188 19110 60240 19116
rect 60200 17746 60228 19110
rect 60384 18426 60412 117098
rect 61016 116612 61068 116618
rect 61016 116554 61068 116560
rect 61028 19310 61056 116554
rect 62960 116346 62988 117098
rect 65248 116680 65300 116686
rect 65248 116622 65300 116628
rect 62948 116340 63000 116346
rect 62948 116282 63000 116288
rect 65260 19310 65288 116622
rect 61016 19304 61068 19310
rect 61016 19246 61068 19252
rect 65248 19304 65300 19310
rect 65248 19246 65300 19252
rect 60372 18420 60424 18426
rect 60372 18362 60424 18368
rect 60188 17740 60240 17746
rect 60188 17682 60240 17688
rect 60556 17536 60608 17542
rect 60556 17478 60608 17484
rect 60568 17338 60596 17478
rect 60556 17332 60608 17338
rect 60556 17274 60608 17280
rect 60096 16788 60148 16794
rect 60096 16730 60148 16736
rect 59728 15564 59780 15570
rect 59728 15506 59780 15512
rect 59544 14952 59596 14958
rect 59544 14894 59596 14900
rect 59740 14890 59768 15506
rect 59728 14884 59780 14890
rect 59728 14826 59780 14832
rect 60096 14884 60148 14890
rect 60096 14826 60148 14832
rect 60108 14006 60136 14826
rect 60096 14000 60148 14006
rect 60096 13942 60148 13948
rect 59912 13932 59964 13938
rect 59912 13874 59964 13880
rect 59924 13530 59952 13874
rect 60372 13864 60424 13870
rect 60372 13806 60424 13812
rect 59912 13524 59964 13530
rect 59912 13466 59964 13472
rect 60280 13252 60332 13258
rect 60280 13194 60332 13200
rect 58716 13184 58768 13190
rect 58716 13126 58768 13132
rect 60096 13184 60148 13190
rect 60096 13126 60148 13132
rect 58532 12980 58584 12986
rect 58532 12922 58584 12928
rect 58072 12640 58124 12646
rect 58072 12582 58124 12588
rect 58084 12102 58112 12582
rect 58072 12096 58124 12102
rect 58072 12038 58124 12044
rect 57980 9648 58032 9654
rect 57980 9590 58032 9596
rect 57980 9444 58032 9450
rect 57980 9386 58032 9392
rect 57336 6724 57388 6730
rect 57336 6666 57388 6672
rect 57348 6322 57376 6666
rect 57704 6656 57756 6662
rect 57704 6598 57756 6604
rect 57886 6624 57942 6633
rect 56692 6316 56744 6322
rect 56692 6258 56744 6264
rect 57244 6316 57296 6322
rect 57244 6258 57296 6264
rect 57336 6316 57388 6322
rect 57336 6258 57388 6264
rect 56232 6180 56284 6186
rect 56232 6122 56284 6128
rect 56048 5568 56100 5574
rect 56048 5510 56100 5516
rect 56060 2514 56088 5510
rect 56244 4214 56272 6122
rect 56704 5914 56732 6258
rect 57060 6248 57112 6254
rect 57060 6190 57112 6196
rect 56692 5908 56744 5914
rect 56692 5850 56744 5856
rect 56232 4208 56284 4214
rect 56232 4150 56284 4156
rect 56968 4072 57020 4078
rect 56968 4014 57020 4020
rect 56324 3596 56376 3602
rect 56324 3538 56376 3544
rect 56048 2508 56100 2514
rect 56048 2450 56100 2456
rect 55956 2304 56008 2310
rect 55956 2246 56008 2252
rect 55968 800 55996 2246
rect 56336 800 56364 3538
rect 56692 2984 56744 2990
rect 56692 2926 56744 2932
rect 56704 800 56732 2926
rect 55772 264 55824 270
rect 55772 206 55824 212
rect 55954 0 56010 800
rect 56322 0 56378 800
rect 56690 0 56746 800
rect 56980 542 57008 4014
rect 57072 2774 57100 6190
rect 57612 5704 57664 5710
rect 57612 5646 57664 5652
rect 57428 3596 57480 3602
rect 57428 3538 57480 3544
rect 57072 2746 57192 2774
rect 57060 2304 57112 2310
rect 57060 2246 57112 2252
rect 57072 800 57100 2246
rect 56968 536 57020 542
rect 56968 478 57020 484
rect 57058 0 57114 800
rect 57164 746 57192 2746
rect 57440 800 57468 3538
rect 57624 1834 57652 5646
rect 57716 2514 57744 6598
rect 57886 6559 57942 6568
rect 57900 6186 57928 6559
rect 57992 6458 58020 9386
rect 58084 8022 58112 12038
rect 58072 8016 58124 8022
rect 58072 7958 58124 7964
rect 58348 6792 58400 6798
rect 58070 6760 58126 6769
rect 58348 6734 58400 6740
rect 58070 6695 58126 6704
rect 58084 6662 58112 6695
rect 58072 6656 58124 6662
rect 58072 6598 58124 6604
rect 57980 6452 58032 6458
rect 57980 6394 58032 6400
rect 57888 6180 57940 6186
rect 57888 6122 57940 6128
rect 57796 2984 57848 2990
rect 57796 2926 57848 2932
rect 57704 2508 57756 2514
rect 57704 2450 57756 2456
rect 57612 1828 57664 1834
rect 57612 1770 57664 1776
rect 57808 800 57836 2926
rect 58084 814 58112 6598
rect 58360 6497 58388 6734
rect 58346 6488 58402 6497
rect 58346 6423 58402 6432
rect 58164 6248 58216 6254
rect 58164 6190 58216 6196
rect 58176 5642 58204 6190
rect 58544 5914 58572 12922
rect 59820 12776 59872 12782
rect 59820 12718 59872 12724
rect 59544 11688 59596 11694
rect 59544 11630 59596 11636
rect 59556 9586 59584 11630
rect 59832 9654 59860 12718
rect 60108 12434 60136 13126
rect 60016 12406 60136 12434
rect 59820 9648 59872 9654
rect 59820 9590 59872 9596
rect 59544 9580 59596 9586
rect 59544 9522 59596 9528
rect 59544 9036 59596 9042
rect 59544 8978 59596 8984
rect 59452 8016 59504 8022
rect 59452 7958 59504 7964
rect 59268 7540 59320 7546
rect 59268 7482 59320 7488
rect 59176 6860 59228 6866
rect 59176 6802 59228 6808
rect 58716 6792 58768 6798
rect 59188 6769 59216 6802
rect 58716 6734 58768 6740
rect 59174 6760 59230 6769
rect 58728 6361 58756 6734
rect 59174 6695 59230 6704
rect 58714 6352 58770 6361
rect 59280 6322 59308 7482
rect 59360 6724 59412 6730
rect 59360 6666 59412 6672
rect 58714 6287 58770 6296
rect 59268 6316 59320 6322
rect 58532 5908 58584 5914
rect 58532 5850 58584 5856
rect 58544 5778 58572 5850
rect 58728 5778 58756 6287
rect 59268 6258 59320 6264
rect 59372 6254 59400 6666
rect 59360 6248 59412 6254
rect 59360 6190 59412 6196
rect 59268 6180 59320 6186
rect 59268 6122 59320 6128
rect 59280 5846 59308 6122
rect 59268 5840 59320 5846
rect 59268 5782 59320 5788
rect 59464 5778 59492 7958
rect 59556 5914 59584 8978
rect 59912 7472 59964 7478
rect 59912 7414 59964 7420
rect 59924 6934 59952 7414
rect 59912 6928 59964 6934
rect 59912 6870 59964 6876
rect 60016 6866 60044 12406
rect 60292 11558 60320 13194
rect 60384 12442 60412 13806
rect 60832 13728 60884 13734
rect 61028 13716 61056 19246
rect 61108 19168 61160 19174
rect 61108 19110 61160 19116
rect 61120 17814 61148 19110
rect 61108 17808 61160 17814
rect 61108 17750 61160 17756
rect 63592 17264 63644 17270
rect 63592 17206 63644 17212
rect 63500 17128 63552 17134
rect 63500 17070 63552 17076
rect 63512 16046 63540 17070
rect 63604 16046 63632 17206
rect 63500 16040 63552 16046
rect 63500 15982 63552 15988
rect 63592 16040 63644 16046
rect 65260 15994 65288 19246
rect 65536 18698 65564 117098
rect 66076 116748 66128 116754
rect 66076 116690 66128 116696
rect 65660 116444 65956 116464
rect 65716 116442 65740 116444
rect 65796 116442 65820 116444
rect 65876 116442 65900 116444
rect 65738 116390 65740 116442
rect 65802 116390 65814 116442
rect 65876 116390 65878 116442
rect 65716 116388 65740 116390
rect 65796 116388 65820 116390
rect 65876 116388 65900 116390
rect 65660 116368 65956 116388
rect 65660 115356 65956 115376
rect 65716 115354 65740 115356
rect 65796 115354 65820 115356
rect 65876 115354 65900 115356
rect 65738 115302 65740 115354
rect 65802 115302 65814 115354
rect 65876 115302 65878 115354
rect 65716 115300 65740 115302
rect 65796 115300 65820 115302
rect 65876 115300 65900 115302
rect 65660 115280 65956 115300
rect 65660 114268 65956 114288
rect 65716 114266 65740 114268
rect 65796 114266 65820 114268
rect 65876 114266 65900 114268
rect 65738 114214 65740 114266
rect 65802 114214 65814 114266
rect 65876 114214 65878 114266
rect 65716 114212 65740 114214
rect 65796 114212 65820 114214
rect 65876 114212 65900 114214
rect 65660 114192 65956 114212
rect 65660 113180 65956 113200
rect 65716 113178 65740 113180
rect 65796 113178 65820 113180
rect 65876 113178 65900 113180
rect 65738 113126 65740 113178
rect 65802 113126 65814 113178
rect 65876 113126 65878 113178
rect 65716 113124 65740 113126
rect 65796 113124 65820 113126
rect 65876 113124 65900 113126
rect 65660 113104 65956 113124
rect 65660 112092 65956 112112
rect 65716 112090 65740 112092
rect 65796 112090 65820 112092
rect 65876 112090 65900 112092
rect 65738 112038 65740 112090
rect 65802 112038 65814 112090
rect 65876 112038 65878 112090
rect 65716 112036 65740 112038
rect 65796 112036 65820 112038
rect 65876 112036 65900 112038
rect 65660 112016 65956 112036
rect 65660 111004 65956 111024
rect 65716 111002 65740 111004
rect 65796 111002 65820 111004
rect 65876 111002 65900 111004
rect 65738 110950 65740 111002
rect 65802 110950 65814 111002
rect 65876 110950 65878 111002
rect 65716 110948 65740 110950
rect 65796 110948 65820 110950
rect 65876 110948 65900 110950
rect 65660 110928 65956 110948
rect 65660 109916 65956 109936
rect 65716 109914 65740 109916
rect 65796 109914 65820 109916
rect 65876 109914 65900 109916
rect 65738 109862 65740 109914
rect 65802 109862 65814 109914
rect 65876 109862 65878 109914
rect 65716 109860 65740 109862
rect 65796 109860 65820 109862
rect 65876 109860 65900 109862
rect 65660 109840 65956 109860
rect 65660 108828 65956 108848
rect 65716 108826 65740 108828
rect 65796 108826 65820 108828
rect 65876 108826 65900 108828
rect 65738 108774 65740 108826
rect 65802 108774 65814 108826
rect 65876 108774 65878 108826
rect 65716 108772 65740 108774
rect 65796 108772 65820 108774
rect 65876 108772 65900 108774
rect 65660 108752 65956 108772
rect 65660 107740 65956 107760
rect 65716 107738 65740 107740
rect 65796 107738 65820 107740
rect 65876 107738 65900 107740
rect 65738 107686 65740 107738
rect 65802 107686 65814 107738
rect 65876 107686 65878 107738
rect 65716 107684 65740 107686
rect 65796 107684 65820 107686
rect 65876 107684 65900 107686
rect 65660 107664 65956 107684
rect 65660 106652 65956 106672
rect 65716 106650 65740 106652
rect 65796 106650 65820 106652
rect 65876 106650 65900 106652
rect 65738 106598 65740 106650
rect 65802 106598 65814 106650
rect 65876 106598 65878 106650
rect 65716 106596 65740 106598
rect 65796 106596 65820 106598
rect 65876 106596 65900 106598
rect 65660 106576 65956 106596
rect 65660 105564 65956 105584
rect 65716 105562 65740 105564
rect 65796 105562 65820 105564
rect 65876 105562 65900 105564
rect 65738 105510 65740 105562
rect 65802 105510 65814 105562
rect 65876 105510 65878 105562
rect 65716 105508 65740 105510
rect 65796 105508 65820 105510
rect 65876 105508 65900 105510
rect 65660 105488 65956 105508
rect 65660 104476 65956 104496
rect 65716 104474 65740 104476
rect 65796 104474 65820 104476
rect 65876 104474 65900 104476
rect 65738 104422 65740 104474
rect 65802 104422 65814 104474
rect 65876 104422 65878 104474
rect 65716 104420 65740 104422
rect 65796 104420 65820 104422
rect 65876 104420 65900 104422
rect 65660 104400 65956 104420
rect 65660 103388 65956 103408
rect 65716 103386 65740 103388
rect 65796 103386 65820 103388
rect 65876 103386 65900 103388
rect 65738 103334 65740 103386
rect 65802 103334 65814 103386
rect 65876 103334 65878 103386
rect 65716 103332 65740 103334
rect 65796 103332 65820 103334
rect 65876 103332 65900 103334
rect 65660 103312 65956 103332
rect 65660 102300 65956 102320
rect 65716 102298 65740 102300
rect 65796 102298 65820 102300
rect 65876 102298 65900 102300
rect 65738 102246 65740 102298
rect 65802 102246 65814 102298
rect 65876 102246 65878 102298
rect 65716 102244 65740 102246
rect 65796 102244 65820 102246
rect 65876 102244 65900 102246
rect 65660 102224 65956 102244
rect 65660 101212 65956 101232
rect 65716 101210 65740 101212
rect 65796 101210 65820 101212
rect 65876 101210 65900 101212
rect 65738 101158 65740 101210
rect 65802 101158 65814 101210
rect 65876 101158 65878 101210
rect 65716 101156 65740 101158
rect 65796 101156 65820 101158
rect 65876 101156 65900 101158
rect 65660 101136 65956 101156
rect 65660 100124 65956 100144
rect 65716 100122 65740 100124
rect 65796 100122 65820 100124
rect 65876 100122 65900 100124
rect 65738 100070 65740 100122
rect 65802 100070 65814 100122
rect 65876 100070 65878 100122
rect 65716 100068 65740 100070
rect 65796 100068 65820 100070
rect 65876 100068 65900 100070
rect 65660 100048 65956 100068
rect 65660 99036 65956 99056
rect 65716 99034 65740 99036
rect 65796 99034 65820 99036
rect 65876 99034 65900 99036
rect 65738 98982 65740 99034
rect 65802 98982 65814 99034
rect 65876 98982 65878 99034
rect 65716 98980 65740 98982
rect 65796 98980 65820 98982
rect 65876 98980 65900 98982
rect 65660 98960 65956 98980
rect 65660 97948 65956 97968
rect 65716 97946 65740 97948
rect 65796 97946 65820 97948
rect 65876 97946 65900 97948
rect 65738 97894 65740 97946
rect 65802 97894 65814 97946
rect 65876 97894 65878 97946
rect 65716 97892 65740 97894
rect 65796 97892 65820 97894
rect 65876 97892 65900 97894
rect 65660 97872 65956 97892
rect 65660 96860 65956 96880
rect 65716 96858 65740 96860
rect 65796 96858 65820 96860
rect 65876 96858 65900 96860
rect 65738 96806 65740 96858
rect 65802 96806 65814 96858
rect 65876 96806 65878 96858
rect 65716 96804 65740 96806
rect 65796 96804 65820 96806
rect 65876 96804 65900 96806
rect 65660 96784 65956 96804
rect 65660 95772 65956 95792
rect 65716 95770 65740 95772
rect 65796 95770 65820 95772
rect 65876 95770 65900 95772
rect 65738 95718 65740 95770
rect 65802 95718 65814 95770
rect 65876 95718 65878 95770
rect 65716 95716 65740 95718
rect 65796 95716 65820 95718
rect 65876 95716 65900 95718
rect 65660 95696 65956 95716
rect 65660 94684 65956 94704
rect 65716 94682 65740 94684
rect 65796 94682 65820 94684
rect 65876 94682 65900 94684
rect 65738 94630 65740 94682
rect 65802 94630 65814 94682
rect 65876 94630 65878 94682
rect 65716 94628 65740 94630
rect 65796 94628 65820 94630
rect 65876 94628 65900 94630
rect 65660 94608 65956 94628
rect 65660 93596 65956 93616
rect 65716 93594 65740 93596
rect 65796 93594 65820 93596
rect 65876 93594 65900 93596
rect 65738 93542 65740 93594
rect 65802 93542 65814 93594
rect 65876 93542 65878 93594
rect 65716 93540 65740 93542
rect 65796 93540 65820 93542
rect 65876 93540 65900 93542
rect 65660 93520 65956 93540
rect 65660 92508 65956 92528
rect 65716 92506 65740 92508
rect 65796 92506 65820 92508
rect 65876 92506 65900 92508
rect 65738 92454 65740 92506
rect 65802 92454 65814 92506
rect 65876 92454 65878 92506
rect 65716 92452 65740 92454
rect 65796 92452 65820 92454
rect 65876 92452 65900 92454
rect 65660 92432 65956 92452
rect 65660 91420 65956 91440
rect 65716 91418 65740 91420
rect 65796 91418 65820 91420
rect 65876 91418 65900 91420
rect 65738 91366 65740 91418
rect 65802 91366 65814 91418
rect 65876 91366 65878 91418
rect 65716 91364 65740 91366
rect 65796 91364 65820 91366
rect 65876 91364 65900 91366
rect 65660 91344 65956 91364
rect 65660 90332 65956 90352
rect 65716 90330 65740 90332
rect 65796 90330 65820 90332
rect 65876 90330 65900 90332
rect 65738 90278 65740 90330
rect 65802 90278 65814 90330
rect 65876 90278 65878 90330
rect 65716 90276 65740 90278
rect 65796 90276 65820 90278
rect 65876 90276 65900 90278
rect 65660 90256 65956 90276
rect 65660 89244 65956 89264
rect 65716 89242 65740 89244
rect 65796 89242 65820 89244
rect 65876 89242 65900 89244
rect 65738 89190 65740 89242
rect 65802 89190 65814 89242
rect 65876 89190 65878 89242
rect 65716 89188 65740 89190
rect 65796 89188 65820 89190
rect 65876 89188 65900 89190
rect 65660 89168 65956 89188
rect 65660 88156 65956 88176
rect 65716 88154 65740 88156
rect 65796 88154 65820 88156
rect 65876 88154 65900 88156
rect 65738 88102 65740 88154
rect 65802 88102 65814 88154
rect 65876 88102 65878 88154
rect 65716 88100 65740 88102
rect 65796 88100 65820 88102
rect 65876 88100 65900 88102
rect 65660 88080 65956 88100
rect 65660 87068 65956 87088
rect 65716 87066 65740 87068
rect 65796 87066 65820 87068
rect 65876 87066 65900 87068
rect 65738 87014 65740 87066
rect 65802 87014 65814 87066
rect 65876 87014 65878 87066
rect 65716 87012 65740 87014
rect 65796 87012 65820 87014
rect 65876 87012 65900 87014
rect 65660 86992 65956 87012
rect 65660 85980 65956 86000
rect 65716 85978 65740 85980
rect 65796 85978 65820 85980
rect 65876 85978 65900 85980
rect 65738 85926 65740 85978
rect 65802 85926 65814 85978
rect 65876 85926 65878 85978
rect 65716 85924 65740 85926
rect 65796 85924 65820 85926
rect 65876 85924 65900 85926
rect 65660 85904 65956 85924
rect 65660 84892 65956 84912
rect 65716 84890 65740 84892
rect 65796 84890 65820 84892
rect 65876 84890 65900 84892
rect 65738 84838 65740 84890
rect 65802 84838 65814 84890
rect 65876 84838 65878 84890
rect 65716 84836 65740 84838
rect 65796 84836 65820 84838
rect 65876 84836 65900 84838
rect 65660 84816 65956 84836
rect 65660 83804 65956 83824
rect 65716 83802 65740 83804
rect 65796 83802 65820 83804
rect 65876 83802 65900 83804
rect 65738 83750 65740 83802
rect 65802 83750 65814 83802
rect 65876 83750 65878 83802
rect 65716 83748 65740 83750
rect 65796 83748 65820 83750
rect 65876 83748 65900 83750
rect 65660 83728 65956 83748
rect 65660 82716 65956 82736
rect 65716 82714 65740 82716
rect 65796 82714 65820 82716
rect 65876 82714 65900 82716
rect 65738 82662 65740 82714
rect 65802 82662 65814 82714
rect 65876 82662 65878 82714
rect 65716 82660 65740 82662
rect 65796 82660 65820 82662
rect 65876 82660 65900 82662
rect 65660 82640 65956 82660
rect 65660 81628 65956 81648
rect 65716 81626 65740 81628
rect 65796 81626 65820 81628
rect 65876 81626 65900 81628
rect 65738 81574 65740 81626
rect 65802 81574 65814 81626
rect 65876 81574 65878 81626
rect 65716 81572 65740 81574
rect 65796 81572 65820 81574
rect 65876 81572 65900 81574
rect 65660 81552 65956 81572
rect 65660 80540 65956 80560
rect 65716 80538 65740 80540
rect 65796 80538 65820 80540
rect 65876 80538 65900 80540
rect 65738 80486 65740 80538
rect 65802 80486 65814 80538
rect 65876 80486 65878 80538
rect 65716 80484 65740 80486
rect 65796 80484 65820 80486
rect 65876 80484 65900 80486
rect 65660 80464 65956 80484
rect 65660 79452 65956 79472
rect 65716 79450 65740 79452
rect 65796 79450 65820 79452
rect 65876 79450 65900 79452
rect 65738 79398 65740 79450
rect 65802 79398 65814 79450
rect 65876 79398 65878 79450
rect 65716 79396 65740 79398
rect 65796 79396 65820 79398
rect 65876 79396 65900 79398
rect 65660 79376 65956 79396
rect 65660 78364 65956 78384
rect 65716 78362 65740 78364
rect 65796 78362 65820 78364
rect 65876 78362 65900 78364
rect 65738 78310 65740 78362
rect 65802 78310 65814 78362
rect 65876 78310 65878 78362
rect 65716 78308 65740 78310
rect 65796 78308 65820 78310
rect 65876 78308 65900 78310
rect 65660 78288 65956 78308
rect 65660 77276 65956 77296
rect 65716 77274 65740 77276
rect 65796 77274 65820 77276
rect 65876 77274 65900 77276
rect 65738 77222 65740 77274
rect 65802 77222 65814 77274
rect 65876 77222 65878 77274
rect 65716 77220 65740 77222
rect 65796 77220 65820 77222
rect 65876 77220 65900 77222
rect 65660 77200 65956 77220
rect 65660 76188 65956 76208
rect 65716 76186 65740 76188
rect 65796 76186 65820 76188
rect 65876 76186 65900 76188
rect 65738 76134 65740 76186
rect 65802 76134 65814 76186
rect 65876 76134 65878 76186
rect 65716 76132 65740 76134
rect 65796 76132 65820 76134
rect 65876 76132 65900 76134
rect 65660 76112 65956 76132
rect 65660 75100 65956 75120
rect 65716 75098 65740 75100
rect 65796 75098 65820 75100
rect 65876 75098 65900 75100
rect 65738 75046 65740 75098
rect 65802 75046 65814 75098
rect 65876 75046 65878 75098
rect 65716 75044 65740 75046
rect 65796 75044 65820 75046
rect 65876 75044 65900 75046
rect 65660 75024 65956 75044
rect 65660 74012 65956 74032
rect 65716 74010 65740 74012
rect 65796 74010 65820 74012
rect 65876 74010 65900 74012
rect 65738 73958 65740 74010
rect 65802 73958 65814 74010
rect 65876 73958 65878 74010
rect 65716 73956 65740 73958
rect 65796 73956 65820 73958
rect 65876 73956 65900 73958
rect 65660 73936 65956 73956
rect 65660 72924 65956 72944
rect 65716 72922 65740 72924
rect 65796 72922 65820 72924
rect 65876 72922 65900 72924
rect 65738 72870 65740 72922
rect 65802 72870 65814 72922
rect 65876 72870 65878 72922
rect 65716 72868 65740 72870
rect 65796 72868 65820 72870
rect 65876 72868 65900 72870
rect 65660 72848 65956 72868
rect 65660 71836 65956 71856
rect 65716 71834 65740 71836
rect 65796 71834 65820 71836
rect 65876 71834 65900 71836
rect 65738 71782 65740 71834
rect 65802 71782 65814 71834
rect 65876 71782 65878 71834
rect 65716 71780 65740 71782
rect 65796 71780 65820 71782
rect 65876 71780 65900 71782
rect 65660 71760 65956 71780
rect 65660 70748 65956 70768
rect 65716 70746 65740 70748
rect 65796 70746 65820 70748
rect 65876 70746 65900 70748
rect 65738 70694 65740 70746
rect 65802 70694 65814 70746
rect 65876 70694 65878 70746
rect 65716 70692 65740 70694
rect 65796 70692 65820 70694
rect 65876 70692 65900 70694
rect 65660 70672 65956 70692
rect 65660 69660 65956 69680
rect 65716 69658 65740 69660
rect 65796 69658 65820 69660
rect 65876 69658 65900 69660
rect 65738 69606 65740 69658
rect 65802 69606 65814 69658
rect 65876 69606 65878 69658
rect 65716 69604 65740 69606
rect 65796 69604 65820 69606
rect 65876 69604 65900 69606
rect 65660 69584 65956 69604
rect 65660 68572 65956 68592
rect 65716 68570 65740 68572
rect 65796 68570 65820 68572
rect 65876 68570 65900 68572
rect 65738 68518 65740 68570
rect 65802 68518 65814 68570
rect 65876 68518 65878 68570
rect 65716 68516 65740 68518
rect 65796 68516 65820 68518
rect 65876 68516 65900 68518
rect 65660 68496 65956 68516
rect 65660 67484 65956 67504
rect 65716 67482 65740 67484
rect 65796 67482 65820 67484
rect 65876 67482 65900 67484
rect 65738 67430 65740 67482
rect 65802 67430 65814 67482
rect 65876 67430 65878 67482
rect 65716 67428 65740 67430
rect 65796 67428 65820 67430
rect 65876 67428 65900 67430
rect 65660 67408 65956 67428
rect 65660 66396 65956 66416
rect 65716 66394 65740 66396
rect 65796 66394 65820 66396
rect 65876 66394 65900 66396
rect 65738 66342 65740 66394
rect 65802 66342 65814 66394
rect 65876 66342 65878 66394
rect 65716 66340 65740 66342
rect 65796 66340 65820 66342
rect 65876 66340 65900 66342
rect 65660 66320 65956 66340
rect 65660 65308 65956 65328
rect 65716 65306 65740 65308
rect 65796 65306 65820 65308
rect 65876 65306 65900 65308
rect 65738 65254 65740 65306
rect 65802 65254 65814 65306
rect 65876 65254 65878 65306
rect 65716 65252 65740 65254
rect 65796 65252 65820 65254
rect 65876 65252 65900 65254
rect 65660 65232 65956 65252
rect 65660 64220 65956 64240
rect 65716 64218 65740 64220
rect 65796 64218 65820 64220
rect 65876 64218 65900 64220
rect 65738 64166 65740 64218
rect 65802 64166 65814 64218
rect 65876 64166 65878 64218
rect 65716 64164 65740 64166
rect 65796 64164 65820 64166
rect 65876 64164 65900 64166
rect 65660 64144 65956 64164
rect 65660 63132 65956 63152
rect 65716 63130 65740 63132
rect 65796 63130 65820 63132
rect 65876 63130 65900 63132
rect 65738 63078 65740 63130
rect 65802 63078 65814 63130
rect 65876 63078 65878 63130
rect 65716 63076 65740 63078
rect 65796 63076 65820 63078
rect 65876 63076 65900 63078
rect 65660 63056 65956 63076
rect 65660 62044 65956 62064
rect 65716 62042 65740 62044
rect 65796 62042 65820 62044
rect 65876 62042 65900 62044
rect 65738 61990 65740 62042
rect 65802 61990 65814 62042
rect 65876 61990 65878 62042
rect 65716 61988 65740 61990
rect 65796 61988 65820 61990
rect 65876 61988 65900 61990
rect 65660 61968 65956 61988
rect 65660 60956 65956 60976
rect 65716 60954 65740 60956
rect 65796 60954 65820 60956
rect 65876 60954 65900 60956
rect 65738 60902 65740 60954
rect 65802 60902 65814 60954
rect 65876 60902 65878 60954
rect 65716 60900 65740 60902
rect 65796 60900 65820 60902
rect 65876 60900 65900 60902
rect 65660 60880 65956 60900
rect 65660 59868 65956 59888
rect 65716 59866 65740 59868
rect 65796 59866 65820 59868
rect 65876 59866 65900 59868
rect 65738 59814 65740 59866
rect 65802 59814 65814 59866
rect 65876 59814 65878 59866
rect 65716 59812 65740 59814
rect 65796 59812 65820 59814
rect 65876 59812 65900 59814
rect 65660 59792 65956 59812
rect 65660 58780 65956 58800
rect 65716 58778 65740 58780
rect 65796 58778 65820 58780
rect 65876 58778 65900 58780
rect 65738 58726 65740 58778
rect 65802 58726 65814 58778
rect 65876 58726 65878 58778
rect 65716 58724 65740 58726
rect 65796 58724 65820 58726
rect 65876 58724 65900 58726
rect 65660 58704 65956 58724
rect 65660 57692 65956 57712
rect 65716 57690 65740 57692
rect 65796 57690 65820 57692
rect 65876 57690 65900 57692
rect 65738 57638 65740 57690
rect 65802 57638 65814 57690
rect 65876 57638 65878 57690
rect 65716 57636 65740 57638
rect 65796 57636 65820 57638
rect 65876 57636 65900 57638
rect 65660 57616 65956 57636
rect 65660 56604 65956 56624
rect 65716 56602 65740 56604
rect 65796 56602 65820 56604
rect 65876 56602 65900 56604
rect 65738 56550 65740 56602
rect 65802 56550 65814 56602
rect 65876 56550 65878 56602
rect 65716 56548 65740 56550
rect 65796 56548 65820 56550
rect 65876 56548 65900 56550
rect 65660 56528 65956 56548
rect 65660 55516 65956 55536
rect 65716 55514 65740 55516
rect 65796 55514 65820 55516
rect 65876 55514 65900 55516
rect 65738 55462 65740 55514
rect 65802 55462 65814 55514
rect 65876 55462 65878 55514
rect 65716 55460 65740 55462
rect 65796 55460 65820 55462
rect 65876 55460 65900 55462
rect 65660 55440 65956 55460
rect 65660 54428 65956 54448
rect 65716 54426 65740 54428
rect 65796 54426 65820 54428
rect 65876 54426 65900 54428
rect 65738 54374 65740 54426
rect 65802 54374 65814 54426
rect 65876 54374 65878 54426
rect 65716 54372 65740 54374
rect 65796 54372 65820 54374
rect 65876 54372 65900 54374
rect 65660 54352 65956 54372
rect 65660 53340 65956 53360
rect 65716 53338 65740 53340
rect 65796 53338 65820 53340
rect 65876 53338 65900 53340
rect 65738 53286 65740 53338
rect 65802 53286 65814 53338
rect 65876 53286 65878 53338
rect 65716 53284 65740 53286
rect 65796 53284 65820 53286
rect 65876 53284 65900 53286
rect 65660 53264 65956 53284
rect 65660 52252 65956 52272
rect 65716 52250 65740 52252
rect 65796 52250 65820 52252
rect 65876 52250 65900 52252
rect 65738 52198 65740 52250
rect 65802 52198 65814 52250
rect 65876 52198 65878 52250
rect 65716 52196 65740 52198
rect 65796 52196 65820 52198
rect 65876 52196 65900 52198
rect 65660 52176 65956 52196
rect 65660 51164 65956 51184
rect 65716 51162 65740 51164
rect 65796 51162 65820 51164
rect 65876 51162 65900 51164
rect 65738 51110 65740 51162
rect 65802 51110 65814 51162
rect 65876 51110 65878 51162
rect 65716 51108 65740 51110
rect 65796 51108 65820 51110
rect 65876 51108 65900 51110
rect 65660 51088 65956 51108
rect 65660 50076 65956 50096
rect 65716 50074 65740 50076
rect 65796 50074 65820 50076
rect 65876 50074 65900 50076
rect 65738 50022 65740 50074
rect 65802 50022 65814 50074
rect 65876 50022 65878 50074
rect 65716 50020 65740 50022
rect 65796 50020 65820 50022
rect 65876 50020 65900 50022
rect 65660 50000 65956 50020
rect 65660 48988 65956 49008
rect 65716 48986 65740 48988
rect 65796 48986 65820 48988
rect 65876 48986 65900 48988
rect 65738 48934 65740 48986
rect 65802 48934 65814 48986
rect 65876 48934 65878 48986
rect 65716 48932 65740 48934
rect 65796 48932 65820 48934
rect 65876 48932 65900 48934
rect 65660 48912 65956 48932
rect 65660 47900 65956 47920
rect 65716 47898 65740 47900
rect 65796 47898 65820 47900
rect 65876 47898 65900 47900
rect 65738 47846 65740 47898
rect 65802 47846 65814 47898
rect 65876 47846 65878 47898
rect 65716 47844 65740 47846
rect 65796 47844 65820 47846
rect 65876 47844 65900 47846
rect 65660 47824 65956 47844
rect 65660 46812 65956 46832
rect 65716 46810 65740 46812
rect 65796 46810 65820 46812
rect 65876 46810 65900 46812
rect 65738 46758 65740 46810
rect 65802 46758 65814 46810
rect 65876 46758 65878 46810
rect 65716 46756 65740 46758
rect 65796 46756 65820 46758
rect 65876 46756 65900 46758
rect 65660 46736 65956 46756
rect 65660 45724 65956 45744
rect 65716 45722 65740 45724
rect 65796 45722 65820 45724
rect 65876 45722 65900 45724
rect 65738 45670 65740 45722
rect 65802 45670 65814 45722
rect 65876 45670 65878 45722
rect 65716 45668 65740 45670
rect 65796 45668 65820 45670
rect 65876 45668 65900 45670
rect 65660 45648 65956 45668
rect 65660 44636 65956 44656
rect 65716 44634 65740 44636
rect 65796 44634 65820 44636
rect 65876 44634 65900 44636
rect 65738 44582 65740 44634
rect 65802 44582 65814 44634
rect 65876 44582 65878 44634
rect 65716 44580 65740 44582
rect 65796 44580 65820 44582
rect 65876 44580 65900 44582
rect 65660 44560 65956 44580
rect 65660 43548 65956 43568
rect 65716 43546 65740 43548
rect 65796 43546 65820 43548
rect 65876 43546 65900 43548
rect 65738 43494 65740 43546
rect 65802 43494 65814 43546
rect 65876 43494 65878 43546
rect 65716 43492 65740 43494
rect 65796 43492 65820 43494
rect 65876 43492 65900 43494
rect 65660 43472 65956 43492
rect 65660 42460 65956 42480
rect 65716 42458 65740 42460
rect 65796 42458 65820 42460
rect 65876 42458 65900 42460
rect 65738 42406 65740 42458
rect 65802 42406 65814 42458
rect 65876 42406 65878 42458
rect 65716 42404 65740 42406
rect 65796 42404 65820 42406
rect 65876 42404 65900 42406
rect 65660 42384 65956 42404
rect 65660 41372 65956 41392
rect 65716 41370 65740 41372
rect 65796 41370 65820 41372
rect 65876 41370 65900 41372
rect 65738 41318 65740 41370
rect 65802 41318 65814 41370
rect 65876 41318 65878 41370
rect 65716 41316 65740 41318
rect 65796 41316 65820 41318
rect 65876 41316 65900 41318
rect 65660 41296 65956 41316
rect 65660 40284 65956 40304
rect 65716 40282 65740 40284
rect 65796 40282 65820 40284
rect 65876 40282 65900 40284
rect 65738 40230 65740 40282
rect 65802 40230 65814 40282
rect 65876 40230 65878 40282
rect 65716 40228 65740 40230
rect 65796 40228 65820 40230
rect 65876 40228 65900 40230
rect 65660 40208 65956 40228
rect 65660 39196 65956 39216
rect 65716 39194 65740 39196
rect 65796 39194 65820 39196
rect 65876 39194 65900 39196
rect 65738 39142 65740 39194
rect 65802 39142 65814 39194
rect 65876 39142 65878 39194
rect 65716 39140 65740 39142
rect 65796 39140 65820 39142
rect 65876 39140 65900 39142
rect 65660 39120 65956 39140
rect 65660 38108 65956 38128
rect 65716 38106 65740 38108
rect 65796 38106 65820 38108
rect 65876 38106 65900 38108
rect 65738 38054 65740 38106
rect 65802 38054 65814 38106
rect 65876 38054 65878 38106
rect 65716 38052 65740 38054
rect 65796 38052 65820 38054
rect 65876 38052 65900 38054
rect 65660 38032 65956 38052
rect 65660 37020 65956 37040
rect 65716 37018 65740 37020
rect 65796 37018 65820 37020
rect 65876 37018 65900 37020
rect 65738 36966 65740 37018
rect 65802 36966 65814 37018
rect 65876 36966 65878 37018
rect 65716 36964 65740 36966
rect 65796 36964 65820 36966
rect 65876 36964 65900 36966
rect 65660 36944 65956 36964
rect 65660 35932 65956 35952
rect 65716 35930 65740 35932
rect 65796 35930 65820 35932
rect 65876 35930 65900 35932
rect 65738 35878 65740 35930
rect 65802 35878 65814 35930
rect 65876 35878 65878 35930
rect 65716 35876 65740 35878
rect 65796 35876 65820 35878
rect 65876 35876 65900 35878
rect 65660 35856 65956 35876
rect 65660 34844 65956 34864
rect 65716 34842 65740 34844
rect 65796 34842 65820 34844
rect 65876 34842 65900 34844
rect 65738 34790 65740 34842
rect 65802 34790 65814 34842
rect 65876 34790 65878 34842
rect 65716 34788 65740 34790
rect 65796 34788 65820 34790
rect 65876 34788 65900 34790
rect 65660 34768 65956 34788
rect 65660 33756 65956 33776
rect 65716 33754 65740 33756
rect 65796 33754 65820 33756
rect 65876 33754 65900 33756
rect 65738 33702 65740 33754
rect 65802 33702 65814 33754
rect 65876 33702 65878 33754
rect 65716 33700 65740 33702
rect 65796 33700 65820 33702
rect 65876 33700 65900 33702
rect 65660 33680 65956 33700
rect 65660 32668 65956 32688
rect 65716 32666 65740 32668
rect 65796 32666 65820 32668
rect 65876 32666 65900 32668
rect 65738 32614 65740 32666
rect 65802 32614 65814 32666
rect 65876 32614 65878 32666
rect 65716 32612 65740 32614
rect 65796 32612 65820 32614
rect 65876 32612 65900 32614
rect 65660 32592 65956 32612
rect 65660 31580 65956 31600
rect 65716 31578 65740 31580
rect 65796 31578 65820 31580
rect 65876 31578 65900 31580
rect 65738 31526 65740 31578
rect 65802 31526 65814 31578
rect 65876 31526 65878 31578
rect 65716 31524 65740 31526
rect 65796 31524 65820 31526
rect 65876 31524 65900 31526
rect 65660 31504 65956 31524
rect 65660 30492 65956 30512
rect 65716 30490 65740 30492
rect 65796 30490 65820 30492
rect 65876 30490 65900 30492
rect 65738 30438 65740 30490
rect 65802 30438 65814 30490
rect 65876 30438 65878 30490
rect 65716 30436 65740 30438
rect 65796 30436 65820 30438
rect 65876 30436 65900 30438
rect 65660 30416 65956 30436
rect 65660 29404 65956 29424
rect 65716 29402 65740 29404
rect 65796 29402 65820 29404
rect 65876 29402 65900 29404
rect 65738 29350 65740 29402
rect 65802 29350 65814 29402
rect 65876 29350 65878 29402
rect 65716 29348 65740 29350
rect 65796 29348 65820 29350
rect 65876 29348 65900 29350
rect 65660 29328 65956 29348
rect 65660 28316 65956 28336
rect 65716 28314 65740 28316
rect 65796 28314 65820 28316
rect 65876 28314 65900 28316
rect 65738 28262 65740 28314
rect 65802 28262 65814 28314
rect 65876 28262 65878 28314
rect 65716 28260 65740 28262
rect 65796 28260 65820 28262
rect 65876 28260 65900 28262
rect 65660 28240 65956 28260
rect 65660 27228 65956 27248
rect 65716 27226 65740 27228
rect 65796 27226 65820 27228
rect 65876 27226 65900 27228
rect 65738 27174 65740 27226
rect 65802 27174 65814 27226
rect 65876 27174 65878 27226
rect 65716 27172 65740 27174
rect 65796 27172 65820 27174
rect 65876 27172 65900 27174
rect 65660 27152 65956 27172
rect 65660 26140 65956 26160
rect 65716 26138 65740 26140
rect 65796 26138 65820 26140
rect 65876 26138 65900 26140
rect 65738 26086 65740 26138
rect 65802 26086 65814 26138
rect 65876 26086 65878 26138
rect 65716 26084 65740 26086
rect 65796 26084 65820 26086
rect 65876 26084 65900 26086
rect 65660 26064 65956 26084
rect 65660 25052 65956 25072
rect 65716 25050 65740 25052
rect 65796 25050 65820 25052
rect 65876 25050 65900 25052
rect 65738 24998 65740 25050
rect 65802 24998 65814 25050
rect 65876 24998 65878 25050
rect 65716 24996 65740 24998
rect 65796 24996 65820 24998
rect 65876 24996 65900 24998
rect 65660 24976 65956 24996
rect 65660 23964 65956 23984
rect 65716 23962 65740 23964
rect 65796 23962 65820 23964
rect 65876 23962 65900 23964
rect 65738 23910 65740 23962
rect 65802 23910 65814 23962
rect 65876 23910 65878 23962
rect 65716 23908 65740 23910
rect 65796 23908 65820 23910
rect 65876 23908 65900 23910
rect 65660 23888 65956 23908
rect 65660 22876 65956 22896
rect 65716 22874 65740 22876
rect 65796 22874 65820 22876
rect 65876 22874 65900 22876
rect 65738 22822 65740 22874
rect 65802 22822 65814 22874
rect 65876 22822 65878 22874
rect 65716 22820 65740 22822
rect 65796 22820 65820 22822
rect 65876 22820 65900 22822
rect 65660 22800 65956 22820
rect 65660 21788 65956 21808
rect 65716 21786 65740 21788
rect 65796 21786 65820 21788
rect 65876 21786 65900 21788
rect 65738 21734 65740 21786
rect 65802 21734 65814 21786
rect 65876 21734 65878 21786
rect 65716 21732 65740 21734
rect 65796 21732 65820 21734
rect 65876 21732 65900 21734
rect 65660 21712 65956 21732
rect 65660 20700 65956 20720
rect 65716 20698 65740 20700
rect 65796 20698 65820 20700
rect 65876 20698 65900 20700
rect 65738 20646 65740 20698
rect 65802 20646 65814 20698
rect 65876 20646 65878 20698
rect 65716 20644 65740 20646
rect 65796 20644 65820 20646
rect 65876 20644 65900 20646
rect 65660 20624 65956 20644
rect 65660 19612 65956 19632
rect 65716 19610 65740 19612
rect 65796 19610 65820 19612
rect 65876 19610 65900 19612
rect 65738 19558 65740 19610
rect 65802 19558 65814 19610
rect 65876 19558 65878 19610
rect 65716 19556 65740 19558
rect 65796 19556 65820 19558
rect 65876 19556 65900 19558
rect 65660 19536 65956 19556
rect 65984 19168 66036 19174
rect 65984 19110 66036 19116
rect 65524 18692 65576 18698
rect 65524 18634 65576 18640
rect 65660 18524 65956 18544
rect 65716 18522 65740 18524
rect 65796 18522 65820 18524
rect 65876 18522 65900 18524
rect 65738 18470 65740 18522
rect 65802 18470 65814 18522
rect 65876 18470 65878 18522
rect 65716 18468 65740 18470
rect 65796 18468 65820 18470
rect 65876 18468 65900 18470
rect 65660 18448 65956 18468
rect 65660 17436 65956 17456
rect 65716 17434 65740 17436
rect 65796 17434 65820 17436
rect 65876 17434 65900 17436
rect 65738 17382 65740 17434
rect 65802 17382 65814 17434
rect 65876 17382 65878 17434
rect 65716 17380 65740 17382
rect 65796 17380 65820 17382
rect 65876 17380 65900 17382
rect 65660 17360 65956 17380
rect 65996 17270 66024 19110
rect 66088 18834 66116 116690
rect 67652 116278 67680 117098
rect 69572 117088 69624 117094
rect 69572 117030 69624 117036
rect 68468 116884 68520 116890
rect 68468 116826 68520 116832
rect 67824 116816 67876 116822
rect 67824 116758 67876 116764
rect 67640 116272 67692 116278
rect 67640 116214 67692 116220
rect 67836 18834 67864 116758
rect 68480 18834 68508 116826
rect 69584 116074 69612 117030
rect 69572 116068 69624 116074
rect 69572 116010 69624 116016
rect 68652 19168 68704 19174
rect 68652 19110 68704 19116
rect 66076 18828 66128 18834
rect 66076 18770 66128 18776
rect 67824 18828 67876 18834
rect 67824 18770 67876 18776
rect 68468 18828 68520 18834
rect 68468 18770 68520 18776
rect 65984 17264 66036 17270
rect 65984 17206 66036 17212
rect 65524 16652 65576 16658
rect 65524 16594 65576 16600
rect 63592 15982 63644 15988
rect 63512 15570 63540 15982
rect 63604 15706 63632 15982
rect 65168 15966 65288 15994
rect 65340 16040 65392 16046
rect 65340 15982 65392 15988
rect 64052 15904 64104 15910
rect 64052 15846 64104 15852
rect 63592 15700 63644 15706
rect 63592 15642 63644 15648
rect 64064 15570 64092 15846
rect 63500 15564 63552 15570
rect 63500 15506 63552 15512
rect 64052 15564 64104 15570
rect 64052 15506 64104 15512
rect 63960 15496 64012 15502
rect 63960 15438 64012 15444
rect 62488 15360 62540 15366
rect 62488 15302 62540 15308
rect 63684 15360 63736 15366
rect 63684 15302 63736 15308
rect 62396 14068 62448 14074
rect 62396 14010 62448 14016
rect 60884 13688 61056 13716
rect 60832 13670 60884 13676
rect 60844 13326 60872 13670
rect 60832 13320 60884 13326
rect 60832 13262 60884 13268
rect 61844 13320 61896 13326
rect 61844 13262 61896 13268
rect 61292 12640 61344 12646
rect 61292 12582 61344 12588
rect 60372 12436 60424 12442
rect 60372 12378 60424 12384
rect 60384 11694 60412 12378
rect 60372 11688 60424 11694
rect 60372 11630 60424 11636
rect 60280 11552 60332 11558
rect 60280 11494 60332 11500
rect 60556 11552 60608 11558
rect 60556 11494 60608 11500
rect 60372 10600 60424 10606
rect 60372 10542 60424 10548
rect 60384 10198 60412 10542
rect 60372 10192 60424 10198
rect 60372 10134 60424 10140
rect 60096 9988 60148 9994
rect 60096 9930 60148 9936
rect 60108 9518 60136 9930
rect 60096 9512 60148 9518
rect 60096 9454 60148 9460
rect 60568 8090 60596 11494
rect 60648 9512 60700 9518
rect 60648 9454 60700 9460
rect 60660 9042 60688 9454
rect 60648 9036 60700 9042
rect 60648 8978 60700 8984
rect 60556 8084 60608 8090
rect 60556 8026 60608 8032
rect 60188 7540 60240 7546
rect 60188 7482 60240 7488
rect 60004 6860 60056 6866
rect 60004 6802 60056 6808
rect 60004 6316 60056 6322
rect 59832 6276 60004 6304
rect 59636 6248 59688 6254
rect 59636 6190 59688 6196
rect 59544 5908 59596 5914
rect 59544 5850 59596 5856
rect 58532 5772 58584 5778
rect 58532 5714 58584 5720
rect 58716 5772 58768 5778
rect 58716 5714 58768 5720
rect 59452 5772 59504 5778
rect 59452 5714 59504 5720
rect 58256 5704 58308 5710
rect 58256 5646 58308 5652
rect 58164 5636 58216 5642
rect 58164 5578 58216 5584
rect 58164 2304 58216 2310
rect 58164 2246 58216 2252
rect 58072 808 58124 814
rect 57152 740 57204 746
rect 57152 682 57204 688
rect 57426 0 57482 800
rect 57794 0 57850 800
rect 58176 800 58204 2246
rect 58268 950 58296 5646
rect 59452 5568 59504 5574
rect 59452 5510 59504 5516
rect 58532 3596 58584 3602
rect 58532 3538 58584 3544
rect 58256 944 58308 950
rect 58256 886 58308 892
rect 58544 800 58572 3538
rect 58900 2984 58952 2990
rect 58900 2926 58952 2932
rect 58912 800 58940 2926
rect 59464 2774 59492 5510
rect 59648 4622 59676 6190
rect 59636 4616 59688 4622
rect 59636 4558 59688 4564
rect 59636 3596 59688 3602
rect 59636 3538 59688 3544
rect 59372 2746 59492 2774
rect 59084 2508 59136 2514
rect 59372 2496 59400 2746
rect 59136 2468 59400 2496
rect 59084 2450 59136 2456
rect 59268 2372 59320 2378
rect 59268 2314 59320 2320
rect 59280 800 59308 2314
rect 59648 800 59676 3538
rect 58072 750 58124 756
rect 58162 0 58218 800
rect 58530 0 58586 800
rect 58898 0 58954 800
rect 59266 0 59322 800
rect 59634 0 59690 800
rect 59832 678 59860 6276
rect 60004 6258 60056 6264
rect 60200 6236 60228 7482
rect 60464 6792 60516 6798
rect 60464 6734 60516 6740
rect 60326 6248 60378 6254
rect 60200 6208 60326 6236
rect 60326 6190 60378 6196
rect 59912 5568 59964 5574
rect 59912 5510 59964 5516
rect 59924 2514 59952 5510
rect 60476 5030 60504 6734
rect 60568 5760 60596 8026
rect 61108 7812 61160 7818
rect 61108 7754 61160 7760
rect 61120 6934 61148 7754
rect 61304 7546 61332 12582
rect 61856 12434 61884 13262
rect 61764 12406 61884 12434
rect 61660 12096 61712 12102
rect 61660 12038 61712 12044
rect 61672 11898 61700 12038
rect 61660 11892 61712 11898
rect 61660 11834 61712 11840
rect 61764 9674 61792 12406
rect 62120 12232 62172 12238
rect 61672 9646 61792 9674
rect 62040 12180 62120 12186
rect 62040 12174 62172 12180
rect 62040 12158 62160 12174
rect 61672 9178 61700 9646
rect 61844 9444 61896 9450
rect 61844 9386 61896 9392
rect 61660 9172 61712 9178
rect 61660 9114 61712 9120
rect 61476 9036 61528 9042
rect 61476 8978 61528 8984
rect 61292 7540 61344 7546
rect 61292 7482 61344 7488
rect 61384 7336 61436 7342
rect 61384 7278 61436 7284
rect 61200 7200 61252 7206
rect 61198 7168 61200 7177
rect 61252 7168 61254 7177
rect 61198 7103 61254 7112
rect 61396 6934 61424 7278
rect 61108 6928 61160 6934
rect 61108 6870 61160 6876
rect 61384 6928 61436 6934
rect 61384 6870 61436 6876
rect 61488 6730 61516 8978
rect 61566 7304 61622 7313
rect 61566 7239 61568 7248
rect 61620 7239 61622 7248
rect 61568 7210 61620 7216
rect 61672 6866 61700 9114
rect 61660 6860 61712 6866
rect 61660 6802 61712 6808
rect 61752 6792 61804 6798
rect 61752 6734 61804 6740
rect 61476 6724 61528 6730
rect 61476 6666 61528 6672
rect 61660 6724 61712 6730
rect 61660 6666 61712 6672
rect 60924 6656 60976 6662
rect 60924 6598 60976 6604
rect 61566 6624 61622 6633
rect 60646 6352 60702 6361
rect 60646 6287 60648 6296
rect 60700 6287 60702 6296
rect 60648 6258 60700 6264
rect 60648 5772 60700 5778
rect 60568 5732 60648 5760
rect 60648 5714 60700 5720
rect 60464 5024 60516 5030
rect 60464 4966 60516 4972
rect 60648 3596 60700 3602
rect 60648 3538 60700 3544
rect 60004 2984 60056 2990
rect 60004 2926 60056 2932
rect 59912 2508 59964 2514
rect 59912 2450 59964 2456
rect 60016 800 60044 2926
rect 60280 2304 60332 2310
rect 60280 2246 60332 2252
rect 60292 800 60320 2246
rect 60660 800 60688 3538
rect 60936 2514 60964 6598
rect 61566 6559 61622 6568
rect 61016 6452 61068 6458
rect 61016 6394 61068 6400
rect 61028 5545 61056 6394
rect 61580 6118 61608 6559
rect 61568 6112 61620 6118
rect 61568 6054 61620 6060
rect 61014 5536 61070 5545
rect 61014 5471 61070 5480
rect 61672 5234 61700 6666
rect 61764 6254 61792 6734
rect 61856 6458 61884 9386
rect 62040 8974 62068 12158
rect 62028 8968 62080 8974
rect 62028 8910 62080 8916
rect 62304 8288 62356 8294
rect 62304 8230 62356 8236
rect 62316 7954 62344 8230
rect 62304 7948 62356 7954
rect 62304 7890 62356 7896
rect 62408 7886 62436 14010
rect 62500 13870 62528 15302
rect 63500 15020 63552 15026
rect 63500 14962 63552 14968
rect 62488 13864 62540 13870
rect 62488 13806 62540 13812
rect 63408 13864 63460 13870
rect 63408 13806 63460 13812
rect 62488 13728 62540 13734
rect 62488 13670 62540 13676
rect 62500 12714 62528 13670
rect 63420 13326 63448 13806
rect 63408 13320 63460 13326
rect 63408 13262 63460 13268
rect 63420 12850 63448 13262
rect 63408 12844 63460 12850
rect 63408 12786 63460 12792
rect 63512 12714 63540 14962
rect 63696 12782 63724 15302
rect 63972 12986 64000 15438
rect 64972 14000 65024 14006
rect 64972 13942 65024 13948
rect 64604 13320 64656 13326
rect 64604 13262 64656 13268
rect 64880 13320 64932 13326
rect 64880 13262 64932 13268
rect 63960 12980 64012 12986
rect 63960 12922 64012 12928
rect 63684 12776 63736 12782
rect 63684 12718 63736 12724
rect 62488 12708 62540 12714
rect 62488 12650 62540 12656
rect 63500 12708 63552 12714
rect 63500 12650 63552 12656
rect 62396 7880 62448 7886
rect 62396 7822 62448 7828
rect 62302 7440 62358 7449
rect 62279 7404 62302 7410
rect 62331 7375 62358 7384
rect 62331 7364 62344 7375
rect 62279 7346 62331 7352
rect 62120 7336 62172 7342
rect 62377 7336 62429 7342
rect 62172 7296 62252 7324
rect 62120 7278 62172 7284
rect 62026 7032 62082 7041
rect 62026 6967 62028 6976
rect 62080 6967 62082 6976
rect 62028 6938 62080 6944
rect 61844 6452 61896 6458
rect 61844 6394 61896 6400
rect 62224 6322 62252 7296
rect 62429 7284 62436 7324
rect 62377 7278 62436 7284
rect 62408 6769 62436 7278
rect 62500 6866 62528 12650
rect 63972 12434 64000 12922
rect 64616 12782 64644 13262
rect 64052 12776 64104 12782
rect 64052 12718 64104 12724
rect 64604 12776 64656 12782
rect 64604 12718 64656 12724
rect 64788 12776 64840 12782
rect 64788 12718 64840 12724
rect 63880 12406 64000 12434
rect 62948 12368 63000 12374
rect 62948 12310 63000 12316
rect 62960 8974 62988 12310
rect 63880 12102 63908 12406
rect 64064 12238 64092 12718
rect 64052 12232 64104 12238
rect 64052 12174 64104 12180
rect 63868 12096 63920 12102
rect 63868 12038 63920 12044
rect 63592 11756 63644 11762
rect 63592 11698 63644 11704
rect 63604 9586 63632 11698
rect 63684 10124 63736 10130
rect 63684 10066 63736 10072
rect 63592 9580 63644 9586
rect 63592 9522 63644 9528
rect 63224 9444 63276 9450
rect 63224 9386 63276 9392
rect 62948 8968 63000 8974
rect 62948 8910 63000 8916
rect 63132 8424 63184 8430
rect 63132 8366 63184 8372
rect 63144 8090 63172 8366
rect 63132 8084 63184 8090
rect 63132 8026 63184 8032
rect 63144 7886 63172 8026
rect 62672 7880 62724 7886
rect 62578 7848 62634 7857
rect 62672 7822 62724 7828
rect 62948 7880 63000 7886
rect 62948 7822 63000 7828
rect 63132 7880 63184 7886
rect 63132 7822 63184 7828
rect 62578 7783 62580 7792
rect 62632 7783 62634 7792
rect 62580 7754 62632 7760
rect 62580 6996 62632 7002
rect 62580 6938 62632 6944
rect 62488 6860 62540 6866
rect 62488 6802 62540 6808
rect 62394 6760 62450 6769
rect 62394 6695 62450 6704
rect 62396 6452 62448 6458
rect 62396 6394 62448 6400
rect 62212 6316 62264 6322
rect 62264 6276 62344 6304
rect 62212 6258 62264 6264
rect 61752 6248 61804 6254
rect 61752 6190 61804 6196
rect 62120 5772 62172 5778
rect 62120 5714 62172 5720
rect 62132 5250 62160 5714
rect 62316 5710 62344 6276
rect 62304 5704 62356 5710
rect 62304 5646 62356 5652
rect 61948 5234 62160 5250
rect 61660 5228 61712 5234
rect 61660 5170 61712 5176
rect 61936 5228 62160 5234
rect 61988 5222 62160 5228
rect 61936 5170 61988 5176
rect 62132 4554 62160 5222
rect 62212 5160 62264 5166
rect 62212 5102 62264 5108
rect 62316 5114 62344 5646
rect 62408 5234 62436 6394
rect 62396 5228 62448 5234
rect 62396 5170 62448 5176
rect 62488 5160 62540 5166
rect 62316 5108 62488 5114
rect 62316 5102 62540 5108
rect 62120 4548 62172 4554
rect 62120 4490 62172 4496
rect 62224 3670 62252 5102
rect 62316 5086 62528 5102
rect 62212 3664 62264 3670
rect 62212 3606 62264 3612
rect 61752 3596 61804 3602
rect 61752 3538 61804 3544
rect 61568 3460 61620 3466
rect 61568 3402 61620 3408
rect 61580 3058 61608 3402
rect 61568 3052 61620 3058
rect 61568 2994 61620 3000
rect 61016 2984 61068 2990
rect 61016 2926 61068 2932
rect 60924 2508 60976 2514
rect 60924 2450 60976 2456
rect 61028 800 61056 2926
rect 61292 2576 61344 2582
rect 61292 2518 61344 2524
rect 61304 2106 61332 2518
rect 61384 2304 61436 2310
rect 61384 2246 61436 2252
rect 61292 2100 61344 2106
rect 61292 2042 61344 2048
rect 61396 800 61424 2246
rect 61764 800 61792 3538
rect 62120 2984 62172 2990
rect 62120 2926 62172 2932
rect 62132 800 62160 2926
rect 62488 2304 62540 2310
rect 62488 2246 62540 2252
rect 62500 800 62528 2246
rect 62592 1766 62620 6938
rect 62684 6458 62712 7822
rect 62856 7812 62908 7818
rect 62856 7754 62908 7760
rect 62764 7404 62816 7410
rect 62764 7346 62816 7352
rect 62776 7290 62804 7346
rect 62868 7290 62896 7754
rect 62776 7262 62896 7290
rect 62764 6656 62816 6662
rect 62764 6598 62816 6604
rect 62672 6452 62724 6458
rect 62672 6394 62724 6400
rect 62672 6248 62724 6254
rect 62672 6190 62724 6196
rect 62684 1902 62712 6190
rect 62776 2582 62804 6598
rect 62868 6372 62896 7262
rect 62960 6474 62988 7822
rect 63130 6488 63186 6497
rect 62960 6446 63080 6474
rect 62948 6384 63000 6390
rect 62868 6344 62948 6372
rect 62948 6326 63000 6332
rect 62960 5778 62988 6326
rect 62948 5772 63000 5778
rect 62948 5714 63000 5720
rect 62856 3596 62908 3602
rect 62856 3538 62908 3544
rect 62764 2576 62816 2582
rect 62764 2518 62816 2524
rect 62672 1896 62724 1902
rect 62672 1838 62724 1844
rect 62580 1760 62632 1766
rect 62580 1702 62632 1708
rect 62868 800 62896 3538
rect 63052 1630 63080 6446
rect 63130 6423 63132 6432
rect 63184 6423 63186 6432
rect 63132 6394 63184 6400
rect 63130 5944 63186 5953
rect 63130 5879 63132 5888
rect 63184 5879 63186 5888
rect 63132 5850 63184 5856
rect 63236 5370 63264 9386
rect 63316 9036 63368 9042
rect 63316 8978 63368 8984
rect 63592 9036 63644 9042
rect 63592 8978 63644 8984
rect 63328 7546 63356 8978
rect 63500 7948 63552 7954
rect 63500 7890 63552 7896
rect 63316 7540 63368 7546
rect 63316 7482 63368 7488
rect 63314 7440 63370 7449
rect 63314 7375 63316 7384
rect 63368 7375 63370 7384
rect 63316 7346 63368 7352
rect 63314 6760 63370 6769
rect 63314 6695 63316 6704
rect 63368 6695 63370 6704
rect 63316 6666 63368 6672
rect 63408 6656 63460 6662
rect 63408 6598 63460 6604
rect 63420 6322 63448 6598
rect 63408 6316 63460 6322
rect 63408 6258 63460 6264
rect 63420 6118 63448 6258
rect 63408 6112 63460 6118
rect 63408 6054 63460 6060
rect 63408 5772 63460 5778
rect 63408 5714 63460 5720
rect 63420 5681 63448 5714
rect 63406 5672 63462 5681
rect 63406 5607 63462 5616
rect 63512 5386 63540 7890
rect 63604 6934 63632 8978
rect 63592 6928 63644 6934
rect 63592 6870 63644 6876
rect 63696 6866 63724 10066
rect 63880 7313 63908 12038
rect 64064 11694 64092 12174
rect 64052 11688 64104 11694
rect 64052 11630 64104 11636
rect 64604 10056 64656 10062
rect 64604 9998 64656 10004
rect 64512 9512 64564 9518
rect 64512 9454 64564 9460
rect 64420 8356 64472 8362
rect 64420 8298 64472 8304
rect 64432 7954 64460 8298
rect 64420 7948 64472 7954
rect 64420 7890 64472 7896
rect 64144 7880 64196 7886
rect 64144 7822 64196 7828
rect 64234 7848 64290 7857
rect 63866 7304 63922 7313
rect 63866 7239 63922 7248
rect 63684 6860 63736 6866
rect 63684 6802 63736 6808
rect 63592 6112 63644 6118
rect 63592 6054 63644 6060
rect 63604 5574 63632 6054
rect 63592 5568 63644 5574
rect 63592 5510 63644 5516
rect 63224 5364 63276 5370
rect 63512 5358 63724 5386
rect 63224 5306 63276 5312
rect 63500 5024 63552 5030
rect 63500 4966 63552 4972
rect 63224 2984 63276 2990
rect 63224 2926 63276 2932
rect 63040 1624 63092 1630
rect 63040 1566 63092 1572
rect 63236 800 63264 2926
rect 63512 2582 63540 4966
rect 63500 2576 63552 2582
rect 63500 2518 63552 2524
rect 63592 2304 63644 2310
rect 63592 2246 63644 2252
rect 63604 800 63632 2246
rect 63696 1970 63724 5358
rect 63880 5166 63908 7239
rect 64156 6798 64184 7822
rect 64234 7783 64236 7792
rect 64288 7783 64290 7792
rect 64236 7754 64288 7760
rect 64418 6896 64474 6905
rect 64418 6831 64474 6840
rect 64432 6798 64460 6831
rect 64144 6792 64196 6798
rect 64064 6752 64144 6780
rect 64064 6254 64092 6752
rect 64144 6734 64196 6740
rect 64420 6792 64472 6798
rect 64420 6734 64472 6740
rect 64524 6390 64552 9454
rect 64616 7546 64644 9998
rect 64800 9382 64828 12718
rect 64892 10198 64920 13262
rect 64880 10192 64932 10198
rect 64880 10134 64932 10140
rect 64984 9674 65012 13942
rect 65168 13734 65196 15966
rect 65248 15904 65300 15910
rect 65248 15846 65300 15852
rect 65156 13728 65208 13734
rect 65156 13670 65208 13676
rect 65260 13530 65288 15846
rect 65248 13524 65300 13530
rect 65248 13466 65300 13472
rect 65352 13394 65380 15982
rect 65536 14958 65564 16594
rect 65660 16348 65956 16368
rect 65716 16346 65740 16348
rect 65796 16346 65820 16348
rect 65876 16346 65900 16348
rect 65738 16294 65740 16346
rect 65802 16294 65814 16346
rect 65876 16294 65878 16346
rect 65716 16292 65740 16294
rect 65796 16292 65820 16294
rect 65876 16292 65900 16294
rect 65660 16272 65956 16292
rect 66088 16130 66116 18770
rect 67088 18692 67140 18698
rect 67088 18634 67140 18640
rect 66168 18624 66220 18630
rect 66168 18566 66220 18572
rect 66904 18624 66956 18630
rect 66904 18566 66956 18572
rect 66180 17202 66208 18566
rect 66168 17196 66220 17202
rect 66168 17138 66220 17144
rect 66916 17134 66944 18566
rect 67100 17134 67128 18634
rect 66904 17128 66956 17134
rect 66904 17070 66956 17076
rect 67088 17128 67140 17134
rect 67088 17070 67140 17076
rect 66168 16992 66220 16998
rect 66168 16934 66220 16940
rect 66352 16992 66404 16998
rect 66352 16934 66404 16940
rect 66180 16454 66208 16934
rect 66364 16726 66392 16934
rect 66352 16720 66404 16726
rect 66352 16662 66404 16668
rect 66260 16584 66312 16590
rect 66260 16526 66312 16532
rect 66168 16448 66220 16454
rect 66168 16390 66220 16396
rect 65708 16108 65760 16114
rect 65708 16050 65760 16056
rect 65996 16102 66116 16130
rect 66180 16114 66208 16390
rect 66168 16108 66220 16114
rect 65720 15434 65748 16050
rect 65996 15570 66024 16102
rect 66168 16050 66220 16056
rect 66076 16040 66128 16046
rect 66272 15994 66300 16526
rect 66128 15988 66300 15994
rect 66076 15982 66300 15988
rect 66088 15966 66300 15982
rect 65984 15564 66036 15570
rect 65984 15506 66036 15512
rect 65708 15428 65760 15434
rect 65708 15370 65760 15376
rect 65660 15260 65956 15280
rect 65716 15258 65740 15260
rect 65796 15258 65820 15260
rect 65876 15258 65900 15260
rect 65738 15206 65740 15258
rect 65802 15206 65814 15258
rect 65876 15206 65878 15258
rect 65716 15204 65740 15206
rect 65796 15204 65820 15206
rect 65876 15204 65900 15206
rect 65660 15184 65956 15204
rect 65524 14952 65576 14958
rect 65524 14894 65576 14900
rect 66364 14890 66392 16662
rect 66916 16590 66944 17070
rect 67100 16658 67128 17070
rect 67088 16652 67140 16658
rect 67088 16594 67140 16600
rect 66904 16584 66956 16590
rect 66904 16526 66956 16532
rect 67836 16182 67864 18770
rect 67824 16176 67876 16182
rect 67824 16118 67876 16124
rect 67640 15360 67692 15366
rect 67640 15302 67692 15308
rect 66352 14884 66404 14890
rect 66352 14826 66404 14832
rect 65524 14816 65576 14822
rect 65524 14758 65576 14764
rect 65536 13938 65564 14758
rect 65660 14172 65956 14192
rect 65716 14170 65740 14172
rect 65796 14170 65820 14172
rect 65876 14170 65900 14172
rect 65738 14118 65740 14170
rect 65802 14118 65814 14170
rect 65876 14118 65878 14170
rect 65716 14116 65740 14118
rect 65796 14116 65820 14118
rect 65876 14116 65900 14118
rect 65660 14096 65956 14116
rect 66904 14000 66956 14006
rect 66904 13942 66956 13948
rect 65524 13932 65576 13938
rect 65524 13874 65576 13880
rect 66260 13728 66312 13734
rect 66260 13670 66312 13676
rect 66272 13530 66300 13670
rect 66260 13524 66312 13530
rect 66260 13466 66312 13472
rect 65340 13388 65392 13394
rect 65340 13330 65392 13336
rect 65064 12640 65116 12646
rect 65064 12582 65116 12588
rect 64892 9646 65012 9674
rect 64788 9376 64840 9382
rect 64788 9318 64840 9324
rect 64604 7540 64656 7546
rect 64604 7482 64656 7488
rect 64788 7404 64840 7410
rect 64892 7392 64920 9646
rect 65076 8974 65104 12582
rect 65352 12102 65380 13330
rect 65660 13084 65956 13104
rect 65716 13082 65740 13084
rect 65796 13082 65820 13084
rect 65876 13082 65900 13084
rect 65738 13030 65740 13082
rect 65802 13030 65814 13082
rect 65876 13030 65878 13082
rect 65716 13028 65740 13030
rect 65796 13028 65820 13030
rect 65876 13028 65900 13030
rect 65660 13008 65956 13028
rect 65524 12776 65576 12782
rect 65524 12718 65576 12724
rect 65156 12096 65208 12102
rect 65156 12038 65208 12044
rect 65340 12096 65392 12102
rect 65340 12038 65392 12044
rect 65064 8968 65116 8974
rect 65064 8910 65116 8916
rect 65076 8498 65104 8910
rect 65064 8492 65116 8498
rect 65064 8434 65116 8440
rect 64840 7364 64920 7392
rect 65064 7404 65116 7410
rect 64788 7346 64840 7352
rect 65064 7346 65116 7352
rect 64788 7200 64840 7206
rect 64788 7142 64840 7148
rect 64800 7002 64828 7142
rect 64604 6996 64656 7002
rect 64604 6938 64656 6944
rect 64788 6996 64840 7002
rect 64788 6938 64840 6944
rect 64616 6798 64644 6938
rect 64786 6896 64842 6905
rect 64786 6831 64842 6840
rect 64800 6798 64828 6831
rect 64604 6792 64656 6798
rect 64604 6734 64656 6740
rect 64788 6792 64840 6798
rect 64788 6734 64840 6740
rect 65076 6730 65104 7346
rect 65168 7177 65196 12038
rect 65432 10600 65484 10606
rect 65432 10542 65484 10548
rect 65444 10062 65472 10542
rect 65432 10056 65484 10062
rect 65432 9998 65484 10004
rect 65444 9518 65472 9998
rect 65432 9512 65484 9518
rect 65432 9454 65484 9460
rect 65248 9444 65300 9450
rect 65248 9386 65300 9392
rect 65154 7168 65210 7177
rect 65154 7103 65210 7112
rect 64880 6724 64932 6730
rect 64880 6666 64932 6672
rect 65064 6724 65116 6730
rect 65064 6666 65116 6672
rect 65156 6724 65208 6730
rect 65156 6666 65208 6672
rect 64512 6384 64564 6390
rect 64512 6326 64564 6332
rect 64602 6352 64658 6361
rect 64420 6316 64472 6322
rect 64602 6287 64658 6296
rect 64420 6258 64472 6264
rect 64052 6248 64104 6254
rect 64052 6190 64104 6196
rect 64064 5710 64092 6190
rect 64432 6089 64460 6258
rect 64616 6186 64644 6287
rect 64604 6180 64656 6186
rect 64604 6122 64656 6128
rect 64418 6080 64474 6089
rect 64418 6015 64474 6024
rect 64234 5808 64290 5817
rect 64234 5743 64236 5752
rect 64288 5743 64290 5752
rect 64236 5714 64288 5720
rect 64052 5704 64104 5710
rect 64052 5646 64104 5652
rect 64328 5704 64380 5710
rect 64328 5646 64380 5652
rect 64602 5672 64658 5681
rect 63868 5160 63920 5166
rect 63868 5102 63920 5108
rect 64340 4298 64368 5646
rect 64892 5642 64920 6666
rect 64602 5607 64604 5616
rect 64656 5607 64658 5616
rect 64880 5636 64932 5642
rect 64604 5578 64656 5584
rect 64880 5578 64932 5584
rect 64788 5568 64840 5574
rect 64788 5510 64840 5516
rect 64800 5234 64828 5510
rect 64788 5228 64840 5234
rect 64788 5170 64840 5176
rect 64248 4270 64368 4298
rect 63960 3596 64012 3602
rect 63960 3538 64012 3544
rect 63684 1964 63736 1970
rect 63684 1906 63736 1912
rect 63972 800 64000 3538
rect 64248 2378 64276 4270
rect 65064 3596 65116 3602
rect 65064 3538 65116 3544
rect 64328 2984 64380 2990
rect 64328 2926 64380 2932
rect 64236 2372 64288 2378
rect 64236 2314 64288 2320
rect 64340 800 64368 2926
rect 64696 2372 64748 2378
rect 64696 2314 64748 2320
rect 64708 800 64736 2314
rect 65076 800 65104 3538
rect 65168 1970 65196 6666
rect 65260 6118 65288 9386
rect 65340 9376 65392 9382
rect 65340 9318 65392 9324
rect 65352 8090 65380 9318
rect 65536 9110 65564 12718
rect 66076 12368 66128 12374
rect 66076 12310 66128 12316
rect 65660 11996 65956 12016
rect 65716 11994 65740 11996
rect 65796 11994 65820 11996
rect 65876 11994 65900 11996
rect 65738 11942 65740 11994
rect 65802 11942 65814 11994
rect 65876 11942 65878 11994
rect 65716 11940 65740 11942
rect 65796 11940 65820 11942
rect 65876 11940 65900 11942
rect 65660 11920 65956 11940
rect 65984 11756 66036 11762
rect 65984 11698 66036 11704
rect 65660 10908 65956 10928
rect 65716 10906 65740 10908
rect 65796 10906 65820 10908
rect 65876 10906 65900 10908
rect 65738 10854 65740 10906
rect 65802 10854 65814 10906
rect 65876 10854 65878 10906
rect 65716 10852 65740 10854
rect 65796 10852 65820 10854
rect 65876 10852 65900 10854
rect 65660 10832 65956 10852
rect 65660 9820 65956 9840
rect 65716 9818 65740 9820
rect 65796 9818 65820 9820
rect 65876 9818 65900 9820
rect 65738 9766 65740 9818
rect 65802 9766 65814 9818
rect 65876 9766 65878 9818
rect 65716 9764 65740 9766
rect 65796 9764 65820 9766
rect 65876 9764 65900 9766
rect 65660 9744 65956 9764
rect 65996 9586 66024 11698
rect 65984 9580 66036 9586
rect 65984 9522 66036 9528
rect 65800 9512 65852 9518
rect 65800 9454 65852 9460
rect 65524 9104 65576 9110
rect 65524 9046 65576 9052
rect 65812 9042 65840 9454
rect 66088 9110 66116 12310
rect 66272 11558 66300 13466
rect 66628 13320 66680 13326
rect 66628 13262 66680 13268
rect 66640 12850 66668 13262
rect 66628 12844 66680 12850
rect 66628 12786 66680 12792
rect 66640 12238 66668 12786
rect 66628 12232 66680 12238
rect 66628 12174 66680 12180
rect 66260 11552 66312 11558
rect 66260 11494 66312 11500
rect 66076 9104 66128 9110
rect 66076 9046 66128 9052
rect 65800 9036 65852 9042
rect 65800 8978 65852 8984
rect 65660 8732 65956 8752
rect 65716 8730 65740 8732
rect 65796 8730 65820 8732
rect 65876 8730 65900 8732
rect 65738 8678 65740 8730
rect 65802 8678 65814 8730
rect 65876 8678 65878 8730
rect 65716 8676 65740 8678
rect 65796 8676 65820 8678
rect 65876 8676 65900 8678
rect 65660 8656 65956 8676
rect 65340 8084 65392 8090
rect 65340 8026 65392 8032
rect 65524 7880 65576 7886
rect 65524 7822 65576 7828
rect 65432 7744 65484 7750
rect 65432 7686 65484 7692
rect 65338 7168 65394 7177
rect 65338 7103 65394 7112
rect 65248 6112 65300 6118
rect 65248 6054 65300 6060
rect 65246 5944 65302 5953
rect 65246 5879 65248 5888
rect 65300 5879 65302 5888
rect 65248 5850 65300 5856
rect 65246 5808 65302 5817
rect 65352 5778 65380 7103
rect 65444 6934 65472 7686
rect 65536 7274 65564 7822
rect 65660 7644 65956 7664
rect 65716 7642 65740 7644
rect 65796 7642 65820 7644
rect 65876 7642 65900 7644
rect 65738 7590 65740 7642
rect 65802 7590 65814 7642
rect 65876 7590 65878 7642
rect 65716 7588 65740 7590
rect 65796 7588 65820 7590
rect 65876 7588 65900 7590
rect 65660 7568 65956 7588
rect 66272 7274 66300 11494
rect 65524 7268 65576 7274
rect 65524 7210 65576 7216
rect 66076 7268 66128 7274
rect 66076 7210 66128 7216
rect 66260 7268 66312 7274
rect 66260 7210 66312 7216
rect 65432 6928 65484 6934
rect 65432 6870 65484 6876
rect 65432 6792 65484 6798
rect 65430 6760 65432 6769
rect 65484 6760 65486 6769
rect 65430 6695 65486 6704
rect 65524 6656 65576 6662
rect 65522 6624 65524 6633
rect 65576 6624 65578 6633
rect 65522 6559 65578 6568
rect 65660 6556 65956 6576
rect 65716 6554 65740 6556
rect 65796 6554 65820 6556
rect 65876 6554 65900 6556
rect 65738 6502 65740 6554
rect 65802 6502 65814 6554
rect 65876 6502 65878 6554
rect 65716 6500 65740 6502
rect 65796 6500 65820 6502
rect 65876 6500 65900 6502
rect 65660 6480 65956 6500
rect 65800 6316 65852 6322
rect 65800 6258 65852 6264
rect 65432 6248 65484 6254
rect 65432 6190 65484 6196
rect 65444 6118 65472 6190
rect 65432 6112 65484 6118
rect 65432 6054 65484 6060
rect 65246 5743 65302 5752
rect 65340 5772 65392 5778
rect 65260 5710 65288 5743
rect 65340 5714 65392 5720
rect 65248 5704 65300 5710
rect 65248 5646 65300 5652
rect 65248 5568 65300 5574
rect 65248 5510 65300 5516
rect 65260 2582 65288 5510
rect 65444 5012 65472 6054
rect 65524 5840 65576 5846
rect 65524 5782 65576 5788
rect 65536 5545 65564 5782
rect 65812 5681 65840 6258
rect 65984 6248 66036 6254
rect 65984 6190 66036 6196
rect 65996 6089 66024 6190
rect 65982 6080 66038 6089
rect 65982 6015 66038 6024
rect 65798 5672 65854 5681
rect 65798 5607 65854 5616
rect 65522 5536 65578 5545
rect 65522 5471 65578 5480
rect 65660 5468 65956 5488
rect 65716 5466 65740 5468
rect 65796 5466 65820 5468
rect 65876 5466 65900 5468
rect 65738 5414 65740 5466
rect 65802 5414 65814 5466
rect 65876 5414 65878 5466
rect 65716 5412 65740 5414
rect 65796 5412 65820 5414
rect 65876 5412 65900 5414
rect 65660 5392 65956 5412
rect 65352 4984 65472 5012
rect 65352 2650 65380 4984
rect 65660 4380 65956 4400
rect 65716 4378 65740 4380
rect 65796 4378 65820 4380
rect 65876 4378 65900 4380
rect 65738 4326 65740 4378
rect 65802 4326 65814 4378
rect 65876 4326 65878 4378
rect 65716 4324 65740 4326
rect 65796 4324 65820 4326
rect 65876 4324 65900 4326
rect 65660 4304 65956 4324
rect 65660 3292 65956 3312
rect 65716 3290 65740 3292
rect 65796 3290 65820 3292
rect 65876 3290 65900 3292
rect 65738 3238 65740 3290
rect 65802 3238 65814 3290
rect 65876 3238 65878 3290
rect 65716 3236 65740 3238
rect 65796 3236 65820 3238
rect 65876 3236 65900 3238
rect 65660 3216 65956 3236
rect 65432 2984 65484 2990
rect 65432 2926 65484 2932
rect 65340 2644 65392 2650
rect 65340 2586 65392 2592
rect 65248 2576 65300 2582
rect 65248 2518 65300 2524
rect 65156 1964 65208 1970
rect 65156 1906 65208 1912
rect 65444 800 65472 2926
rect 65984 2304 66036 2310
rect 65984 2246 66036 2252
rect 65660 2204 65956 2224
rect 65716 2202 65740 2204
rect 65796 2202 65820 2204
rect 65876 2202 65900 2204
rect 65738 2150 65740 2202
rect 65802 2150 65814 2202
rect 65876 2150 65878 2202
rect 65716 2148 65740 2150
rect 65796 2148 65820 2150
rect 65876 2148 65900 2150
rect 65660 2128 65956 2148
rect 65996 1170 66024 2246
rect 66088 1698 66116 7210
rect 66272 7041 66300 7210
rect 66258 7032 66314 7041
rect 66258 6967 66314 6976
rect 66916 6361 66944 13942
rect 67652 13870 67680 15302
rect 68192 14272 68244 14278
rect 68192 14214 68244 14220
rect 68284 14272 68336 14278
rect 68284 14214 68336 14220
rect 67640 13864 67692 13870
rect 67640 13806 67692 13812
rect 68008 13728 68060 13734
rect 68008 13670 68060 13676
rect 67456 13320 67508 13326
rect 67456 13262 67508 13268
rect 67088 13184 67140 13190
rect 67088 13126 67140 13132
rect 66996 8968 67048 8974
rect 66996 8910 67048 8916
rect 66902 6352 66958 6361
rect 66902 6287 66958 6296
rect 67008 6254 67036 8910
rect 67100 6662 67128 13126
rect 67272 12980 67324 12986
rect 67272 12922 67324 12928
rect 67180 12096 67232 12102
rect 67180 12038 67232 12044
rect 67192 11694 67220 12038
rect 67180 11688 67232 11694
rect 67180 11630 67232 11636
rect 67192 11218 67220 11630
rect 67180 11212 67232 11218
rect 67180 11154 67232 11160
rect 67284 8430 67312 12922
rect 67468 9586 67496 13262
rect 68020 12850 68048 13670
rect 68008 12844 68060 12850
rect 68008 12786 68060 12792
rect 67548 11144 67600 11150
rect 67548 11086 67600 11092
rect 67560 10198 67588 11086
rect 67548 10192 67600 10198
rect 67548 10134 67600 10140
rect 67456 9580 67508 9586
rect 67456 9522 67508 9528
rect 67640 8628 67692 8634
rect 67640 8570 67692 8576
rect 67272 8424 67324 8430
rect 67272 8366 67324 8372
rect 67088 6656 67140 6662
rect 67088 6598 67140 6604
rect 66996 6248 67048 6254
rect 66996 6190 67048 6196
rect 66812 6112 66864 6118
rect 66812 6054 66864 6060
rect 66168 4072 66220 4078
rect 66168 4014 66220 4020
rect 66076 1692 66128 1698
rect 66076 1634 66128 1640
rect 65812 1142 66024 1170
rect 65812 800 65840 1142
rect 66180 800 66208 4014
rect 66536 3596 66588 3602
rect 66536 3538 66588 3544
rect 66548 800 66576 3538
rect 66628 2984 66680 2990
rect 66628 2926 66680 2932
rect 66640 1222 66668 2926
rect 66824 2582 66852 6054
rect 67272 4072 67324 4078
rect 67272 4014 67324 4020
rect 66812 2576 66864 2582
rect 66812 2518 66864 2524
rect 66904 2304 66956 2310
rect 66904 2246 66956 2252
rect 66628 1216 66680 1222
rect 66628 1158 66680 1164
rect 66916 800 66944 2246
rect 67284 800 67312 4014
rect 67548 3392 67600 3398
rect 67548 3334 67600 3340
rect 67560 3194 67588 3334
rect 67652 3194 67680 8570
rect 67916 6112 67968 6118
rect 67916 6054 67968 6060
rect 67824 5568 67876 5574
rect 67824 5510 67876 5516
rect 67732 3596 67784 3602
rect 67732 3538 67784 3544
rect 67548 3188 67600 3194
rect 67548 3130 67600 3136
rect 67640 3188 67692 3194
rect 67640 3130 67692 3136
rect 67744 1154 67772 3538
rect 67836 2582 67864 5510
rect 67824 2576 67876 2582
rect 67824 2518 67876 2524
rect 67928 2514 67956 6054
rect 68020 5914 68048 12786
rect 68100 7268 68152 7274
rect 68100 7210 68152 7216
rect 68112 6254 68140 7210
rect 68100 6248 68152 6254
rect 68100 6190 68152 6196
rect 68008 5908 68060 5914
rect 68008 5850 68060 5856
rect 68204 5710 68232 14214
rect 68296 7206 68324 14214
rect 68480 12646 68508 18770
rect 68560 14952 68612 14958
rect 68560 14894 68612 14900
rect 68572 14482 68600 14894
rect 68560 14476 68612 14482
rect 68560 14418 68612 14424
rect 68468 12640 68520 12646
rect 68468 12582 68520 12588
rect 68572 11558 68600 14418
rect 68664 13734 68692 19110
rect 69676 18290 69704 117098
rect 72436 116278 72464 117098
rect 73068 117088 73120 117094
rect 73068 117030 73120 117036
rect 72424 116272 72476 116278
rect 72424 116214 72476 116220
rect 72424 116068 72476 116074
rect 72424 116010 72476 116016
rect 72148 20052 72200 20058
rect 72148 19994 72200 20000
rect 71320 19236 71372 19242
rect 71320 19178 71372 19184
rect 71136 18692 71188 18698
rect 71136 18634 71188 18640
rect 70860 18624 70912 18630
rect 70860 18566 70912 18572
rect 69664 18284 69716 18290
rect 69664 18226 69716 18232
rect 70768 18080 70820 18086
rect 70768 18022 70820 18028
rect 70400 17332 70452 17338
rect 70400 17274 70452 17280
rect 69848 17128 69900 17134
rect 69848 17070 69900 17076
rect 69860 16726 69888 17070
rect 69940 17060 69992 17066
rect 69940 17002 69992 17008
rect 69848 16720 69900 16726
rect 69848 16662 69900 16668
rect 68928 16448 68980 16454
rect 68928 16390 68980 16396
rect 68940 15502 68968 16390
rect 69020 16244 69072 16250
rect 69020 16186 69072 16192
rect 68928 15496 68980 15502
rect 68928 15438 68980 15444
rect 68940 14890 68968 15438
rect 68928 14884 68980 14890
rect 68928 14826 68980 14832
rect 69032 13870 69060 16186
rect 69848 15904 69900 15910
rect 69848 15846 69900 15852
rect 69860 15570 69888 15846
rect 69848 15564 69900 15570
rect 69848 15506 69900 15512
rect 69388 15496 69440 15502
rect 69388 15438 69440 15444
rect 69112 14408 69164 14414
rect 69112 14350 69164 14356
rect 69124 13938 69152 14350
rect 69112 13932 69164 13938
rect 69112 13874 69164 13880
rect 69020 13864 69072 13870
rect 69020 13806 69072 13812
rect 68652 13728 68704 13734
rect 68652 13670 68704 13676
rect 68664 12102 68692 13670
rect 69400 12850 69428 15438
rect 69756 14476 69808 14482
rect 69756 14418 69808 14424
rect 69572 14000 69624 14006
rect 69572 13942 69624 13948
rect 69388 12844 69440 12850
rect 69388 12786 69440 12792
rect 68652 12096 68704 12102
rect 68652 12038 68704 12044
rect 68560 11552 68612 11558
rect 68560 11494 68612 11500
rect 68572 7954 68600 11494
rect 68664 8294 68692 12038
rect 68652 8288 68704 8294
rect 68652 8230 68704 8236
rect 68560 7948 68612 7954
rect 68560 7890 68612 7896
rect 68284 7200 68336 7206
rect 68284 7142 68336 7148
rect 69112 6384 69164 6390
rect 69112 6326 69164 6332
rect 69020 6112 69072 6118
rect 69020 6054 69072 6060
rect 68928 5908 68980 5914
rect 68928 5850 68980 5856
rect 68940 5778 68968 5850
rect 68928 5772 68980 5778
rect 68928 5714 68980 5720
rect 68192 5704 68244 5710
rect 68192 5646 68244 5652
rect 68008 4548 68060 4554
rect 68008 4490 68060 4496
rect 68020 3058 68048 4490
rect 68376 4072 68428 4078
rect 68376 4014 68428 4020
rect 68282 3768 68338 3777
rect 68282 3703 68338 3712
rect 68296 3670 68324 3703
rect 68284 3664 68336 3670
rect 68284 3606 68336 3612
rect 68008 3052 68060 3058
rect 68008 2994 68060 3000
rect 67916 2508 67968 2514
rect 67916 2450 67968 2456
rect 68008 2508 68060 2514
rect 68008 2450 68060 2456
rect 68020 2394 68048 2450
rect 67836 2366 68048 2394
rect 67732 1148 67784 1154
rect 67732 1090 67784 1096
rect 67836 1034 67864 2366
rect 68008 2304 68060 2310
rect 68008 2246 68060 2252
rect 67652 1006 67864 1034
rect 67652 800 67680 1006
rect 68020 800 68048 2246
rect 68388 800 68416 4014
rect 68558 3360 68614 3369
rect 68558 3295 68614 3304
rect 68572 3194 68600 3295
rect 68560 3188 68612 3194
rect 68560 3130 68612 3136
rect 68650 2952 68706 2961
rect 68650 2887 68652 2896
rect 68704 2887 68706 2896
rect 68652 2858 68704 2864
rect 68836 2848 68888 2854
rect 68836 2790 68888 2796
rect 68744 1148 68796 1154
rect 68744 1090 68796 1096
rect 68756 800 68784 1090
rect 59820 672 59872 678
rect 59820 614 59872 620
rect 60002 0 60058 800
rect 60278 0 60334 800
rect 60646 0 60702 800
rect 61014 0 61070 800
rect 61382 0 61438 800
rect 61750 0 61806 800
rect 62118 0 62174 800
rect 62486 0 62542 800
rect 62854 0 62910 800
rect 63222 0 63278 800
rect 63590 0 63646 800
rect 63958 0 64014 800
rect 64326 0 64382 800
rect 64694 0 64750 800
rect 65062 0 65118 800
rect 65430 0 65486 800
rect 65798 0 65854 800
rect 66166 0 66222 800
rect 66534 0 66590 800
rect 66902 0 66958 800
rect 67270 0 67326 800
rect 67638 0 67694 800
rect 68006 0 68062 800
rect 68374 0 68430 800
rect 68742 0 68798 800
rect 68848 610 68876 2790
rect 69032 2582 69060 6054
rect 69124 3602 69152 6326
rect 69584 6322 69612 13942
rect 69768 13258 69796 14418
rect 69848 13864 69900 13870
rect 69952 13852 69980 17002
rect 70216 16992 70268 16998
rect 70216 16934 70268 16940
rect 70228 16046 70256 16934
rect 70412 16590 70440 17274
rect 70780 17134 70808 18022
rect 70872 17338 70900 18566
rect 70860 17332 70912 17338
rect 70860 17274 70912 17280
rect 71148 17134 71176 18634
rect 71332 17134 71360 19178
rect 72160 18222 72188 19994
rect 72436 18834 72464 116010
rect 73080 22094 73108 117030
rect 76944 116346 76972 117166
rect 77116 117156 77168 117162
rect 77116 117098 77168 117104
rect 79048 117156 79100 117162
rect 79048 117098 79100 117104
rect 81808 117156 81860 117162
rect 81808 117098 81860 117104
rect 86592 117156 86644 117162
rect 86592 117098 86644 117104
rect 88432 117156 88484 117162
rect 88432 117098 88484 117104
rect 91376 117156 91428 117162
rect 91376 117098 91428 117104
rect 93216 117156 93268 117162
rect 93216 117098 93268 117104
rect 96068 117156 96120 117162
rect 96068 117098 96120 117104
rect 77128 116346 77156 117098
rect 76932 116340 76984 116346
rect 76932 116282 76984 116288
rect 77116 116340 77168 116346
rect 77116 116282 77168 116288
rect 79060 116278 79088 117098
rect 81020 116988 81316 117008
rect 81076 116986 81100 116988
rect 81156 116986 81180 116988
rect 81236 116986 81260 116988
rect 81098 116934 81100 116986
rect 81162 116934 81174 116986
rect 81236 116934 81238 116986
rect 81076 116932 81100 116934
rect 81156 116932 81180 116934
rect 81236 116932 81260 116934
rect 81020 116912 81316 116932
rect 81820 116346 81848 117098
rect 86604 116346 86632 117098
rect 88444 116550 88472 117098
rect 88432 116544 88484 116550
rect 88432 116486 88484 116492
rect 91388 116346 91416 117098
rect 93228 116618 93256 117098
rect 93216 116612 93268 116618
rect 93216 116554 93268 116560
rect 96080 116346 96108 117098
rect 97644 117094 97672 117166
rect 101220 117156 101272 117162
rect 101220 117098 101272 117104
rect 103060 117156 103112 117162
rect 103060 117098 103112 117104
rect 105360 117156 105412 117162
rect 105360 117098 105412 117104
rect 107200 117156 107252 117162
rect 107200 117098 107252 117104
rect 110236 117156 110288 117162
rect 110236 117098 110288 117104
rect 111156 117156 111208 117162
rect 111156 117098 111208 117104
rect 114928 117156 114980 117162
rect 114928 117098 114980 117104
rect 116676 117156 116728 117162
rect 116676 117098 116728 117104
rect 119620 117156 119672 117162
rect 119620 117098 119672 117104
rect 121736 117156 121788 117162
rect 121736 117098 121788 117104
rect 124312 117156 124364 117162
rect 124312 117098 124364 117104
rect 128912 117156 128964 117162
rect 128912 117098 128964 117104
rect 130752 117156 130804 117162
rect 130752 117098 130804 117104
rect 133512 117156 133564 117162
rect 133512 117098 133564 117104
rect 135444 117156 135496 117162
rect 135444 117098 135496 117104
rect 138020 117156 138072 117162
rect 138020 117098 138072 117104
rect 140412 117156 140464 117162
rect 140412 117098 140464 117104
rect 143172 117156 143224 117162
rect 143172 117098 143224 117104
rect 144552 117156 144604 117162
rect 144552 117098 144604 117104
rect 146760 117156 146812 117162
rect 146760 117098 146812 117104
rect 149520 117156 149572 117162
rect 149520 117098 149572 117104
rect 150900 117156 150952 117162
rect 150900 117098 150952 117104
rect 154120 117156 154172 117162
rect 154120 117098 154172 117104
rect 154856 117156 154908 117162
rect 154856 117098 154908 117104
rect 159088 117156 159140 117162
rect 159088 117098 159140 117104
rect 162032 117156 162084 117162
rect 162032 117098 162084 117104
rect 164332 117156 164384 117162
rect 164332 117098 164384 117104
rect 168196 117156 168248 117162
rect 168196 117098 168248 117104
rect 171232 117156 171284 117162
rect 171232 117098 171284 117104
rect 172888 117156 172940 117162
rect 172888 117098 172940 117104
rect 176016 117156 176068 117162
rect 176016 117098 176068 117104
rect 176936 117156 176988 117162
rect 176936 117098 176988 117104
rect 97632 117088 97684 117094
rect 97632 117030 97684 117036
rect 97644 116686 97672 117030
rect 97632 116680 97684 116686
rect 97632 116622 97684 116628
rect 96380 116444 96676 116464
rect 96436 116442 96460 116444
rect 96516 116442 96540 116444
rect 96596 116442 96620 116444
rect 96458 116390 96460 116442
rect 96522 116390 96534 116442
rect 96596 116390 96598 116442
rect 96436 116388 96460 116390
rect 96516 116388 96540 116390
rect 96596 116388 96620 116390
rect 96380 116368 96676 116388
rect 101232 116346 101260 117098
rect 103072 116754 103100 117098
rect 103060 116748 103112 116754
rect 103060 116690 103112 116696
rect 105372 116346 105400 117098
rect 107212 116822 107240 117098
rect 107200 116816 107252 116822
rect 107200 116758 107252 116764
rect 110248 116346 110276 117098
rect 111168 116890 111196 117098
rect 111740 116988 112036 117008
rect 111796 116986 111820 116988
rect 111876 116986 111900 116988
rect 111956 116986 111980 116988
rect 111818 116934 111820 116986
rect 111882 116934 111894 116986
rect 111956 116934 111958 116986
rect 111796 116932 111820 116934
rect 111876 116932 111900 116934
rect 111956 116932 111980 116934
rect 111740 116912 112036 116932
rect 111156 116884 111208 116890
rect 111156 116826 111208 116832
rect 114940 116346 114968 117098
rect 81808 116340 81860 116346
rect 81808 116282 81860 116288
rect 86592 116340 86644 116346
rect 86592 116282 86644 116288
rect 91376 116340 91428 116346
rect 91376 116282 91428 116288
rect 96068 116340 96120 116346
rect 96068 116282 96120 116288
rect 101220 116340 101272 116346
rect 101220 116282 101272 116288
rect 105360 116340 105412 116346
rect 105360 116282 105412 116288
rect 110236 116340 110288 116346
rect 110236 116282 110288 116288
rect 114928 116340 114980 116346
rect 114928 116282 114980 116288
rect 79048 116272 79100 116278
rect 79048 116214 79100 116220
rect 116688 116074 116716 117098
rect 119632 116346 119660 117098
rect 119620 116340 119672 116346
rect 119620 116282 119672 116288
rect 116676 116068 116728 116074
rect 116676 116010 116728 116016
rect 81020 115900 81316 115920
rect 81076 115898 81100 115900
rect 81156 115898 81180 115900
rect 81236 115898 81260 115900
rect 81098 115846 81100 115898
rect 81162 115846 81174 115898
rect 81236 115846 81238 115898
rect 81076 115844 81100 115846
rect 81156 115844 81180 115846
rect 81236 115844 81260 115846
rect 81020 115824 81316 115844
rect 111740 115900 112036 115920
rect 111796 115898 111820 115900
rect 111876 115898 111900 115900
rect 111956 115898 111980 115900
rect 111818 115846 111820 115898
rect 111882 115846 111894 115898
rect 111956 115846 111958 115898
rect 111796 115844 111820 115846
rect 111876 115844 111900 115846
rect 111956 115844 111980 115846
rect 111740 115824 112036 115844
rect 96380 115356 96676 115376
rect 96436 115354 96460 115356
rect 96516 115354 96540 115356
rect 96596 115354 96620 115356
rect 96458 115302 96460 115354
rect 96522 115302 96534 115354
rect 96596 115302 96598 115354
rect 96436 115300 96460 115302
rect 96516 115300 96540 115302
rect 96596 115300 96620 115302
rect 96380 115280 96676 115300
rect 81020 114812 81316 114832
rect 81076 114810 81100 114812
rect 81156 114810 81180 114812
rect 81236 114810 81260 114812
rect 81098 114758 81100 114810
rect 81162 114758 81174 114810
rect 81236 114758 81238 114810
rect 81076 114756 81100 114758
rect 81156 114756 81180 114758
rect 81236 114756 81260 114758
rect 81020 114736 81316 114756
rect 111740 114812 112036 114832
rect 111796 114810 111820 114812
rect 111876 114810 111900 114812
rect 111956 114810 111980 114812
rect 111818 114758 111820 114810
rect 111882 114758 111894 114810
rect 111956 114758 111958 114810
rect 111796 114756 111820 114758
rect 111876 114756 111900 114758
rect 111956 114756 111980 114758
rect 111740 114736 112036 114756
rect 96380 114268 96676 114288
rect 96436 114266 96460 114268
rect 96516 114266 96540 114268
rect 96596 114266 96620 114268
rect 96458 114214 96460 114266
rect 96522 114214 96534 114266
rect 96596 114214 96598 114266
rect 96436 114212 96460 114214
rect 96516 114212 96540 114214
rect 96596 114212 96620 114214
rect 96380 114192 96676 114212
rect 81020 113724 81316 113744
rect 81076 113722 81100 113724
rect 81156 113722 81180 113724
rect 81236 113722 81260 113724
rect 81098 113670 81100 113722
rect 81162 113670 81174 113722
rect 81236 113670 81238 113722
rect 81076 113668 81100 113670
rect 81156 113668 81180 113670
rect 81236 113668 81260 113670
rect 81020 113648 81316 113668
rect 111740 113724 112036 113744
rect 111796 113722 111820 113724
rect 111876 113722 111900 113724
rect 111956 113722 111980 113724
rect 111818 113670 111820 113722
rect 111882 113670 111894 113722
rect 111956 113670 111958 113722
rect 111796 113668 111820 113670
rect 111876 113668 111900 113670
rect 111956 113668 111980 113670
rect 111740 113648 112036 113668
rect 96380 113180 96676 113200
rect 96436 113178 96460 113180
rect 96516 113178 96540 113180
rect 96596 113178 96620 113180
rect 96458 113126 96460 113178
rect 96522 113126 96534 113178
rect 96596 113126 96598 113178
rect 96436 113124 96460 113126
rect 96516 113124 96540 113126
rect 96596 113124 96620 113126
rect 96380 113104 96676 113124
rect 81020 112636 81316 112656
rect 81076 112634 81100 112636
rect 81156 112634 81180 112636
rect 81236 112634 81260 112636
rect 81098 112582 81100 112634
rect 81162 112582 81174 112634
rect 81236 112582 81238 112634
rect 81076 112580 81100 112582
rect 81156 112580 81180 112582
rect 81236 112580 81260 112582
rect 81020 112560 81316 112580
rect 111740 112636 112036 112656
rect 111796 112634 111820 112636
rect 111876 112634 111900 112636
rect 111956 112634 111980 112636
rect 111818 112582 111820 112634
rect 111882 112582 111894 112634
rect 111956 112582 111958 112634
rect 111796 112580 111820 112582
rect 111876 112580 111900 112582
rect 111956 112580 111980 112582
rect 111740 112560 112036 112580
rect 96380 112092 96676 112112
rect 96436 112090 96460 112092
rect 96516 112090 96540 112092
rect 96596 112090 96620 112092
rect 96458 112038 96460 112090
rect 96522 112038 96534 112090
rect 96596 112038 96598 112090
rect 96436 112036 96460 112038
rect 96516 112036 96540 112038
rect 96596 112036 96620 112038
rect 96380 112016 96676 112036
rect 81020 111548 81316 111568
rect 81076 111546 81100 111548
rect 81156 111546 81180 111548
rect 81236 111546 81260 111548
rect 81098 111494 81100 111546
rect 81162 111494 81174 111546
rect 81236 111494 81238 111546
rect 81076 111492 81100 111494
rect 81156 111492 81180 111494
rect 81236 111492 81260 111494
rect 81020 111472 81316 111492
rect 111740 111548 112036 111568
rect 111796 111546 111820 111548
rect 111876 111546 111900 111548
rect 111956 111546 111980 111548
rect 111818 111494 111820 111546
rect 111882 111494 111894 111546
rect 111956 111494 111958 111546
rect 111796 111492 111820 111494
rect 111876 111492 111900 111494
rect 111956 111492 111980 111494
rect 111740 111472 112036 111492
rect 96380 111004 96676 111024
rect 96436 111002 96460 111004
rect 96516 111002 96540 111004
rect 96596 111002 96620 111004
rect 96458 110950 96460 111002
rect 96522 110950 96534 111002
rect 96596 110950 96598 111002
rect 96436 110948 96460 110950
rect 96516 110948 96540 110950
rect 96596 110948 96620 110950
rect 96380 110928 96676 110948
rect 81020 110460 81316 110480
rect 81076 110458 81100 110460
rect 81156 110458 81180 110460
rect 81236 110458 81260 110460
rect 81098 110406 81100 110458
rect 81162 110406 81174 110458
rect 81236 110406 81238 110458
rect 81076 110404 81100 110406
rect 81156 110404 81180 110406
rect 81236 110404 81260 110406
rect 81020 110384 81316 110404
rect 111740 110460 112036 110480
rect 111796 110458 111820 110460
rect 111876 110458 111900 110460
rect 111956 110458 111980 110460
rect 111818 110406 111820 110458
rect 111882 110406 111894 110458
rect 111956 110406 111958 110458
rect 111796 110404 111820 110406
rect 111876 110404 111900 110406
rect 111956 110404 111980 110406
rect 111740 110384 112036 110404
rect 96380 109916 96676 109936
rect 96436 109914 96460 109916
rect 96516 109914 96540 109916
rect 96596 109914 96620 109916
rect 96458 109862 96460 109914
rect 96522 109862 96534 109914
rect 96596 109862 96598 109914
rect 96436 109860 96460 109862
rect 96516 109860 96540 109862
rect 96596 109860 96620 109862
rect 96380 109840 96676 109860
rect 81020 109372 81316 109392
rect 81076 109370 81100 109372
rect 81156 109370 81180 109372
rect 81236 109370 81260 109372
rect 81098 109318 81100 109370
rect 81162 109318 81174 109370
rect 81236 109318 81238 109370
rect 81076 109316 81100 109318
rect 81156 109316 81180 109318
rect 81236 109316 81260 109318
rect 81020 109296 81316 109316
rect 111740 109372 112036 109392
rect 111796 109370 111820 109372
rect 111876 109370 111900 109372
rect 111956 109370 111980 109372
rect 111818 109318 111820 109370
rect 111882 109318 111894 109370
rect 111956 109318 111958 109370
rect 111796 109316 111820 109318
rect 111876 109316 111900 109318
rect 111956 109316 111980 109318
rect 111740 109296 112036 109316
rect 96380 108828 96676 108848
rect 96436 108826 96460 108828
rect 96516 108826 96540 108828
rect 96596 108826 96620 108828
rect 96458 108774 96460 108826
rect 96522 108774 96534 108826
rect 96596 108774 96598 108826
rect 96436 108772 96460 108774
rect 96516 108772 96540 108774
rect 96596 108772 96620 108774
rect 96380 108752 96676 108772
rect 81020 108284 81316 108304
rect 81076 108282 81100 108284
rect 81156 108282 81180 108284
rect 81236 108282 81260 108284
rect 81098 108230 81100 108282
rect 81162 108230 81174 108282
rect 81236 108230 81238 108282
rect 81076 108228 81100 108230
rect 81156 108228 81180 108230
rect 81236 108228 81260 108230
rect 81020 108208 81316 108228
rect 111740 108284 112036 108304
rect 111796 108282 111820 108284
rect 111876 108282 111900 108284
rect 111956 108282 111980 108284
rect 111818 108230 111820 108282
rect 111882 108230 111894 108282
rect 111956 108230 111958 108282
rect 111796 108228 111820 108230
rect 111876 108228 111900 108230
rect 111956 108228 111980 108230
rect 111740 108208 112036 108228
rect 96380 107740 96676 107760
rect 96436 107738 96460 107740
rect 96516 107738 96540 107740
rect 96596 107738 96620 107740
rect 96458 107686 96460 107738
rect 96522 107686 96534 107738
rect 96596 107686 96598 107738
rect 96436 107684 96460 107686
rect 96516 107684 96540 107686
rect 96596 107684 96620 107686
rect 96380 107664 96676 107684
rect 81020 107196 81316 107216
rect 81076 107194 81100 107196
rect 81156 107194 81180 107196
rect 81236 107194 81260 107196
rect 81098 107142 81100 107194
rect 81162 107142 81174 107194
rect 81236 107142 81238 107194
rect 81076 107140 81100 107142
rect 81156 107140 81180 107142
rect 81236 107140 81260 107142
rect 81020 107120 81316 107140
rect 111740 107196 112036 107216
rect 111796 107194 111820 107196
rect 111876 107194 111900 107196
rect 111956 107194 111980 107196
rect 111818 107142 111820 107194
rect 111882 107142 111894 107194
rect 111956 107142 111958 107194
rect 111796 107140 111820 107142
rect 111876 107140 111900 107142
rect 111956 107140 111980 107142
rect 111740 107120 112036 107140
rect 96380 106652 96676 106672
rect 96436 106650 96460 106652
rect 96516 106650 96540 106652
rect 96596 106650 96620 106652
rect 96458 106598 96460 106650
rect 96522 106598 96534 106650
rect 96596 106598 96598 106650
rect 96436 106596 96460 106598
rect 96516 106596 96540 106598
rect 96596 106596 96620 106598
rect 96380 106576 96676 106596
rect 81020 106108 81316 106128
rect 81076 106106 81100 106108
rect 81156 106106 81180 106108
rect 81236 106106 81260 106108
rect 81098 106054 81100 106106
rect 81162 106054 81174 106106
rect 81236 106054 81238 106106
rect 81076 106052 81100 106054
rect 81156 106052 81180 106054
rect 81236 106052 81260 106054
rect 81020 106032 81316 106052
rect 111740 106108 112036 106128
rect 111796 106106 111820 106108
rect 111876 106106 111900 106108
rect 111956 106106 111980 106108
rect 111818 106054 111820 106106
rect 111882 106054 111894 106106
rect 111956 106054 111958 106106
rect 111796 106052 111820 106054
rect 111876 106052 111900 106054
rect 111956 106052 111980 106054
rect 111740 106032 112036 106052
rect 96380 105564 96676 105584
rect 96436 105562 96460 105564
rect 96516 105562 96540 105564
rect 96596 105562 96620 105564
rect 96458 105510 96460 105562
rect 96522 105510 96534 105562
rect 96596 105510 96598 105562
rect 96436 105508 96460 105510
rect 96516 105508 96540 105510
rect 96596 105508 96620 105510
rect 96380 105488 96676 105508
rect 81020 105020 81316 105040
rect 81076 105018 81100 105020
rect 81156 105018 81180 105020
rect 81236 105018 81260 105020
rect 81098 104966 81100 105018
rect 81162 104966 81174 105018
rect 81236 104966 81238 105018
rect 81076 104964 81100 104966
rect 81156 104964 81180 104966
rect 81236 104964 81260 104966
rect 81020 104944 81316 104964
rect 111740 105020 112036 105040
rect 111796 105018 111820 105020
rect 111876 105018 111900 105020
rect 111956 105018 111980 105020
rect 111818 104966 111820 105018
rect 111882 104966 111894 105018
rect 111956 104966 111958 105018
rect 111796 104964 111820 104966
rect 111876 104964 111900 104966
rect 111956 104964 111980 104966
rect 111740 104944 112036 104964
rect 96380 104476 96676 104496
rect 96436 104474 96460 104476
rect 96516 104474 96540 104476
rect 96596 104474 96620 104476
rect 96458 104422 96460 104474
rect 96522 104422 96534 104474
rect 96596 104422 96598 104474
rect 96436 104420 96460 104422
rect 96516 104420 96540 104422
rect 96596 104420 96620 104422
rect 96380 104400 96676 104420
rect 81020 103932 81316 103952
rect 81076 103930 81100 103932
rect 81156 103930 81180 103932
rect 81236 103930 81260 103932
rect 81098 103878 81100 103930
rect 81162 103878 81174 103930
rect 81236 103878 81238 103930
rect 81076 103876 81100 103878
rect 81156 103876 81180 103878
rect 81236 103876 81260 103878
rect 81020 103856 81316 103876
rect 111740 103932 112036 103952
rect 111796 103930 111820 103932
rect 111876 103930 111900 103932
rect 111956 103930 111980 103932
rect 111818 103878 111820 103930
rect 111882 103878 111894 103930
rect 111956 103878 111958 103930
rect 111796 103876 111820 103878
rect 111876 103876 111900 103878
rect 111956 103876 111980 103878
rect 111740 103856 112036 103876
rect 96380 103388 96676 103408
rect 96436 103386 96460 103388
rect 96516 103386 96540 103388
rect 96596 103386 96620 103388
rect 96458 103334 96460 103386
rect 96522 103334 96534 103386
rect 96596 103334 96598 103386
rect 96436 103332 96460 103334
rect 96516 103332 96540 103334
rect 96596 103332 96620 103334
rect 96380 103312 96676 103332
rect 81020 102844 81316 102864
rect 81076 102842 81100 102844
rect 81156 102842 81180 102844
rect 81236 102842 81260 102844
rect 81098 102790 81100 102842
rect 81162 102790 81174 102842
rect 81236 102790 81238 102842
rect 81076 102788 81100 102790
rect 81156 102788 81180 102790
rect 81236 102788 81260 102790
rect 81020 102768 81316 102788
rect 111740 102844 112036 102864
rect 111796 102842 111820 102844
rect 111876 102842 111900 102844
rect 111956 102842 111980 102844
rect 111818 102790 111820 102842
rect 111882 102790 111894 102842
rect 111956 102790 111958 102842
rect 111796 102788 111820 102790
rect 111876 102788 111900 102790
rect 111956 102788 111980 102790
rect 111740 102768 112036 102788
rect 96380 102300 96676 102320
rect 96436 102298 96460 102300
rect 96516 102298 96540 102300
rect 96596 102298 96620 102300
rect 96458 102246 96460 102298
rect 96522 102246 96534 102298
rect 96596 102246 96598 102298
rect 96436 102244 96460 102246
rect 96516 102244 96540 102246
rect 96596 102244 96620 102246
rect 96380 102224 96676 102244
rect 81020 101756 81316 101776
rect 81076 101754 81100 101756
rect 81156 101754 81180 101756
rect 81236 101754 81260 101756
rect 81098 101702 81100 101754
rect 81162 101702 81174 101754
rect 81236 101702 81238 101754
rect 81076 101700 81100 101702
rect 81156 101700 81180 101702
rect 81236 101700 81260 101702
rect 81020 101680 81316 101700
rect 111740 101756 112036 101776
rect 111796 101754 111820 101756
rect 111876 101754 111900 101756
rect 111956 101754 111980 101756
rect 111818 101702 111820 101754
rect 111882 101702 111894 101754
rect 111956 101702 111958 101754
rect 111796 101700 111820 101702
rect 111876 101700 111900 101702
rect 111956 101700 111980 101702
rect 111740 101680 112036 101700
rect 96380 101212 96676 101232
rect 96436 101210 96460 101212
rect 96516 101210 96540 101212
rect 96596 101210 96620 101212
rect 96458 101158 96460 101210
rect 96522 101158 96534 101210
rect 96596 101158 96598 101210
rect 96436 101156 96460 101158
rect 96516 101156 96540 101158
rect 96596 101156 96620 101158
rect 96380 101136 96676 101156
rect 81020 100668 81316 100688
rect 81076 100666 81100 100668
rect 81156 100666 81180 100668
rect 81236 100666 81260 100668
rect 81098 100614 81100 100666
rect 81162 100614 81174 100666
rect 81236 100614 81238 100666
rect 81076 100612 81100 100614
rect 81156 100612 81180 100614
rect 81236 100612 81260 100614
rect 81020 100592 81316 100612
rect 111740 100668 112036 100688
rect 111796 100666 111820 100668
rect 111876 100666 111900 100668
rect 111956 100666 111980 100668
rect 111818 100614 111820 100666
rect 111882 100614 111894 100666
rect 111956 100614 111958 100666
rect 111796 100612 111820 100614
rect 111876 100612 111900 100614
rect 111956 100612 111980 100614
rect 111740 100592 112036 100612
rect 96380 100124 96676 100144
rect 96436 100122 96460 100124
rect 96516 100122 96540 100124
rect 96596 100122 96620 100124
rect 96458 100070 96460 100122
rect 96522 100070 96534 100122
rect 96596 100070 96598 100122
rect 96436 100068 96460 100070
rect 96516 100068 96540 100070
rect 96596 100068 96620 100070
rect 96380 100048 96676 100068
rect 81020 99580 81316 99600
rect 81076 99578 81100 99580
rect 81156 99578 81180 99580
rect 81236 99578 81260 99580
rect 81098 99526 81100 99578
rect 81162 99526 81174 99578
rect 81236 99526 81238 99578
rect 81076 99524 81100 99526
rect 81156 99524 81180 99526
rect 81236 99524 81260 99526
rect 81020 99504 81316 99524
rect 111740 99580 112036 99600
rect 111796 99578 111820 99580
rect 111876 99578 111900 99580
rect 111956 99578 111980 99580
rect 111818 99526 111820 99578
rect 111882 99526 111894 99578
rect 111956 99526 111958 99578
rect 111796 99524 111820 99526
rect 111876 99524 111900 99526
rect 111956 99524 111980 99526
rect 111740 99504 112036 99524
rect 96380 99036 96676 99056
rect 96436 99034 96460 99036
rect 96516 99034 96540 99036
rect 96596 99034 96620 99036
rect 96458 98982 96460 99034
rect 96522 98982 96534 99034
rect 96596 98982 96598 99034
rect 96436 98980 96460 98982
rect 96516 98980 96540 98982
rect 96596 98980 96620 98982
rect 96380 98960 96676 98980
rect 81020 98492 81316 98512
rect 81076 98490 81100 98492
rect 81156 98490 81180 98492
rect 81236 98490 81260 98492
rect 81098 98438 81100 98490
rect 81162 98438 81174 98490
rect 81236 98438 81238 98490
rect 81076 98436 81100 98438
rect 81156 98436 81180 98438
rect 81236 98436 81260 98438
rect 81020 98416 81316 98436
rect 111740 98492 112036 98512
rect 111796 98490 111820 98492
rect 111876 98490 111900 98492
rect 111956 98490 111980 98492
rect 111818 98438 111820 98490
rect 111882 98438 111894 98490
rect 111956 98438 111958 98490
rect 111796 98436 111820 98438
rect 111876 98436 111900 98438
rect 111956 98436 111980 98438
rect 111740 98416 112036 98436
rect 96380 97948 96676 97968
rect 96436 97946 96460 97948
rect 96516 97946 96540 97948
rect 96596 97946 96620 97948
rect 96458 97894 96460 97946
rect 96522 97894 96534 97946
rect 96596 97894 96598 97946
rect 96436 97892 96460 97894
rect 96516 97892 96540 97894
rect 96596 97892 96620 97894
rect 96380 97872 96676 97892
rect 81020 97404 81316 97424
rect 81076 97402 81100 97404
rect 81156 97402 81180 97404
rect 81236 97402 81260 97404
rect 81098 97350 81100 97402
rect 81162 97350 81174 97402
rect 81236 97350 81238 97402
rect 81076 97348 81100 97350
rect 81156 97348 81180 97350
rect 81236 97348 81260 97350
rect 81020 97328 81316 97348
rect 111740 97404 112036 97424
rect 111796 97402 111820 97404
rect 111876 97402 111900 97404
rect 111956 97402 111980 97404
rect 111818 97350 111820 97402
rect 111882 97350 111894 97402
rect 111956 97350 111958 97402
rect 111796 97348 111820 97350
rect 111876 97348 111900 97350
rect 111956 97348 111980 97350
rect 111740 97328 112036 97348
rect 96380 96860 96676 96880
rect 96436 96858 96460 96860
rect 96516 96858 96540 96860
rect 96596 96858 96620 96860
rect 96458 96806 96460 96858
rect 96522 96806 96534 96858
rect 96596 96806 96598 96858
rect 96436 96804 96460 96806
rect 96516 96804 96540 96806
rect 96596 96804 96620 96806
rect 96380 96784 96676 96804
rect 81020 96316 81316 96336
rect 81076 96314 81100 96316
rect 81156 96314 81180 96316
rect 81236 96314 81260 96316
rect 81098 96262 81100 96314
rect 81162 96262 81174 96314
rect 81236 96262 81238 96314
rect 81076 96260 81100 96262
rect 81156 96260 81180 96262
rect 81236 96260 81260 96262
rect 81020 96240 81316 96260
rect 111740 96316 112036 96336
rect 111796 96314 111820 96316
rect 111876 96314 111900 96316
rect 111956 96314 111980 96316
rect 111818 96262 111820 96314
rect 111882 96262 111894 96314
rect 111956 96262 111958 96314
rect 111796 96260 111820 96262
rect 111876 96260 111900 96262
rect 111956 96260 111980 96262
rect 111740 96240 112036 96260
rect 96380 95772 96676 95792
rect 96436 95770 96460 95772
rect 96516 95770 96540 95772
rect 96596 95770 96620 95772
rect 96458 95718 96460 95770
rect 96522 95718 96534 95770
rect 96596 95718 96598 95770
rect 96436 95716 96460 95718
rect 96516 95716 96540 95718
rect 96596 95716 96620 95718
rect 96380 95696 96676 95716
rect 81020 95228 81316 95248
rect 81076 95226 81100 95228
rect 81156 95226 81180 95228
rect 81236 95226 81260 95228
rect 81098 95174 81100 95226
rect 81162 95174 81174 95226
rect 81236 95174 81238 95226
rect 81076 95172 81100 95174
rect 81156 95172 81180 95174
rect 81236 95172 81260 95174
rect 81020 95152 81316 95172
rect 111740 95228 112036 95248
rect 111796 95226 111820 95228
rect 111876 95226 111900 95228
rect 111956 95226 111980 95228
rect 111818 95174 111820 95226
rect 111882 95174 111894 95226
rect 111956 95174 111958 95226
rect 111796 95172 111820 95174
rect 111876 95172 111900 95174
rect 111956 95172 111980 95174
rect 111740 95152 112036 95172
rect 96380 94684 96676 94704
rect 96436 94682 96460 94684
rect 96516 94682 96540 94684
rect 96596 94682 96620 94684
rect 96458 94630 96460 94682
rect 96522 94630 96534 94682
rect 96596 94630 96598 94682
rect 96436 94628 96460 94630
rect 96516 94628 96540 94630
rect 96596 94628 96620 94630
rect 96380 94608 96676 94628
rect 81020 94140 81316 94160
rect 81076 94138 81100 94140
rect 81156 94138 81180 94140
rect 81236 94138 81260 94140
rect 81098 94086 81100 94138
rect 81162 94086 81174 94138
rect 81236 94086 81238 94138
rect 81076 94084 81100 94086
rect 81156 94084 81180 94086
rect 81236 94084 81260 94086
rect 81020 94064 81316 94084
rect 111740 94140 112036 94160
rect 111796 94138 111820 94140
rect 111876 94138 111900 94140
rect 111956 94138 111980 94140
rect 111818 94086 111820 94138
rect 111882 94086 111894 94138
rect 111956 94086 111958 94138
rect 111796 94084 111820 94086
rect 111876 94084 111900 94086
rect 111956 94084 111980 94086
rect 111740 94064 112036 94084
rect 96380 93596 96676 93616
rect 96436 93594 96460 93596
rect 96516 93594 96540 93596
rect 96596 93594 96620 93596
rect 96458 93542 96460 93594
rect 96522 93542 96534 93594
rect 96596 93542 96598 93594
rect 96436 93540 96460 93542
rect 96516 93540 96540 93542
rect 96596 93540 96620 93542
rect 96380 93520 96676 93540
rect 81020 93052 81316 93072
rect 81076 93050 81100 93052
rect 81156 93050 81180 93052
rect 81236 93050 81260 93052
rect 81098 92998 81100 93050
rect 81162 92998 81174 93050
rect 81236 92998 81238 93050
rect 81076 92996 81100 92998
rect 81156 92996 81180 92998
rect 81236 92996 81260 92998
rect 81020 92976 81316 92996
rect 111740 93052 112036 93072
rect 111796 93050 111820 93052
rect 111876 93050 111900 93052
rect 111956 93050 111980 93052
rect 111818 92998 111820 93050
rect 111882 92998 111894 93050
rect 111956 92998 111958 93050
rect 111796 92996 111820 92998
rect 111876 92996 111900 92998
rect 111956 92996 111980 92998
rect 111740 92976 112036 92996
rect 96380 92508 96676 92528
rect 96436 92506 96460 92508
rect 96516 92506 96540 92508
rect 96596 92506 96620 92508
rect 96458 92454 96460 92506
rect 96522 92454 96534 92506
rect 96596 92454 96598 92506
rect 96436 92452 96460 92454
rect 96516 92452 96540 92454
rect 96596 92452 96620 92454
rect 96380 92432 96676 92452
rect 81020 91964 81316 91984
rect 81076 91962 81100 91964
rect 81156 91962 81180 91964
rect 81236 91962 81260 91964
rect 81098 91910 81100 91962
rect 81162 91910 81174 91962
rect 81236 91910 81238 91962
rect 81076 91908 81100 91910
rect 81156 91908 81180 91910
rect 81236 91908 81260 91910
rect 81020 91888 81316 91908
rect 111740 91964 112036 91984
rect 111796 91962 111820 91964
rect 111876 91962 111900 91964
rect 111956 91962 111980 91964
rect 111818 91910 111820 91962
rect 111882 91910 111894 91962
rect 111956 91910 111958 91962
rect 111796 91908 111820 91910
rect 111876 91908 111900 91910
rect 111956 91908 111980 91910
rect 111740 91888 112036 91908
rect 96380 91420 96676 91440
rect 96436 91418 96460 91420
rect 96516 91418 96540 91420
rect 96596 91418 96620 91420
rect 96458 91366 96460 91418
rect 96522 91366 96534 91418
rect 96596 91366 96598 91418
rect 96436 91364 96460 91366
rect 96516 91364 96540 91366
rect 96596 91364 96620 91366
rect 96380 91344 96676 91364
rect 81020 90876 81316 90896
rect 81076 90874 81100 90876
rect 81156 90874 81180 90876
rect 81236 90874 81260 90876
rect 81098 90822 81100 90874
rect 81162 90822 81174 90874
rect 81236 90822 81238 90874
rect 81076 90820 81100 90822
rect 81156 90820 81180 90822
rect 81236 90820 81260 90822
rect 81020 90800 81316 90820
rect 111740 90876 112036 90896
rect 111796 90874 111820 90876
rect 111876 90874 111900 90876
rect 111956 90874 111980 90876
rect 111818 90822 111820 90874
rect 111882 90822 111894 90874
rect 111956 90822 111958 90874
rect 111796 90820 111820 90822
rect 111876 90820 111900 90822
rect 111956 90820 111980 90822
rect 111740 90800 112036 90820
rect 96380 90332 96676 90352
rect 96436 90330 96460 90332
rect 96516 90330 96540 90332
rect 96596 90330 96620 90332
rect 96458 90278 96460 90330
rect 96522 90278 96534 90330
rect 96596 90278 96598 90330
rect 96436 90276 96460 90278
rect 96516 90276 96540 90278
rect 96596 90276 96620 90278
rect 96380 90256 96676 90276
rect 81020 89788 81316 89808
rect 81076 89786 81100 89788
rect 81156 89786 81180 89788
rect 81236 89786 81260 89788
rect 81098 89734 81100 89786
rect 81162 89734 81174 89786
rect 81236 89734 81238 89786
rect 81076 89732 81100 89734
rect 81156 89732 81180 89734
rect 81236 89732 81260 89734
rect 81020 89712 81316 89732
rect 111740 89788 112036 89808
rect 111796 89786 111820 89788
rect 111876 89786 111900 89788
rect 111956 89786 111980 89788
rect 111818 89734 111820 89786
rect 111882 89734 111894 89786
rect 111956 89734 111958 89786
rect 111796 89732 111820 89734
rect 111876 89732 111900 89734
rect 111956 89732 111980 89734
rect 111740 89712 112036 89732
rect 96380 89244 96676 89264
rect 96436 89242 96460 89244
rect 96516 89242 96540 89244
rect 96596 89242 96620 89244
rect 96458 89190 96460 89242
rect 96522 89190 96534 89242
rect 96596 89190 96598 89242
rect 96436 89188 96460 89190
rect 96516 89188 96540 89190
rect 96596 89188 96620 89190
rect 96380 89168 96676 89188
rect 81020 88700 81316 88720
rect 81076 88698 81100 88700
rect 81156 88698 81180 88700
rect 81236 88698 81260 88700
rect 81098 88646 81100 88698
rect 81162 88646 81174 88698
rect 81236 88646 81238 88698
rect 81076 88644 81100 88646
rect 81156 88644 81180 88646
rect 81236 88644 81260 88646
rect 81020 88624 81316 88644
rect 111740 88700 112036 88720
rect 111796 88698 111820 88700
rect 111876 88698 111900 88700
rect 111956 88698 111980 88700
rect 111818 88646 111820 88698
rect 111882 88646 111894 88698
rect 111956 88646 111958 88698
rect 111796 88644 111820 88646
rect 111876 88644 111900 88646
rect 111956 88644 111980 88646
rect 111740 88624 112036 88644
rect 96380 88156 96676 88176
rect 96436 88154 96460 88156
rect 96516 88154 96540 88156
rect 96596 88154 96620 88156
rect 96458 88102 96460 88154
rect 96522 88102 96534 88154
rect 96596 88102 96598 88154
rect 96436 88100 96460 88102
rect 96516 88100 96540 88102
rect 96596 88100 96620 88102
rect 96380 88080 96676 88100
rect 81020 87612 81316 87632
rect 81076 87610 81100 87612
rect 81156 87610 81180 87612
rect 81236 87610 81260 87612
rect 81098 87558 81100 87610
rect 81162 87558 81174 87610
rect 81236 87558 81238 87610
rect 81076 87556 81100 87558
rect 81156 87556 81180 87558
rect 81236 87556 81260 87558
rect 81020 87536 81316 87556
rect 111740 87612 112036 87632
rect 111796 87610 111820 87612
rect 111876 87610 111900 87612
rect 111956 87610 111980 87612
rect 111818 87558 111820 87610
rect 111882 87558 111894 87610
rect 111956 87558 111958 87610
rect 111796 87556 111820 87558
rect 111876 87556 111900 87558
rect 111956 87556 111980 87558
rect 111740 87536 112036 87556
rect 96380 87068 96676 87088
rect 96436 87066 96460 87068
rect 96516 87066 96540 87068
rect 96596 87066 96620 87068
rect 96458 87014 96460 87066
rect 96522 87014 96534 87066
rect 96596 87014 96598 87066
rect 96436 87012 96460 87014
rect 96516 87012 96540 87014
rect 96596 87012 96620 87014
rect 96380 86992 96676 87012
rect 81020 86524 81316 86544
rect 81076 86522 81100 86524
rect 81156 86522 81180 86524
rect 81236 86522 81260 86524
rect 81098 86470 81100 86522
rect 81162 86470 81174 86522
rect 81236 86470 81238 86522
rect 81076 86468 81100 86470
rect 81156 86468 81180 86470
rect 81236 86468 81260 86470
rect 81020 86448 81316 86468
rect 111740 86524 112036 86544
rect 111796 86522 111820 86524
rect 111876 86522 111900 86524
rect 111956 86522 111980 86524
rect 111818 86470 111820 86522
rect 111882 86470 111894 86522
rect 111956 86470 111958 86522
rect 111796 86468 111820 86470
rect 111876 86468 111900 86470
rect 111956 86468 111980 86470
rect 111740 86448 112036 86468
rect 96380 85980 96676 86000
rect 96436 85978 96460 85980
rect 96516 85978 96540 85980
rect 96596 85978 96620 85980
rect 96458 85926 96460 85978
rect 96522 85926 96534 85978
rect 96596 85926 96598 85978
rect 96436 85924 96460 85926
rect 96516 85924 96540 85926
rect 96596 85924 96620 85926
rect 96380 85904 96676 85924
rect 81020 85436 81316 85456
rect 81076 85434 81100 85436
rect 81156 85434 81180 85436
rect 81236 85434 81260 85436
rect 81098 85382 81100 85434
rect 81162 85382 81174 85434
rect 81236 85382 81238 85434
rect 81076 85380 81100 85382
rect 81156 85380 81180 85382
rect 81236 85380 81260 85382
rect 81020 85360 81316 85380
rect 111740 85436 112036 85456
rect 111796 85434 111820 85436
rect 111876 85434 111900 85436
rect 111956 85434 111980 85436
rect 111818 85382 111820 85434
rect 111882 85382 111894 85434
rect 111956 85382 111958 85434
rect 111796 85380 111820 85382
rect 111876 85380 111900 85382
rect 111956 85380 111980 85382
rect 111740 85360 112036 85380
rect 96380 84892 96676 84912
rect 96436 84890 96460 84892
rect 96516 84890 96540 84892
rect 96596 84890 96620 84892
rect 96458 84838 96460 84890
rect 96522 84838 96534 84890
rect 96596 84838 96598 84890
rect 96436 84836 96460 84838
rect 96516 84836 96540 84838
rect 96596 84836 96620 84838
rect 96380 84816 96676 84836
rect 81020 84348 81316 84368
rect 81076 84346 81100 84348
rect 81156 84346 81180 84348
rect 81236 84346 81260 84348
rect 81098 84294 81100 84346
rect 81162 84294 81174 84346
rect 81236 84294 81238 84346
rect 81076 84292 81100 84294
rect 81156 84292 81180 84294
rect 81236 84292 81260 84294
rect 81020 84272 81316 84292
rect 111740 84348 112036 84368
rect 111796 84346 111820 84348
rect 111876 84346 111900 84348
rect 111956 84346 111980 84348
rect 111818 84294 111820 84346
rect 111882 84294 111894 84346
rect 111956 84294 111958 84346
rect 111796 84292 111820 84294
rect 111876 84292 111900 84294
rect 111956 84292 111980 84294
rect 111740 84272 112036 84292
rect 96380 83804 96676 83824
rect 96436 83802 96460 83804
rect 96516 83802 96540 83804
rect 96596 83802 96620 83804
rect 96458 83750 96460 83802
rect 96522 83750 96534 83802
rect 96596 83750 96598 83802
rect 96436 83748 96460 83750
rect 96516 83748 96540 83750
rect 96596 83748 96620 83750
rect 96380 83728 96676 83748
rect 81020 83260 81316 83280
rect 81076 83258 81100 83260
rect 81156 83258 81180 83260
rect 81236 83258 81260 83260
rect 81098 83206 81100 83258
rect 81162 83206 81174 83258
rect 81236 83206 81238 83258
rect 81076 83204 81100 83206
rect 81156 83204 81180 83206
rect 81236 83204 81260 83206
rect 81020 83184 81316 83204
rect 111740 83260 112036 83280
rect 111796 83258 111820 83260
rect 111876 83258 111900 83260
rect 111956 83258 111980 83260
rect 111818 83206 111820 83258
rect 111882 83206 111894 83258
rect 111956 83206 111958 83258
rect 111796 83204 111820 83206
rect 111876 83204 111900 83206
rect 111956 83204 111980 83206
rect 111740 83184 112036 83204
rect 96380 82716 96676 82736
rect 96436 82714 96460 82716
rect 96516 82714 96540 82716
rect 96596 82714 96620 82716
rect 96458 82662 96460 82714
rect 96522 82662 96534 82714
rect 96596 82662 96598 82714
rect 96436 82660 96460 82662
rect 96516 82660 96540 82662
rect 96596 82660 96620 82662
rect 96380 82640 96676 82660
rect 81020 82172 81316 82192
rect 81076 82170 81100 82172
rect 81156 82170 81180 82172
rect 81236 82170 81260 82172
rect 81098 82118 81100 82170
rect 81162 82118 81174 82170
rect 81236 82118 81238 82170
rect 81076 82116 81100 82118
rect 81156 82116 81180 82118
rect 81236 82116 81260 82118
rect 81020 82096 81316 82116
rect 111740 82172 112036 82192
rect 111796 82170 111820 82172
rect 111876 82170 111900 82172
rect 111956 82170 111980 82172
rect 111818 82118 111820 82170
rect 111882 82118 111894 82170
rect 111956 82118 111958 82170
rect 111796 82116 111820 82118
rect 111876 82116 111900 82118
rect 111956 82116 111980 82118
rect 111740 82096 112036 82116
rect 96380 81628 96676 81648
rect 96436 81626 96460 81628
rect 96516 81626 96540 81628
rect 96596 81626 96620 81628
rect 96458 81574 96460 81626
rect 96522 81574 96534 81626
rect 96596 81574 96598 81626
rect 96436 81572 96460 81574
rect 96516 81572 96540 81574
rect 96596 81572 96620 81574
rect 96380 81552 96676 81572
rect 81020 81084 81316 81104
rect 81076 81082 81100 81084
rect 81156 81082 81180 81084
rect 81236 81082 81260 81084
rect 81098 81030 81100 81082
rect 81162 81030 81174 81082
rect 81236 81030 81238 81082
rect 81076 81028 81100 81030
rect 81156 81028 81180 81030
rect 81236 81028 81260 81030
rect 81020 81008 81316 81028
rect 111740 81084 112036 81104
rect 111796 81082 111820 81084
rect 111876 81082 111900 81084
rect 111956 81082 111980 81084
rect 111818 81030 111820 81082
rect 111882 81030 111894 81082
rect 111956 81030 111958 81082
rect 111796 81028 111820 81030
rect 111876 81028 111900 81030
rect 111956 81028 111980 81030
rect 111740 81008 112036 81028
rect 96380 80540 96676 80560
rect 96436 80538 96460 80540
rect 96516 80538 96540 80540
rect 96596 80538 96620 80540
rect 96458 80486 96460 80538
rect 96522 80486 96534 80538
rect 96596 80486 96598 80538
rect 96436 80484 96460 80486
rect 96516 80484 96540 80486
rect 96596 80484 96620 80486
rect 96380 80464 96676 80484
rect 81020 79996 81316 80016
rect 81076 79994 81100 79996
rect 81156 79994 81180 79996
rect 81236 79994 81260 79996
rect 81098 79942 81100 79994
rect 81162 79942 81174 79994
rect 81236 79942 81238 79994
rect 81076 79940 81100 79942
rect 81156 79940 81180 79942
rect 81236 79940 81260 79942
rect 81020 79920 81316 79940
rect 111740 79996 112036 80016
rect 111796 79994 111820 79996
rect 111876 79994 111900 79996
rect 111956 79994 111980 79996
rect 111818 79942 111820 79994
rect 111882 79942 111894 79994
rect 111956 79942 111958 79994
rect 111796 79940 111820 79942
rect 111876 79940 111900 79942
rect 111956 79940 111980 79942
rect 111740 79920 112036 79940
rect 96380 79452 96676 79472
rect 96436 79450 96460 79452
rect 96516 79450 96540 79452
rect 96596 79450 96620 79452
rect 96458 79398 96460 79450
rect 96522 79398 96534 79450
rect 96596 79398 96598 79450
rect 96436 79396 96460 79398
rect 96516 79396 96540 79398
rect 96596 79396 96620 79398
rect 96380 79376 96676 79396
rect 81020 78908 81316 78928
rect 81076 78906 81100 78908
rect 81156 78906 81180 78908
rect 81236 78906 81260 78908
rect 81098 78854 81100 78906
rect 81162 78854 81174 78906
rect 81236 78854 81238 78906
rect 81076 78852 81100 78854
rect 81156 78852 81180 78854
rect 81236 78852 81260 78854
rect 81020 78832 81316 78852
rect 111740 78908 112036 78928
rect 111796 78906 111820 78908
rect 111876 78906 111900 78908
rect 111956 78906 111980 78908
rect 111818 78854 111820 78906
rect 111882 78854 111894 78906
rect 111956 78854 111958 78906
rect 111796 78852 111820 78854
rect 111876 78852 111900 78854
rect 111956 78852 111980 78854
rect 111740 78832 112036 78852
rect 96380 78364 96676 78384
rect 96436 78362 96460 78364
rect 96516 78362 96540 78364
rect 96596 78362 96620 78364
rect 96458 78310 96460 78362
rect 96522 78310 96534 78362
rect 96596 78310 96598 78362
rect 96436 78308 96460 78310
rect 96516 78308 96540 78310
rect 96596 78308 96620 78310
rect 96380 78288 96676 78308
rect 81020 77820 81316 77840
rect 81076 77818 81100 77820
rect 81156 77818 81180 77820
rect 81236 77818 81260 77820
rect 81098 77766 81100 77818
rect 81162 77766 81174 77818
rect 81236 77766 81238 77818
rect 81076 77764 81100 77766
rect 81156 77764 81180 77766
rect 81236 77764 81260 77766
rect 81020 77744 81316 77764
rect 111740 77820 112036 77840
rect 111796 77818 111820 77820
rect 111876 77818 111900 77820
rect 111956 77818 111980 77820
rect 111818 77766 111820 77818
rect 111882 77766 111894 77818
rect 111956 77766 111958 77818
rect 111796 77764 111820 77766
rect 111876 77764 111900 77766
rect 111956 77764 111980 77766
rect 111740 77744 112036 77764
rect 96380 77276 96676 77296
rect 96436 77274 96460 77276
rect 96516 77274 96540 77276
rect 96596 77274 96620 77276
rect 96458 77222 96460 77274
rect 96522 77222 96534 77274
rect 96596 77222 96598 77274
rect 96436 77220 96460 77222
rect 96516 77220 96540 77222
rect 96596 77220 96620 77222
rect 96380 77200 96676 77220
rect 81020 76732 81316 76752
rect 81076 76730 81100 76732
rect 81156 76730 81180 76732
rect 81236 76730 81260 76732
rect 81098 76678 81100 76730
rect 81162 76678 81174 76730
rect 81236 76678 81238 76730
rect 81076 76676 81100 76678
rect 81156 76676 81180 76678
rect 81236 76676 81260 76678
rect 81020 76656 81316 76676
rect 111740 76732 112036 76752
rect 111796 76730 111820 76732
rect 111876 76730 111900 76732
rect 111956 76730 111980 76732
rect 111818 76678 111820 76730
rect 111882 76678 111894 76730
rect 111956 76678 111958 76730
rect 111796 76676 111820 76678
rect 111876 76676 111900 76678
rect 111956 76676 111980 76678
rect 111740 76656 112036 76676
rect 96380 76188 96676 76208
rect 96436 76186 96460 76188
rect 96516 76186 96540 76188
rect 96596 76186 96620 76188
rect 96458 76134 96460 76186
rect 96522 76134 96534 76186
rect 96596 76134 96598 76186
rect 96436 76132 96460 76134
rect 96516 76132 96540 76134
rect 96596 76132 96620 76134
rect 96380 76112 96676 76132
rect 81020 75644 81316 75664
rect 81076 75642 81100 75644
rect 81156 75642 81180 75644
rect 81236 75642 81260 75644
rect 81098 75590 81100 75642
rect 81162 75590 81174 75642
rect 81236 75590 81238 75642
rect 81076 75588 81100 75590
rect 81156 75588 81180 75590
rect 81236 75588 81260 75590
rect 81020 75568 81316 75588
rect 111740 75644 112036 75664
rect 111796 75642 111820 75644
rect 111876 75642 111900 75644
rect 111956 75642 111980 75644
rect 111818 75590 111820 75642
rect 111882 75590 111894 75642
rect 111956 75590 111958 75642
rect 111796 75588 111820 75590
rect 111876 75588 111900 75590
rect 111956 75588 111980 75590
rect 111740 75568 112036 75588
rect 96380 75100 96676 75120
rect 96436 75098 96460 75100
rect 96516 75098 96540 75100
rect 96596 75098 96620 75100
rect 96458 75046 96460 75098
rect 96522 75046 96534 75098
rect 96596 75046 96598 75098
rect 96436 75044 96460 75046
rect 96516 75044 96540 75046
rect 96596 75044 96620 75046
rect 96380 75024 96676 75044
rect 81020 74556 81316 74576
rect 81076 74554 81100 74556
rect 81156 74554 81180 74556
rect 81236 74554 81260 74556
rect 81098 74502 81100 74554
rect 81162 74502 81174 74554
rect 81236 74502 81238 74554
rect 81076 74500 81100 74502
rect 81156 74500 81180 74502
rect 81236 74500 81260 74502
rect 81020 74480 81316 74500
rect 111740 74556 112036 74576
rect 111796 74554 111820 74556
rect 111876 74554 111900 74556
rect 111956 74554 111980 74556
rect 111818 74502 111820 74554
rect 111882 74502 111894 74554
rect 111956 74502 111958 74554
rect 111796 74500 111820 74502
rect 111876 74500 111900 74502
rect 111956 74500 111980 74502
rect 111740 74480 112036 74500
rect 96380 74012 96676 74032
rect 96436 74010 96460 74012
rect 96516 74010 96540 74012
rect 96596 74010 96620 74012
rect 96458 73958 96460 74010
rect 96522 73958 96534 74010
rect 96596 73958 96598 74010
rect 96436 73956 96460 73958
rect 96516 73956 96540 73958
rect 96596 73956 96620 73958
rect 96380 73936 96676 73956
rect 81020 73468 81316 73488
rect 81076 73466 81100 73468
rect 81156 73466 81180 73468
rect 81236 73466 81260 73468
rect 81098 73414 81100 73466
rect 81162 73414 81174 73466
rect 81236 73414 81238 73466
rect 81076 73412 81100 73414
rect 81156 73412 81180 73414
rect 81236 73412 81260 73414
rect 81020 73392 81316 73412
rect 111740 73468 112036 73488
rect 111796 73466 111820 73468
rect 111876 73466 111900 73468
rect 111956 73466 111980 73468
rect 111818 73414 111820 73466
rect 111882 73414 111894 73466
rect 111956 73414 111958 73466
rect 111796 73412 111820 73414
rect 111876 73412 111900 73414
rect 111956 73412 111980 73414
rect 111740 73392 112036 73412
rect 96380 72924 96676 72944
rect 96436 72922 96460 72924
rect 96516 72922 96540 72924
rect 96596 72922 96620 72924
rect 96458 72870 96460 72922
rect 96522 72870 96534 72922
rect 96596 72870 96598 72922
rect 96436 72868 96460 72870
rect 96516 72868 96540 72870
rect 96596 72868 96620 72870
rect 96380 72848 96676 72868
rect 81020 72380 81316 72400
rect 81076 72378 81100 72380
rect 81156 72378 81180 72380
rect 81236 72378 81260 72380
rect 81098 72326 81100 72378
rect 81162 72326 81174 72378
rect 81236 72326 81238 72378
rect 81076 72324 81100 72326
rect 81156 72324 81180 72326
rect 81236 72324 81260 72326
rect 81020 72304 81316 72324
rect 111740 72380 112036 72400
rect 111796 72378 111820 72380
rect 111876 72378 111900 72380
rect 111956 72378 111980 72380
rect 111818 72326 111820 72378
rect 111882 72326 111894 72378
rect 111956 72326 111958 72378
rect 111796 72324 111820 72326
rect 111876 72324 111900 72326
rect 111956 72324 111980 72326
rect 111740 72304 112036 72324
rect 96380 71836 96676 71856
rect 96436 71834 96460 71836
rect 96516 71834 96540 71836
rect 96596 71834 96620 71836
rect 96458 71782 96460 71834
rect 96522 71782 96534 71834
rect 96596 71782 96598 71834
rect 96436 71780 96460 71782
rect 96516 71780 96540 71782
rect 96596 71780 96620 71782
rect 96380 71760 96676 71780
rect 81020 71292 81316 71312
rect 81076 71290 81100 71292
rect 81156 71290 81180 71292
rect 81236 71290 81260 71292
rect 81098 71238 81100 71290
rect 81162 71238 81174 71290
rect 81236 71238 81238 71290
rect 81076 71236 81100 71238
rect 81156 71236 81180 71238
rect 81236 71236 81260 71238
rect 81020 71216 81316 71236
rect 111740 71292 112036 71312
rect 111796 71290 111820 71292
rect 111876 71290 111900 71292
rect 111956 71290 111980 71292
rect 111818 71238 111820 71290
rect 111882 71238 111894 71290
rect 111956 71238 111958 71290
rect 111796 71236 111820 71238
rect 111876 71236 111900 71238
rect 111956 71236 111980 71238
rect 111740 71216 112036 71236
rect 96380 70748 96676 70768
rect 96436 70746 96460 70748
rect 96516 70746 96540 70748
rect 96596 70746 96620 70748
rect 96458 70694 96460 70746
rect 96522 70694 96534 70746
rect 96596 70694 96598 70746
rect 96436 70692 96460 70694
rect 96516 70692 96540 70694
rect 96596 70692 96620 70694
rect 96380 70672 96676 70692
rect 81020 70204 81316 70224
rect 81076 70202 81100 70204
rect 81156 70202 81180 70204
rect 81236 70202 81260 70204
rect 81098 70150 81100 70202
rect 81162 70150 81174 70202
rect 81236 70150 81238 70202
rect 81076 70148 81100 70150
rect 81156 70148 81180 70150
rect 81236 70148 81260 70150
rect 81020 70128 81316 70148
rect 111740 70204 112036 70224
rect 111796 70202 111820 70204
rect 111876 70202 111900 70204
rect 111956 70202 111980 70204
rect 111818 70150 111820 70202
rect 111882 70150 111894 70202
rect 111956 70150 111958 70202
rect 111796 70148 111820 70150
rect 111876 70148 111900 70150
rect 111956 70148 111980 70150
rect 111740 70128 112036 70148
rect 96380 69660 96676 69680
rect 96436 69658 96460 69660
rect 96516 69658 96540 69660
rect 96596 69658 96620 69660
rect 96458 69606 96460 69658
rect 96522 69606 96534 69658
rect 96596 69606 96598 69658
rect 96436 69604 96460 69606
rect 96516 69604 96540 69606
rect 96596 69604 96620 69606
rect 96380 69584 96676 69604
rect 81020 69116 81316 69136
rect 81076 69114 81100 69116
rect 81156 69114 81180 69116
rect 81236 69114 81260 69116
rect 81098 69062 81100 69114
rect 81162 69062 81174 69114
rect 81236 69062 81238 69114
rect 81076 69060 81100 69062
rect 81156 69060 81180 69062
rect 81236 69060 81260 69062
rect 81020 69040 81316 69060
rect 111740 69116 112036 69136
rect 111796 69114 111820 69116
rect 111876 69114 111900 69116
rect 111956 69114 111980 69116
rect 111818 69062 111820 69114
rect 111882 69062 111894 69114
rect 111956 69062 111958 69114
rect 111796 69060 111820 69062
rect 111876 69060 111900 69062
rect 111956 69060 111980 69062
rect 111740 69040 112036 69060
rect 96380 68572 96676 68592
rect 96436 68570 96460 68572
rect 96516 68570 96540 68572
rect 96596 68570 96620 68572
rect 96458 68518 96460 68570
rect 96522 68518 96534 68570
rect 96596 68518 96598 68570
rect 96436 68516 96460 68518
rect 96516 68516 96540 68518
rect 96596 68516 96620 68518
rect 96380 68496 96676 68516
rect 81020 68028 81316 68048
rect 81076 68026 81100 68028
rect 81156 68026 81180 68028
rect 81236 68026 81260 68028
rect 81098 67974 81100 68026
rect 81162 67974 81174 68026
rect 81236 67974 81238 68026
rect 81076 67972 81100 67974
rect 81156 67972 81180 67974
rect 81236 67972 81260 67974
rect 81020 67952 81316 67972
rect 111740 68028 112036 68048
rect 111796 68026 111820 68028
rect 111876 68026 111900 68028
rect 111956 68026 111980 68028
rect 111818 67974 111820 68026
rect 111882 67974 111894 68026
rect 111956 67974 111958 68026
rect 111796 67972 111820 67974
rect 111876 67972 111900 67974
rect 111956 67972 111980 67974
rect 111740 67952 112036 67972
rect 96380 67484 96676 67504
rect 96436 67482 96460 67484
rect 96516 67482 96540 67484
rect 96596 67482 96620 67484
rect 96458 67430 96460 67482
rect 96522 67430 96534 67482
rect 96596 67430 96598 67482
rect 96436 67428 96460 67430
rect 96516 67428 96540 67430
rect 96596 67428 96620 67430
rect 96380 67408 96676 67428
rect 81020 66940 81316 66960
rect 81076 66938 81100 66940
rect 81156 66938 81180 66940
rect 81236 66938 81260 66940
rect 81098 66886 81100 66938
rect 81162 66886 81174 66938
rect 81236 66886 81238 66938
rect 81076 66884 81100 66886
rect 81156 66884 81180 66886
rect 81236 66884 81260 66886
rect 81020 66864 81316 66884
rect 111740 66940 112036 66960
rect 111796 66938 111820 66940
rect 111876 66938 111900 66940
rect 111956 66938 111980 66940
rect 111818 66886 111820 66938
rect 111882 66886 111894 66938
rect 111956 66886 111958 66938
rect 111796 66884 111820 66886
rect 111876 66884 111900 66886
rect 111956 66884 111980 66886
rect 111740 66864 112036 66884
rect 96380 66396 96676 66416
rect 96436 66394 96460 66396
rect 96516 66394 96540 66396
rect 96596 66394 96620 66396
rect 96458 66342 96460 66394
rect 96522 66342 96534 66394
rect 96596 66342 96598 66394
rect 96436 66340 96460 66342
rect 96516 66340 96540 66342
rect 96596 66340 96620 66342
rect 96380 66320 96676 66340
rect 81020 65852 81316 65872
rect 81076 65850 81100 65852
rect 81156 65850 81180 65852
rect 81236 65850 81260 65852
rect 81098 65798 81100 65850
rect 81162 65798 81174 65850
rect 81236 65798 81238 65850
rect 81076 65796 81100 65798
rect 81156 65796 81180 65798
rect 81236 65796 81260 65798
rect 81020 65776 81316 65796
rect 111740 65852 112036 65872
rect 111796 65850 111820 65852
rect 111876 65850 111900 65852
rect 111956 65850 111980 65852
rect 111818 65798 111820 65850
rect 111882 65798 111894 65850
rect 111956 65798 111958 65850
rect 111796 65796 111820 65798
rect 111876 65796 111900 65798
rect 111956 65796 111980 65798
rect 111740 65776 112036 65796
rect 96380 65308 96676 65328
rect 96436 65306 96460 65308
rect 96516 65306 96540 65308
rect 96596 65306 96620 65308
rect 96458 65254 96460 65306
rect 96522 65254 96534 65306
rect 96596 65254 96598 65306
rect 96436 65252 96460 65254
rect 96516 65252 96540 65254
rect 96596 65252 96620 65254
rect 96380 65232 96676 65252
rect 81020 64764 81316 64784
rect 81076 64762 81100 64764
rect 81156 64762 81180 64764
rect 81236 64762 81260 64764
rect 81098 64710 81100 64762
rect 81162 64710 81174 64762
rect 81236 64710 81238 64762
rect 81076 64708 81100 64710
rect 81156 64708 81180 64710
rect 81236 64708 81260 64710
rect 81020 64688 81316 64708
rect 111740 64764 112036 64784
rect 111796 64762 111820 64764
rect 111876 64762 111900 64764
rect 111956 64762 111980 64764
rect 111818 64710 111820 64762
rect 111882 64710 111894 64762
rect 111956 64710 111958 64762
rect 111796 64708 111820 64710
rect 111876 64708 111900 64710
rect 111956 64708 111980 64710
rect 111740 64688 112036 64708
rect 96380 64220 96676 64240
rect 96436 64218 96460 64220
rect 96516 64218 96540 64220
rect 96596 64218 96620 64220
rect 96458 64166 96460 64218
rect 96522 64166 96534 64218
rect 96596 64166 96598 64218
rect 96436 64164 96460 64166
rect 96516 64164 96540 64166
rect 96596 64164 96620 64166
rect 96380 64144 96676 64164
rect 81020 63676 81316 63696
rect 81076 63674 81100 63676
rect 81156 63674 81180 63676
rect 81236 63674 81260 63676
rect 81098 63622 81100 63674
rect 81162 63622 81174 63674
rect 81236 63622 81238 63674
rect 81076 63620 81100 63622
rect 81156 63620 81180 63622
rect 81236 63620 81260 63622
rect 81020 63600 81316 63620
rect 111740 63676 112036 63696
rect 111796 63674 111820 63676
rect 111876 63674 111900 63676
rect 111956 63674 111980 63676
rect 111818 63622 111820 63674
rect 111882 63622 111894 63674
rect 111956 63622 111958 63674
rect 111796 63620 111820 63622
rect 111876 63620 111900 63622
rect 111956 63620 111980 63622
rect 111740 63600 112036 63620
rect 96380 63132 96676 63152
rect 96436 63130 96460 63132
rect 96516 63130 96540 63132
rect 96596 63130 96620 63132
rect 96458 63078 96460 63130
rect 96522 63078 96534 63130
rect 96596 63078 96598 63130
rect 96436 63076 96460 63078
rect 96516 63076 96540 63078
rect 96596 63076 96620 63078
rect 96380 63056 96676 63076
rect 81020 62588 81316 62608
rect 81076 62586 81100 62588
rect 81156 62586 81180 62588
rect 81236 62586 81260 62588
rect 81098 62534 81100 62586
rect 81162 62534 81174 62586
rect 81236 62534 81238 62586
rect 81076 62532 81100 62534
rect 81156 62532 81180 62534
rect 81236 62532 81260 62534
rect 81020 62512 81316 62532
rect 111740 62588 112036 62608
rect 111796 62586 111820 62588
rect 111876 62586 111900 62588
rect 111956 62586 111980 62588
rect 111818 62534 111820 62586
rect 111882 62534 111894 62586
rect 111956 62534 111958 62586
rect 111796 62532 111820 62534
rect 111876 62532 111900 62534
rect 111956 62532 111980 62534
rect 111740 62512 112036 62532
rect 96380 62044 96676 62064
rect 96436 62042 96460 62044
rect 96516 62042 96540 62044
rect 96596 62042 96620 62044
rect 96458 61990 96460 62042
rect 96522 61990 96534 62042
rect 96596 61990 96598 62042
rect 96436 61988 96460 61990
rect 96516 61988 96540 61990
rect 96596 61988 96620 61990
rect 96380 61968 96676 61988
rect 81020 61500 81316 61520
rect 81076 61498 81100 61500
rect 81156 61498 81180 61500
rect 81236 61498 81260 61500
rect 81098 61446 81100 61498
rect 81162 61446 81174 61498
rect 81236 61446 81238 61498
rect 81076 61444 81100 61446
rect 81156 61444 81180 61446
rect 81236 61444 81260 61446
rect 81020 61424 81316 61444
rect 111740 61500 112036 61520
rect 111796 61498 111820 61500
rect 111876 61498 111900 61500
rect 111956 61498 111980 61500
rect 111818 61446 111820 61498
rect 111882 61446 111894 61498
rect 111956 61446 111958 61498
rect 111796 61444 111820 61446
rect 111876 61444 111900 61446
rect 111956 61444 111980 61446
rect 111740 61424 112036 61444
rect 96380 60956 96676 60976
rect 96436 60954 96460 60956
rect 96516 60954 96540 60956
rect 96596 60954 96620 60956
rect 96458 60902 96460 60954
rect 96522 60902 96534 60954
rect 96596 60902 96598 60954
rect 96436 60900 96460 60902
rect 96516 60900 96540 60902
rect 96596 60900 96620 60902
rect 96380 60880 96676 60900
rect 81020 60412 81316 60432
rect 81076 60410 81100 60412
rect 81156 60410 81180 60412
rect 81236 60410 81260 60412
rect 81098 60358 81100 60410
rect 81162 60358 81174 60410
rect 81236 60358 81238 60410
rect 81076 60356 81100 60358
rect 81156 60356 81180 60358
rect 81236 60356 81260 60358
rect 81020 60336 81316 60356
rect 111740 60412 112036 60432
rect 111796 60410 111820 60412
rect 111876 60410 111900 60412
rect 111956 60410 111980 60412
rect 111818 60358 111820 60410
rect 111882 60358 111894 60410
rect 111956 60358 111958 60410
rect 111796 60356 111820 60358
rect 111876 60356 111900 60358
rect 111956 60356 111980 60358
rect 111740 60336 112036 60356
rect 96380 59868 96676 59888
rect 96436 59866 96460 59868
rect 96516 59866 96540 59868
rect 96596 59866 96620 59868
rect 96458 59814 96460 59866
rect 96522 59814 96534 59866
rect 96596 59814 96598 59866
rect 96436 59812 96460 59814
rect 96516 59812 96540 59814
rect 96596 59812 96620 59814
rect 96380 59792 96676 59812
rect 81020 59324 81316 59344
rect 81076 59322 81100 59324
rect 81156 59322 81180 59324
rect 81236 59322 81260 59324
rect 81098 59270 81100 59322
rect 81162 59270 81174 59322
rect 81236 59270 81238 59322
rect 81076 59268 81100 59270
rect 81156 59268 81180 59270
rect 81236 59268 81260 59270
rect 81020 59248 81316 59268
rect 111740 59324 112036 59344
rect 111796 59322 111820 59324
rect 111876 59322 111900 59324
rect 111956 59322 111980 59324
rect 111818 59270 111820 59322
rect 111882 59270 111894 59322
rect 111956 59270 111958 59322
rect 111796 59268 111820 59270
rect 111876 59268 111900 59270
rect 111956 59268 111980 59270
rect 111740 59248 112036 59268
rect 96380 58780 96676 58800
rect 96436 58778 96460 58780
rect 96516 58778 96540 58780
rect 96596 58778 96620 58780
rect 96458 58726 96460 58778
rect 96522 58726 96534 58778
rect 96596 58726 96598 58778
rect 96436 58724 96460 58726
rect 96516 58724 96540 58726
rect 96596 58724 96620 58726
rect 96380 58704 96676 58724
rect 81020 58236 81316 58256
rect 81076 58234 81100 58236
rect 81156 58234 81180 58236
rect 81236 58234 81260 58236
rect 81098 58182 81100 58234
rect 81162 58182 81174 58234
rect 81236 58182 81238 58234
rect 81076 58180 81100 58182
rect 81156 58180 81180 58182
rect 81236 58180 81260 58182
rect 81020 58160 81316 58180
rect 111740 58236 112036 58256
rect 111796 58234 111820 58236
rect 111876 58234 111900 58236
rect 111956 58234 111980 58236
rect 111818 58182 111820 58234
rect 111882 58182 111894 58234
rect 111956 58182 111958 58234
rect 111796 58180 111820 58182
rect 111876 58180 111900 58182
rect 111956 58180 111980 58182
rect 111740 58160 112036 58180
rect 96380 57692 96676 57712
rect 96436 57690 96460 57692
rect 96516 57690 96540 57692
rect 96596 57690 96620 57692
rect 96458 57638 96460 57690
rect 96522 57638 96534 57690
rect 96596 57638 96598 57690
rect 96436 57636 96460 57638
rect 96516 57636 96540 57638
rect 96596 57636 96620 57638
rect 96380 57616 96676 57636
rect 81020 57148 81316 57168
rect 81076 57146 81100 57148
rect 81156 57146 81180 57148
rect 81236 57146 81260 57148
rect 81098 57094 81100 57146
rect 81162 57094 81174 57146
rect 81236 57094 81238 57146
rect 81076 57092 81100 57094
rect 81156 57092 81180 57094
rect 81236 57092 81260 57094
rect 81020 57072 81316 57092
rect 111740 57148 112036 57168
rect 111796 57146 111820 57148
rect 111876 57146 111900 57148
rect 111956 57146 111980 57148
rect 111818 57094 111820 57146
rect 111882 57094 111894 57146
rect 111956 57094 111958 57146
rect 111796 57092 111820 57094
rect 111876 57092 111900 57094
rect 111956 57092 111980 57094
rect 111740 57072 112036 57092
rect 96380 56604 96676 56624
rect 96436 56602 96460 56604
rect 96516 56602 96540 56604
rect 96596 56602 96620 56604
rect 96458 56550 96460 56602
rect 96522 56550 96534 56602
rect 96596 56550 96598 56602
rect 96436 56548 96460 56550
rect 96516 56548 96540 56550
rect 96596 56548 96620 56550
rect 96380 56528 96676 56548
rect 81020 56060 81316 56080
rect 81076 56058 81100 56060
rect 81156 56058 81180 56060
rect 81236 56058 81260 56060
rect 81098 56006 81100 56058
rect 81162 56006 81174 56058
rect 81236 56006 81238 56058
rect 81076 56004 81100 56006
rect 81156 56004 81180 56006
rect 81236 56004 81260 56006
rect 81020 55984 81316 56004
rect 111740 56060 112036 56080
rect 111796 56058 111820 56060
rect 111876 56058 111900 56060
rect 111956 56058 111980 56060
rect 111818 56006 111820 56058
rect 111882 56006 111894 56058
rect 111956 56006 111958 56058
rect 111796 56004 111820 56006
rect 111876 56004 111900 56006
rect 111956 56004 111980 56006
rect 111740 55984 112036 56004
rect 96380 55516 96676 55536
rect 96436 55514 96460 55516
rect 96516 55514 96540 55516
rect 96596 55514 96620 55516
rect 96458 55462 96460 55514
rect 96522 55462 96534 55514
rect 96596 55462 96598 55514
rect 96436 55460 96460 55462
rect 96516 55460 96540 55462
rect 96596 55460 96620 55462
rect 96380 55440 96676 55460
rect 81020 54972 81316 54992
rect 81076 54970 81100 54972
rect 81156 54970 81180 54972
rect 81236 54970 81260 54972
rect 81098 54918 81100 54970
rect 81162 54918 81174 54970
rect 81236 54918 81238 54970
rect 81076 54916 81100 54918
rect 81156 54916 81180 54918
rect 81236 54916 81260 54918
rect 81020 54896 81316 54916
rect 111740 54972 112036 54992
rect 111796 54970 111820 54972
rect 111876 54970 111900 54972
rect 111956 54970 111980 54972
rect 111818 54918 111820 54970
rect 111882 54918 111894 54970
rect 111956 54918 111958 54970
rect 111796 54916 111820 54918
rect 111876 54916 111900 54918
rect 111956 54916 111980 54918
rect 111740 54896 112036 54916
rect 96380 54428 96676 54448
rect 96436 54426 96460 54428
rect 96516 54426 96540 54428
rect 96596 54426 96620 54428
rect 96458 54374 96460 54426
rect 96522 54374 96534 54426
rect 96596 54374 96598 54426
rect 96436 54372 96460 54374
rect 96516 54372 96540 54374
rect 96596 54372 96620 54374
rect 96380 54352 96676 54372
rect 81020 53884 81316 53904
rect 81076 53882 81100 53884
rect 81156 53882 81180 53884
rect 81236 53882 81260 53884
rect 81098 53830 81100 53882
rect 81162 53830 81174 53882
rect 81236 53830 81238 53882
rect 81076 53828 81100 53830
rect 81156 53828 81180 53830
rect 81236 53828 81260 53830
rect 81020 53808 81316 53828
rect 111740 53884 112036 53904
rect 111796 53882 111820 53884
rect 111876 53882 111900 53884
rect 111956 53882 111980 53884
rect 111818 53830 111820 53882
rect 111882 53830 111894 53882
rect 111956 53830 111958 53882
rect 111796 53828 111820 53830
rect 111876 53828 111900 53830
rect 111956 53828 111980 53830
rect 111740 53808 112036 53828
rect 96380 53340 96676 53360
rect 96436 53338 96460 53340
rect 96516 53338 96540 53340
rect 96596 53338 96620 53340
rect 96458 53286 96460 53338
rect 96522 53286 96534 53338
rect 96596 53286 96598 53338
rect 96436 53284 96460 53286
rect 96516 53284 96540 53286
rect 96596 53284 96620 53286
rect 96380 53264 96676 53284
rect 81020 52796 81316 52816
rect 81076 52794 81100 52796
rect 81156 52794 81180 52796
rect 81236 52794 81260 52796
rect 81098 52742 81100 52794
rect 81162 52742 81174 52794
rect 81236 52742 81238 52794
rect 81076 52740 81100 52742
rect 81156 52740 81180 52742
rect 81236 52740 81260 52742
rect 81020 52720 81316 52740
rect 111740 52796 112036 52816
rect 111796 52794 111820 52796
rect 111876 52794 111900 52796
rect 111956 52794 111980 52796
rect 111818 52742 111820 52794
rect 111882 52742 111894 52794
rect 111956 52742 111958 52794
rect 111796 52740 111820 52742
rect 111876 52740 111900 52742
rect 111956 52740 111980 52742
rect 111740 52720 112036 52740
rect 96380 52252 96676 52272
rect 96436 52250 96460 52252
rect 96516 52250 96540 52252
rect 96596 52250 96620 52252
rect 96458 52198 96460 52250
rect 96522 52198 96534 52250
rect 96596 52198 96598 52250
rect 96436 52196 96460 52198
rect 96516 52196 96540 52198
rect 96596 52196 96620 52198
rect 96380 52176 96676 52196
rect 81020 51708 81316 51728
rect 81076 51706 81100 51708
rect 81156 51706 81180 51708
rect 81236 51706 81260 51708
rect 81098 51654 81100 51706
rect 81162 51654 81174 51706
rect 81236 51654 81238 51706
rect 81076 51652 81100 51654
rect 81156 51652 81180 51654
rect 81236 51652 81260 51654
rect 81020 51632 81316 51652
rect 111740 51708 112036 51728
rect 111796 51706 111820 51708
rect 111876 51706 111900 51708
rect 111956 51706 111980 51708
rect 111818 51654 111820 51706
rect 111882 51654 111894 51706
rect 111956 51654 111958 51706
rect 111796 51652 111820 51654
rect 111876 51652 111900 51654
rect 111956 51652 111980 51654
rect 111740 51632 112036 51652
rect 96380 51164 96676 51184
rect 96436 51162 96460 51164
rect 96516 51162 96540 51164
rect 96596 51162 96620 51164
rect 96458 51110 96460 51162
rect 96522 51110 96534 51162
rect 96596 51110 96598 51162
rect 96436 51108 96460 51110
rect 96516 51108 96540 51110
rect 96596 51108 96620 51110
rect 96380 51088 96676 51108
rect 81020 50620 81316 50640
rect 81076 50618 81100 50620
rect 81156 50618 81180 50620
rect 81236 50618 81260 50620
rect 81098 50566 81100 50618
rect 81162 50566 81174 50618
rect 81236 50566 81238 50618
rect 81076 50564 81100 50566
rect 81156 50564 81180 50566
rect 81236 50564 81260 50566
rect 81020 50544 81316 50564
rect 111740 50620 112036 50640
rect 111796 50618 111820 50620
rect 111876 50618 111900 50620
rect 111956 50618 111980 50620
rect 111818 50566 111820 50618
rect 111882 50566 111894 50618
rect 111956 50566 111958 50618
rect 111796 50564 111820 50566
rect 111876 50564 111900 50566
rect 111956 50564 111980 50566
rect 111740 50544 112036 50564
rect 96380 50076 96676 50096
rect 96436 50074 96460 50076
rect 96516 50074 96540 50076
rect 96596 50074 96620 50076
rect 96458 50022 96460 50074
rect 96522 50022 96534 50074
rect 96596 50022 96598 50074
rect 96436 50020 96460 50022
rect 96516 50020 96540 50022
rect 96596 50020 96620 50022
rect 96380 50000 96676 50020
rect 81020 49532 81316 49552
rect 81076 49530 81100 49532
rect 81156 49530 81180 49532
rect 81236 49530 81260 49532
rect 81098 49478 81100 49530
rect 81162 49478 81174 49530
rect 81236 49478 81238 49530
rect 81076 49476 81100 49478
rect 81156 49476 81180 49478
rect 81236 49476 81260 49478
rect 81020 49456 81316 49476
rect 111740 49532 112036 49552
rect 111796 49530 111820 49532
rect 111876 49530 111900 49532
rect 111956 49530 111980 49532
rect 111818 49478 111820 49530
rect 111882 49478 111894 49530
rect 111956 49478 111958 49530
rect 111796 49476 111820 49478
rect 111876 49476 111900 49478
rect 111956 49476 111980 49478
rect 111740 49456 112036 49476
rect 96380 48988 96676 49008
rect 96436 48986 96460 48988
rect 96516 48986 96540 48988
rect 96596 48986 96620 48988
rect 96458 48934 96460 48986
rect 96522 48934 96534 48986
rect 96596 48934 96598 48986
rect 96436 48932 96460 48934
rect 96516 48932 96540 48934
rect 96596 48932 96620 48934
rect 96380 48912 96676 48932
rect 81020 48444 81316 48464
rect 81076 48442 81100 48444
rect 81156 48442 81180 48444
rect 81236 48442 81260 48444
rect 81098 48390 81100 48442
rect 81162 48390 81174 48442
rect 81236 48390 81238 48442
rect 81076 48388 81100 48390
rect 81156 48388 81180 48390
rect 81236 48388 81260 48390
rect 81020 48368 81316 48388
rect 111740 48444 112036 48464
rect 111796 48442 111820 48444
rect 111876 48442 111900 48444
rect 111956 48442 111980 48444
rect 111818 48390 111820 48442
rect 111882 48390 111894 48442
rect 111956 48390 111958 48442
rect 111796 48388 111820 48390
rect 111876 48388 111900 48390
rect 111956 48388 111980 48390
rect 111740 48368 112036 48388
rect 96380 47900 96676 47920
rect 96436 47898 96460 47900
rect 96516 47898 96540 47900
rect 96596 47898 96620 47900
rect 96458 47846 96460 47898
rect 96522 47846 96534 47898
rect 96596 47846 96598 47898
rect 96436 47844 96460 47846
rect 96516 47844 96540 47846
rect 96596 47844 96620 47846
rect 96380 47824 96676 47844
rect 81020 47356 81316 47376
rect 81076 47354 81100 47356
rect 81156 47354 81180 47356
rect 81236 47354 81260 47356
rect 81098 47302 81100 47354
rect 81162 47302 81174 47354
rect 81236 47302 81238 47354
rect 81076 47300 81100 47302
rect 81156 47300 81180 47302
rect 81236 47300 81260 47302
rect 81020 47280 81316 47300
rect 111740 47356 112036 47376
rect 111796 47354 111820 47356
rect 111876 47354 111900 47356
rect 111956 47354 111980 47356
rect 111818 47302 111820 47354
rect 111882 47302 111894 47354
rect 111956 47302 111958 47354
rect 111796 47300 111820 47302
rect 111876 47300 111900 47302
rect 111956 47300 111980 47302
rect 111740 47280 112036 47300
rect 96380 46812 96676 46832
rect 96436 46810 96460 46812
rect 96516 46810 96540 46812
rect 96596 46810 96620 46812
rect 96458 46758 96460 46810
rect 96522 46758 96534 46810
rect 96596 46758 96598 46810
rect 96436 46756 96460 46758
rect 96516 46756 96540 46758
rect 96596 46756 96620 46758
rect 96380 46736 96676 46756
rect 81020 46268 81316 46288
rect 81076 46266 81100 46268
rect 81156 46266 81180 46268
rect 81236 46266 81260 46268
rect 81098 46214 81100 46266
rect 81162 46214 81174 46266
rect 81236 46214 81238 46266
rect 81076 46212 81100 46214
rect 81156 46212 81180 46214
rect 81236 46212 81260 46214
rect 81020 46192 81316 46212
rect 111740 46268 112036 46288
rect 111796 46266 111820 46268
rect 111876 46266 111900 46268
rect 111956 46266 111980 46268
rect 111818 46214 111820 46266
rect 111882 46214 111894 46266
rect 111956 46214 111958 46266
rect 111796 46212 111820 46214
rect 111876 46212 111900 46214
rect 111956 46212 111980 46214
rect 111740 46192 112036 46212
rect 96380 45724 96676 45744
rect 96436 45722 96460 45724
rect 96516 45722 96540 45724
rect 96596 45722 96620 45724
rect 96458 45670 96460 45722
rect 96522 45670 96534 45722
rect 96596 45670 96598 45722
rect 96436 45668 96460 45670
rect 96516 45668 96540 45670
rect 96596 45668 96620 45670
rect 96380 45648 96676 45668
rect 81020 45180 81316 45200
rect 81076 45178 81100 45180
rect 81156 45178 81180 45180
rect 81236 45178 81260 45180
rect 81098 45126 81100 45178
rect 81162 45126 81174 45178
rect 81236 45126 81238 45178
rect 81076 45124 81100 45126
rect 81156 45124 81180 45126
rect 81236 45124 81260 45126
rect 81020 45104 81316 45124
rect 111740 45180 112036 45200
rect 111796 45178 111820 45180
rect 111876 45178 111900 45180
rect 111956 45178 111980 45180
rect 111818 45126 111820 45178
rect 111882 45126 111894 45178
rect 111956 45126 111958 45178
rect 111796 45124 111820 45126
rect 111876 45124 111900 45126
rect 111956 45124 111980 45126
rect 111740 45104 112036 45124
rect 96380 44636 96676 44656
rect 96436 44634 96460 44636
rect 96516 44634 96540 44636
rect 96596 44634 96620 44636
rect 96458 44582 96460 44634
rect 96522 44582 96534 44634
rect 96596 44582 96598 44634
rect 96436 44580 96460 44582
rect 96516 44580 96540 44582
rect 96596 44580 96620 44582
rect 96380 44560 96676 44580
rect 81020 44092 81316 44112
rect 81076 44090 81100 44092
rect 81156 44090 81180 44092
rect 81236 44090 81260 44092
rect 81098 44038 81100 44090
rect 81162 44038 81174 44090
rect 81236 44038 81238 44090
rect 81076 44036 81100 44038
rect 81156 44036 81180 44038
rect 81236 44036 81260 44038
rect 81020 44016 81316 44036
rect 111740 44092 112036 44112
rect 111796 44090 111820 44092
rect 111876 44090 111900 44092
rect 111956 44090 111980 44092
rect 111818 44038 111820 44090
rect 111882 44038 111894 44090
rect 111956 44038 111958 44090
rect 111796 44036 111820 44038
rect 111876 44036 111900 44038
rect 111956 44036 111980 44038
rect 111740 44016 112036 44036
rect 96380 43548 96676 43568
rect 96436 43546 96460 43548
rect 96516 43546 96540 43548
rect 96596 43546 96620 43548
rect 96458 43494 96460 43546
rect 96522 43494 96534 43546
rect 96596 43494 96598 43546
rect 96436 43492 96460 43494
rect 96516 43492 96540 43494
rect 96596 43492 96620 43494
rect 96380 43472 96676 43492
rect 81020 43004 81316 43024
rect 81076 43002 81100 43004
rect 81156 43002 81180 43004
rect 81236 43002 81260 43004
rect 81098 42950 81100 43002
rect 81162 42950 81174 43002
rect 81236 42950 81238 43002
rect 81076 42948 81100 42950
rect 81156 42948 81180 42950
rect 81236 42948 81260 42950
rect 81020 42928 81316 42948
rect 111740 43004 112036 43024
rect 111796 43002 111820 43004
rect 111876 43002 111900 43004
rect 111956 43002 111980 43004
rect 111818 42950 111820 43002
rect 111882 42950 111894 43002
rect 111956 42950 111958 43002
rect 111796 42948 111820 42950
rect 111876 42948 111900 42950
rect 111956 42948 111980 42950
rect 111740 42928 112036 42948
rect 96380 42460 96676 42480
rect 96436 42458 96460 42460
rect 96516 42458 96540 42460
rect 96596 42458 96620 42460
rect 96458 42406 96460 42458
rect 96522 42406 96534 42458
rect 96596 42406 96598 42458
rect 96436 42404 96460 42406
rect 96516 42404 96540 42406
rect 96596 42404 96620 42406
rect 96380 42384 96676 42404
rect 81020 41916 81316 41936
rect 81076 41914 81100 41916
rect 81156 41914 81180 41916
rect 81236 41914 81260 41916
rect 81098 41862 81100 41914
rect 81162 41862 81174 41914
rect 81236 41862 81238 41914
rect 81076 41860 81100 41862
rect 81156 41860 81180 41862
rect 81236 41860 81260 41862
rect 81020 41840 81316 41860
rect 111740 41916 112036 41936
rect 111796 41914 111820 41916
rect 111876 41914 111900 41916
rect 111956 41914 111980 41916
rect 111818 41862 111820 41914
rect 111882 41862 111894 41914
rect 111956 41862 111958 41914
rect 111796 41860 111820 41862
rect 111876 41860 111900 41862
rect 111956 41860 111980 41862
rect 111740 41840 112036 41860
rect 96380 41372 96676 41392
rect 96436 41370 96460 41372
rect 96516 41370 96540 41372
rect 96596 41370 96620 41372
rect 96458 41318 96460 41370
rect 96522 41318 96534 41370
rect 96596 41318 96598 41370
rect 96436 41316 96460 41318
rect 96516 41316 96540 41318
rect 96596 41316 96620 41318
rect 96380 41296 96676 41316
rect 81020 40828 81316 40848
rect 81076 40826 81100 40828
rect 81156 40826 81180 40828
rect 81236 40826 81260 40828
rect 81098 40774 81100 40826
rect 81162 40774 81174 40826
rect 81236 40774 81238 40826
rect 81076 40772 81100 40774
rect 81156 40772 81180 40774
rect 81236 40772 81260 40774
rect 81020 40752 81316 40772
rect 111740 40828 112036 40848
rect 111796 40826 111820 40828
rect 111876 40826 111900 40828
rect 111956 40826 111980 40828
rect 111818 40774 111820 40826
rect 111882 40774 111894 40826
rect 111956 40774 111958 40826
rect 111796 40772 111820 40774
rect 111876 40772 111900 40774
rect 111956 40772 111980 40774
rect 111740 40752 112036 40772
rect 96380 40284 96676 40304
rect 96436 40282 96460 40284
rect 96516 40282 96540 40284
rect 96596 40282 96620 40284
rect 96458 40230 96460 40282
rect 96522 40230 96534 40282
rect 96596 40230 96598 40282
rect 96436 40228 96460 40230
rect 96516 40228 96540 40230
rect 96596 40228 96620 40230
rect 96380 40208 96676 40228
rect 81020 39740 81316 39760
rect 81076 39738 81100 39740
rect 81156 39738 81180 39740
rect 81236 39738 81260 39740
rect 81098 39686 81100 39738
rect 81162 39686 81174 39738
rect 81236 39686 81238 39738
rect 81076 39684 81100 39686
rect 81156 39684 81180 39686
rect 81236 39684 81260 39686
rect 81020 39664 81316 39684
rect 111740 39740 112036 39760
rect 111796 39738 111820 39740
rect 111876 39738 111900 39740
rect 111956 39738 111980 39740
rect 111818 39686 111820 39738
rect 111882 39686 111894 39738
rect 111956 39686 111958 39738
rect 111796 39684 111820 39686
rect 111876 39684 111900 39686
rect 111956 39684 111980 39686
rect 111740 39664 112036 39684
rect 96380 39196 96676 39216
rect 96436 39194 96460 39196
rect 96516 39194 96540 39196
rect 96596 39194 96620 39196
rect 96458 39142 96460 39194
rect 96522 39142 96534 39194
rect 96596 39142 96598 39194
rect 96436 39140 96460 39142
rect 96516 39140 96540 39142
rect 96596 39140 96620 39142
rect 96380 39120 96676 39140
rect 81020 38652 81316 38672
rect 81076 38650 81100 38652
rect 81156 38650 81180 38652
rect 81236 38650 81260 38652
rect 81098 38598 81100 38650
rect 81162 38598 81174 38650
rect 81236 38598 81238 38650
rect 81076 38596 81100 38598
rect 81156 38596 81180 38598
rect 81236 38596 81260 38598
rect 81020 38576 81316 38596
rect 111740 38652 112036 38672
rect 111796 38650 111820 38652
rect 111876 38650 111900 38652
rect 111956 38650 111980 38652
rect 111818 38598 111820 38650
rect 111882 38598 111894 38650
rect 111956 38598 111958 38650
rect 111796 38596 111820 38598
rect 111876 38596 111900 38598
rect 111956 38596 111980 38598
rect 111740 38576 112036 38596
rect 96380 38108 96676 38128
rect 96436 38106 96460 38108
rect 96516 38106 96540 38108
rect 96596 38106 96620 38108
rect 96458 38054 96460 38106
rect 96522 38054 96534 38106
rect 96596 38054 96598 38106
rect 96436 38052 96460 38054
rect 96516 38052 96540 38054
rect 96596 38052 96620 38054
rect 96380 38032 96676 38052
rect 81020 37564 81316 37584
rect 81076 37562 81100 37564
rect 81156 37562 81180 37564
rect 81236 37562 81260 37564
rect 81098 37510 81100 37562
rect 81162 37510 81174 37562
rect 81236 37510 81238 37562
rect 81076 37508 81100 37510
rect 81156 37508 81180 37510
rect 81236 37508 81260 37510
rect 81020 37488 81316 37508
rect 111740 37564 112036 37584
rect 111796 37562 111820 37564
rect 111876 37562 111900 37564
rect 111956 37562 111980 37564
rect 111818 37510 111820 37562
rect 111882 37510 111894 37562
rect 111956 37510 111958 37562
rect 111796 37508 111820 37510
rect 111876 37508 111900 37510
rect 111956 37508 111980 37510
rect 111740 37488 112036 37508
rect 96380 37020 96676 37040
rect 96436 37018 96460 37020
rect 96516 37018 96540 37020
rect 96596 37018 96620 37020
rect 96458 36966 96460 37018
rect 96522 36966 96534 37018
rect 96596 36966 96598 37018
rect 96436 36964 96460 36966
rect 96516 36964 96540 36966
rect 96596 36964 96620 36966
rect 96380 36944 96676 36964
rect 81020 36476 81316 36496
rect 81076 36474 81100 36476
rect 81156 36474 81180 36476
rect 81236 36474 81260 36476
rect 81098 36422 81100 36474
rect 81162 36422 81174 36474
rect 81236 36422 81238 36474
rect 81076 36420 81100 36422
rect 81156 36420 81180 36422
rect 81236 36420 81260 36422
rect 81020 36400 81316 36420
rect 111740 36476 112036 36496
rect 111796 36474 111820 36476
rect 111876 36474 111900 36476
rect 111956 36474 111980 36476
rect 111818 36422 111820 36474
rect 111882 36422 111894 36474
rect 111956 36422 111958 36474
rect 111796 36420 111820 36422
rect 111876 36420 111900 36422
rect 111956 36420 111980 36422
rect 111740 36400 112036 36420
rect 96380 35932 96676 35952
rect 96436 35930 96460 35932
rect 96516 35930 96540 35932
rect 96596 35930 96620 35932
rect 96458 35878 96460 35930
rect 96522 35878 96534 35930
rect 96596 35878 96598 35930
rect 96436 35876 96460 35878
rect 96516 35876 96540 35878
rect 96596 35876 96620 35878
rect 96380 35856 96676 35876
rect 81020 35388 81316 35408
rect 81076 35386 81100 35388
rect 81156 35386 81180 35388
rect 81236 35386 81260 35388
rect 81098 35334 81100 35386
rect 81162 35334 81174 35386
rect 81236 35334 81238 35386
rect 81076 35332 81100 35334
rect 81156 35332 81180 35334
rect 81236 35332 81260 35334
rect 81020 35312 81316 35332
rect 111740 35388 112036 35408
rect 111796 35386 111820 35388
rect 111876 35386 111900 35388
rect 111956 35386 111980 35388
rect 111818 35334 111820 35386
rect 111882 35334 111894 35386
rect 111956 35334 111958 35386
rect 111796 35332 111820 35334
rect 111876 35332 111900 35334
rect 111956 35332 111980 35334
rect 111740 35312 112036 35332
rect 96380 34844 96676 34864
rect 96436 34842 96460 34844
rect 96516 34842 96540 34844
rect 96596 34842 96620 34844
rect 96458 34790 96460 34842
rect 96522 34790 96534 34842
rect 96596 34790 96598 34842
rect 96436 34788 96460 34790
rect 96516 34788 96540 34790
rect 96596 34788 96620 34790
rect 96380 34768 96676 34788
rect 81020 34300 81316 34320
rect 81076 34298 81100 34300
rect 81156 34298 81180 34300
rect 81236 34298 81260 34300
rect 81098 34246 81100 34298
rect 81162 34246 81174 34298
rect 81236 34246 81238 34298
rect 81076 34244 81100 34246
rect 81156 34244 81180 34246
rect 81236 34244 81260 34246
rect 81020 34224 81316 34244
rect 111740 34300 112036 34320
rect 111796 34298 111820 34300
rect 111876 34298 111900 34300
rect 111956 34298 111980 34300
rect 111818 34246 111820 34298
rect 111882 34246 111894 34298
rect 111956 34246 111958 34298
rect 111796 34244 111820 34246
rect 111876 34244 111900 34246
rect 111956 34244 111980 34246
rect 111740 34224 112036 34244
rect 96380 33756 96676 33776
rect 96436 33754 96460 33756
rect 96516 33754 96540 33756
rect 96596 33754 96620 33756
rect 96458 33702 96460 33754
rect 96522 33702 96534 33754
rect 96596 33702 96598 33754
rect 96436 33700 96460 33702
rect 96516 33700 96540 33702
rect 96596 33700 96620 33702
rect 96380 33680 96676 33700
rect 81020 33212 81316 33232
rect 81076 33210 81100 33212
rect 81156 33210 81180 33212
rect 81236 33210 81260 33212
rect 81098 33158 81100 33210
rect 81162 33158 81174 33210
rect 81236 33158 81238 33210
rect 81076 33156 81100 33158
rect 81156 33156 81180 33158
rect 81236 33156 81260 33158
rect 81020 33136 81316 33156
rect 111740 33212 112036 33232
rect 111796 33210 111820 33212
rect 111876 33210 111900 33212
rect 111956 33210 111980 33212
rect 111818 33158 111820 33210
rect 111882 33158 111894 33210
rect 111956 33158 111958 33210
rect 111796 33156 111820 33158
rect 111876 33156 111900 33158
rect 111956 33156 111980 33158
rect 111740 33136 112036 33156
rect 96380 32668 96676 32688
rect 96436 32666 96460 32668
rect 96516 32666 96540 32668
rect 96596 32666 96620 32668
rect 96458 32614 96460 32666
rect 96522 32614 96534 32666
rect 96596 32614 96598 32666
rect 96436 32612 96460 32614
rect 96516 32612 96540 32614
rect 96596 32612 96620 32614
rect 96380 32592 96676 32612
rect 81020 32124 81316 32144
rect 81076 32122 81100 32124
rect 81156 32122 81180 32124
rect 81236 32122 81260 32124
rect 81098 32070 81100 32122
rect 81162 32070 81174 32122
rect 81236 32070 81238 32122
rect 81076 32068 81100 32070
rect 81156 32068 81180 32070
rect 81236 32068 81260 32070
rect 81020 32048 81316 32068
rect 111740 32124 112036 32144
rect 111796 32122 111820 32124
rect 111876 32122 111900 32124
rect 111956 32122 111980 32124
rect 111818 32070 111820 32122
rect 111882 32070 111894 32122
rect 111956 32070 111958 32122
rect 111796 32068 111820 32070
rect 111876 32068 111900 32070
rect 111956 32068 111980 32070
rect 111740 32048 112036 32068
rect 96380 31580 96676 31600
rect 96436 31578 96460 31580
rect 96516 31578 96540 31580
rect 96596 31578 96620 31580
rect 96458 31526 96460 31578
rect 96522 31526 96534 31578
rect 96596 31526 96598 31578
rect 96436 31524 96460 31526
rect 96516 31524 96540 31526
rect 96596 31524 96620 31526
rect 96380 31504 96676 31524
rect 81020 31036 81316 31056
rect 81076 31034 81100 31036
rect 81156 31034 81180 31036
rect 81236 31034 81260 31036
rect 81098 30982 81100 31034
rect 81162 30982 81174 31034
rect 81236 30982 81238 31034
rect 81076 30980 81100 30982
rect 81156 30980 81180 30982
rect 81236 30980 81260 30982
rect 81020 30960 81316 30980
rect 111740 31036 112036 31056
rect 111796 31034 111820 31036
rect 111876 31034 111900 31036
rect 111956 31034 111980 31036
rect 111818 30982 111820 31034
rect 111882 30982 111894 31034
rect 111956 30982 111958 31034
rect 111796 30980 111820 30982
rect 111876 30980 111900 30982
rect 111956 30980 111980 30982
rect 111740 30960 112036 30980
rect 96380 30492 96676 30512
rect 96436 30490 96460 30492
rect 96516 30490 96540 30492
rect 96596 30490 96620 30492
rect 96458 30438 96460 30490
rect 96522 30438 96534 30490
rect 96596 30438 96598 30490
rect 96436 30436 96460 30438
rect 96516 30436 96540 30438
rect 96596 30436 96620 30438
rect 96380 30416 96676 30436
rect 81020 29948 81316 29968
rect 81076 29946 81100 29948
rect 81156 29946 81180 29948
rect 81236 29946 81260 29948
rect 81098 29894 81100 29946
rect 81162 29894 81174 29946
rect 81236 29894 81238 29946
rect 81076 29892 81100 29894
rect 81156 29892 81180 29894
rect 81236 29892 81260 29894
rect 81020 29872 81316 29892
rect 111740 29948 112036 29968
rect 111796 29946 111820 29948
rect 111876 29946 111900 29948
rect 111956 29946 111980 29948
rect 111818 29894 111820 29946
rect 111882 29894 111894 29946
rect 111956 29894 111958 29946
rect 111796 29892 111820 29894
rect 111876 29892 111900 29894
rect 111956 29892 111980 29894
rect 111740 29872 112036 29892
rect 96380 29404 96676 29424
rect 96436 29402 96460 29404
rect 96516 29402 96540 29404
rect 96596 29402 96620 29404
rect 96458 29350 96460 29402
rect 96522 29350 96534 29402
rect 96596 29350 96598 29402
rect 96436 29348 96460 29350
rect 96516 29348 96540 29350
rect 96596 29348 96620 29350
rect 96380 29328 96676 29348
rect 81020 28860 81316 28880
rect 81076 28858 81100 28860
rect 81156 28858 81180 28860
rect 81236 28858 81260 28860
rect 81098 28806 81100 28858
rect 81162 28806 81174 28858
rect 81236 28806 81238 28858
rect 81076 28804 81100 28806
rect 81156 28804 81180 28806
rect 81236 28804 81260 28806
rect 81020 28784 81316 28804
rect 111740 28860 112036 28880
rect 111796 28858 111820 28860
rect 111876 28858 111900 28860
rect 111956 28858 111980 28860
rect 111818 28806 111820 28858
rect 111882 28806 111894 28858
rect 111956 28806 111958 28858
rect 111796 28804 111820 28806
rect 111876 28804 111900 28806
rect 111956 28804 111980 28806
rect 111740 28784 112036 28804
rect 96380 28316 96676 28336
rect 96436 28314 96460 28316
rect 96516 28314 96540 28316
rect 96596 28314 96620 28316
rect 96458 28262 96460 28314
rect 96522 28262 96534 28314
rect 96596 28262 96598 28314
rect 96436 28260 96460 28262
rect 96516 28260 96540 28262
rect 96596 28260 96620 28262
rect 96380 28240 96676 28260
rect 81020 27772 81316 27792
rect 81076 27770 81100 27772
rect 81156 27770 81180 27772
rect 81236 27770 81260 27772
rect 81098 27718 81100 27770
rect 81162 27718 81174 27770
rect 81236 27718 81238 27770
rect 81076 27716 81100 27718
rect 81156 27716 81180 27718
rect 81236 27716 81260 27718
rect 81020 27696 81316 27716
rect 111740 27772 112036 27792
rect 111796 27770 111820 27772
rect 111876 27770 111900 27772
rect 111956 27770 111980 27772
rect 111818 27718 111820 27770
rect 111882 27718 111894 27770
rect 111956 27718 111958 27770
rect 111796 27716 111820 27718
rect 111876 27716 111900 27718
rect 111956 27716 111980 27718
rect 111740 27696 112036 27716
rect 96380 27228 96676 27248
rect 96436 27226 96460 27228
rect 96516 27226 96540 27228
rect 96596 27226 96620 27228
rect 96458 27174 96460 27226
rect 96522 27174 96534 27226
rect 96596 27174 96598 27226
rect 96436 27172 96460 27174
rect 96516 27172 96540 27174
rect 96596 27172 96620 27174
rect 96380 27152 96676 27172
rect 81020 26684 81316 26704
rect 81076 26682 81100 26684
rect 81156 26682 81180 26684
rect 81236 26682 81260 26684
rect 81098 26630 81100 26682
rect 81162 26630 81174 26682
rect 81236 26630 81238 26682
rect 81076 26628 81100 26630
rect 81156 26628 81180 26630
rect 81236 26628 81260 26630
rect 81020 26608 81316 26628
rect 111740 26684 112036 26704
rect 111796 26682 111820 26684
rect 111876 26682 111900 26684
rect 111956 26682 111980 26684
rect 111818 26630 111820 26682
rect 111882 26630 111894 26682
rect 111956 26630 111958 26682
rect 111796 26628 111820 26630
rect 111876 26628 111900 26630
rect 111956 26628 111980 26630
rect 111740 26608 112036 26628
rect 96380 26140 96676 26160
rect 96436 26138 96460 26140
rect 96516 26138 96540 26140
rect 96596 26138 96620 26140
rect 96458 26086 96460 26138
rect 96522 26086 96534 26138
rect 96596 26086 96598 26138
rect 96436 26084 96460 26086
rect 96516 26084 96540 26086
rect 96596 26084 96620 26086
rect 96380 26064 96676 26084
rect 81020 25596 81316 25616
rect 81076 25594 81100 25596
rect 81156 25594 81180 25596
rect 81236 25594 81260 25596
rect 81098 25542 81100 25594
rect 81162 25542 81174 25594
rect 81236 25542 81238 25594
rect 81076 25540 81100 25542
rect 81156 25540 81180 25542
rect 81236 25540 81260 25542
rect 81020 25520 81316 25540
rect 111740 25596 112036 25616
rect 111796 25594 111820 25596
rect 111876 25594 111900 25596
rect 111956 25594 111980 25596
rect 111818 25542 111820 25594
rect 111882 25542 111894 25594
rect 111956 25542 111958 25594
rect 111796 25540 111820 25542
rect 111876 25540 111900 25542
rect 111956 25540 111980 25542
rect 111740 25520 112036 25540
rect 96380 25052 96676 25072
rect 96436 25050 96460 25052
rect 96516 25050 96540 25052
rect 96596 25050 96620 25052
rect 96458 24998 96460 25050
rect 96522 24998 96534 25050
rect 96596 24998 96598 25050
rect 96436 24996 96460 24998
rect 96516 24996 96540 24998
rect 96596 24996 96620 24998
rect 96380 24976 96676 24996
rect 81020 24508 81316 24528
rect 81076 24506 81100 24508
rect 81156 24506 81180 24508
rect 81236 24506 81260 24508
rect 81098 24454 81100 24506
rect 81162 24454 81174 24506
rect 81236 24454 81238 24506
rect 81076 24452 81100 24454
rect 81156 24452 81180 24454
rect 81236 24452 81260 24454
rect 81020 24432 81316 24452
rect 111740 24508 112036 24528
rect 111796 24506 111820 24508
rect 111876 24506 111900 24508
rect 111956 24506 111980 24508
rect 111818 24454 111820 24506
rect 111882 24454 111894 24506
rect 111956 24454 111958 24506
rect 111796 24452 111820 24454
rect 111876 24452 111900 24454
rect 111956 24452 111980 24454
rect 111740 24432 112036 24452
rect 96380 23964 96676 23984
rect 96436 23962 96460 23964
rect 96516 23962 96540 23964
rect 96596 23962 96620 23964
rect 96458 23910 96460 23962
rect 96522 23910 96534 23962
rect 96596 23910 96598 23962
rect 96436 23908 96460 23910
rect 96516 23908 96540 23910
rect 96596 23908 96620 23910
rect 96380 23888 96676 23908
rect 81020 23420 81316 23440
rect 81076 23418 81100 23420
rect 81156 23418 81180 23420
rect 81236 23418 81260 23420
rect 81098 23366 81100 23418
rect 81162 23366 81174 23418
rect 81236 23366 81238 23418
rect 81076 23364 81100 23366
rect 81156 23364 81180 23366
rect 81236 23364 81260 23366
rect 81020 23344 81316 23364
rect 111740 23420 112036 23440
rect 111796 23418 111820 23420
rect 111876 23418 111900 23420
rect 111956 23418 111980 23420
rect 111818 23366 111820 23418
rect 111882 23366 111894 23418
rect 111956 23366 111958 23418
rect 111796 23364 111820 23366
rect 111876 23364 111900 23366
rect 111956 23364 111980 23366
rect 111740 23344 112036 23364
rect 96380 22876 96676 22896
rect 96436 22874 96460 22876
rect 96516 22874 96540 22876
rect 96596 22874 96620 22876
rect 96458 22822 96460 22874
rect 96522 22822 96534 22874
rect 96596 22822 96598 22874
rect 96436 22820 96460 22822
rect 96516 22820 96540 22822
rect 96596 22820 96620 22822
rect 96380 22800 96676 22820
rect 81020 22332 81316 22352
rect 81076 22330 81100 22332
rect 81156 22330 81180 22332
rect 81236 22330 81260 22332
rect 81098 22278 81100 22330
rect 81162 22278 81174 22330
rect 81236 22278 81238 22330
rect 81076 22276 81100 22278
rect 81156 22276 81180 22278
rect 81236 22276 81260 22278
rect 81020 22256 81316 22276
rect 111740 22332 112036 22352
rect 111796 22330 111820 22332
rect 111876 22330 111900 22332
rect 111956 22330 111980 22332
rect 111818 22278 111820 22330
rect 111882 22278 111894 22330
rect 111956 22278 111958 22330
rect 111796 22276 111820 22278
rect 111876 22276 111900 22278
rect 111956 22276 111980 22278
rect 111740 22256 112036 22276
rect 72988 22066 73108 22094
rect 72884 19304 72936 19310
rect 72884 19246 72936 19252
rect 72896 19174 72924 19246
rect 72884 19168 72936 19174
rect 72884 19110 72936 19116
rect 72988 18834 73016 22066
rect 96380 21788 96676 21808
rect 96436 21786 96460 21788
rect 96516 21786 96540 21788
rect 96596 21786 96620 21788
rect 96458 21734 96460 21786
rect 96522 21734 96534 21786
rect 96596 21734 96598 21786
rect 96436 21732 96460 21734
rect 96516 21732 96540 21734
rect 96596 21732 96620 21734
rect 96380 21712 96676 21732
rect 81020 21244 81316 21264
rect 81076 21242 81100 21244
rect 81156 21242 81180 21244
rect 81236 21242 81260 21244
rect 81098 21190 81100 21242
rect 81162 21190 81174 21242
rect 81236 21190 81238 21242
rect 81076 21188 81100 21190
rect 81156 21188 81180 21190
rect 81236 21188 81260 21190
rect 81020 21168 81316 21188
rect 111740 21244 112036 21264
rect 111796 21242 111820 21244
rect 111876 21242 111900 21244
rect 111956 21242 111980 21244
rect 111818 21190 111820 21242
rect 111882 21190 111894 21242
rect 111956 21190 111958 21242
rect 111796 21188 111820 21190
rect 111876 21188 111900 21190
rect 111956 21188 111980 21190
rect 111740 21168 112036 21188
rect 96380 20700 96676 20720
rect 96436 20698 96460 20700
rect 96516 20698 96540 20700
rect 96596 20698 96620 20700
rect 96458 20646 96460 20698
rect 96522 20646 96534 20698
rect 96596 20646 96598 20698
rect 96436 20644 96460 20646
rect 96516 20644 96540 20646
rect 96596 20644 96620 20646
rect 96380 20624 96676 20644
rect 74540 20256 74592 20262
rect 74540 20198 74592 20204
rect 75828 20256 75880 20262
rect 75828 20198 75880 20204
rect 73252 19984 73304 19990
rect 73252 19926 73304 19932
rect 73264 19310 73292 19926
rect 73252 19304 73304 19310
rect 74552 19258 74580 20198
rect 73252 19246 73304 19252
rect 74368 19230 74580 19258
rect 75276 19236 75328 19242
rect 73160 19168 73212 19174
rect 73080 19116 73160 19122
rect 73080 19110 73212 19116
rect 73528 19168 73580 19174
rect 73528 19110 73580 19116
rect 73080 19094 73200 19110
rect 72240 18828 72292 18834
rect 72240 18770 72292 18776
rect 72424 18828 72476 18834
rect 72424 18770 72476 18776
rect 72976 18828 73028 18834
rect 72976 18770 73028 18776
rect 72148 18216 72200 18222
rect 72148 18158 72200 18164
rect 70768 17128 70820 17134
rect 70768 17070 70820 17076
rect 71136 17128 71188 17134
rect 71136 17070 71188 17076
rect 71320 17128 71372 17134
rect 71320 17070 71372 17076
rect 71688 17128 71740 17134
rect 71688 17070 71740 17076
rect 70780 16590 70808 17070
rect 70400 16584 70452 16590
rect 70400 16526 70452 16532
rect 70768 16584 70820 16590
rect 70768 16526 70820 16532
rect 70216 16040 70268 16046
rect 70216 15982 70268 15988
rect 70228 15570 70256 15982
rect 70216 15564 70268 15570
rect 70216 15506 70268 15512
rect 70032 15360 70084 15366
rect 70032 15302 70084 15308
rect 70124 15360 70176 15366
rect 70124 15302 70176 15308
rect 69900 13824 69980 13852
rect 69848 13806 69900 13812
rect 69756 13252 69808 13258
rect 69756 13194 69808 13200
rect 69664 12232 69716 12238
rect 69664 12174 69716 12180
rect 69676 9518 69704 12174
rect 69860 12102 69888 13806
rect 70044 12714 70072 15302
rect 70136 14618 70164 15302
rect 70412 14822 70440 16526
rect 71148 16114 71176 17070
rect 71136 16108 71188 16114
rect 71136 16050 71188 16056
rect 70492 16040 70544 16046
rect 70492 15982 70544 15988
rect 70504 15706 70532 15982
rect 71332 15978 71360 17070
rect 71504 16992 71556 16998
rect 71504 16934 71556 16940
rect 71516 16658 71544 16934
rect 71504 16652 71556 16658
rect 71504 16594 71556 16600
rect 71700 16590 71728 17070
rect 71688 16584 71740 16590
rect 71688 16526 71740 16532
rect 71700 16046 71728 16526
rect 71872 16244 71924 16250
rect 71872 16186 71924 16192
rect 71688 16040 71740 16046
rect 71688 15982 71740 15988
rect 71320 15972 71372 15978
rect 71320 15914 71372 15920
rect 70492 15700 70544 15706
rect 70492 15642 70544 15648
rect 71700 15570 71728 15982
rect 71884 15638 71912 16186
rect 72056 16040 72108 16046
rect 72056 15982 72108 15988
rect 72068 15706 72096 15982
rect 72056 15700 72108 15706
rect 72056 15642 72108 15648
rect 71872 15632 71924 15638
rect 71872 15574 71924 15580
rect 71688 15564 71740 15570
rect 71688 15506 71740 15512
rect 72160 15502 72188 18158
rect 72148 15496 72200 15502
rect 72148 15438 72200 15444
rect 70400 14816 70452 14822
rect 70400 14758 70452 14764
rect 70124 14612 70176 14618
rect 70124 14554 70176 14560
rect 70308 14408 70360 14414
rect 70308 14350 70360 14356
rect 70216 14000 70268 14006
rect 70216 13942 70268 13948
rect 70228 13326 70256 13942
rect 70320 13938 70348 14350
rect 70308 13932 70360 13938
rect 70308 13874 70360 13880
rect 70320 13394 70348 13874
rect 72252 13462 72280 18770
rect 72332 17332 72384 17338
rect 72332 17274 72384 17280
rect 72344 15910 72372 17274
rect 72516 16992 72568 16998
rect 72516 16934 72568 16940
rect 72424 16652 72476 16658
rect 72424 16594 72476 16600
rect 72332 15904 72384 15910
rect 72332 15846 72384 15852
rect 72436 13530 72464 16594
rect 72528 13870 72556 16934
rect 72884 16652 72936 16658
rect 72884 16594 72936 16600
rect 72896 16250 72924 16594
rect 72884 16244 72936 16250
rect 72884 16186 72936 16192
rect 72516 13864 72568 13870
rect 72516 13806 72568 13812
rect 72424 13524 72476 13530
rect 72424 13466 72476 13472
rect 72240 13456 72292 13462
rect 72240 13398 72292 13404
rect 70308 13388 70360 13394
rect 70308 13330 70360 13336
rect 71136 13388 71188 13394
rect 71136 13330 71188 13336
rect 70216 13320 70268 13326
rect 70216 13262 70268 13268
rect 70124 13184 70176 13190
rect 70124 13126 70176 13132
rect 70136 12782 70164 13126
rect 70228 12850 70256 13262
rect 70676 13184 70728 13190
rect 70676 13126 70728 13132
rect 70216 12844 70268 12850
rect 70216 12786 70268 12792
rect 70124 12776 70176 12782
rect 70124 12718 70176 12724
rect 70032 12708 70084 12714
rect 70032 12650 70084 12656
rect 69848 12096 69900 12102
rect 69848 12038 69900 12044
rect 69664 9512 69716 9518
rect 69664 9454 69716 9460
rect 70032 8560 70084 8566
rect 70032 8502 70084 8508
rect 69756 6656 69808 6662
rect 69756 6598 69808 6604
rect 69848 6656 69900 6662
rect 69848 6598 69900 6604
rect 69768 6322 69796 6598
rect 69572 6316 69624 6322
rect 69572 6258 69624 6264
rect 69756 6316 69808 6322
rect 69756 6258 69808 6264
rect 69664 5772 69716 5778
rect 69664 5714 69716 5720
rect 69386 4720 69442 4729
rect 69386 4655 69442 4664
rect 69400 3602 69428 4655
rect 69480 4072 69532 4078
rect 69480 4014 69532 4020
rect 69112 3596 69164 3602
rect 69112 3538 69164 3544
rect 69388 3596 69440 3602
rect 69388 3538 69440 3544
rect 69020 2576 69072 2582
rect 69020 2518 69072 2524
rect 69112 2304 69164 2310
rect 69112 2246 69164 2252
rect 69124 800 69152 2246
rect 69492 800 69520 4014
rect 69676 3670 69704 5714
rect 69860 3670 69888 6598
rect 69664 3664 69716 3670
rect 69664 3606 69716 3612
rect 69848 3664 69900 3670
rect 69848 3606 69900 3612
rect 69940 3664 69992 3670
rect 69940 3606 69992 3612
rect 69572 3596 69624 3602
rect 69572 3538 69624 3544
rect 69584 1154 69612 3538
rect 69754 3496 69810 3505
rect 69754 3431 69810 3440
rect 69768 3398 69796 3431
rect 69756 3392 69808 3398
rect 69756 3334 69808 3340
rect 69952 3194 69980 3606
rect 70044 3398 70072 8502
rect 70136 7818 70164 12718
rect 70400 11348 70452 11354
rect 70400 11290 70452 11296
rect 70124 7812 70176 7818
rect 70124 7754 70176 7760
rect 70308 7812 70360 7818
rect 70308 7754 70360 7760
rect 70320 6254 70348 7754
rect 70308 6248 70360 6254
rect 70412 6225 70440 11290
rect 70688 6866 70716 13126
rect 70952 12096 71004 12102
rect 70952 12038 71004 12044
rect 70964 6934 70992 12038
rect 71148 11354 71176 13330
rect 72988 12782 73016 18770
rect 73080 17338 73108 19094
rect 73252 18896 73304 18902
rect 73252 18838 73304 18844
rect 73068 17332 73120 17338
rect 73068 17274 73120 17280
rect 73264 17134 73292 18838
rect 73540 18222 73568 19110
rect 74368 18902 74396 19230
rect 75276 19178 75328 19184
rect 75000 19168 75052 19174
rect 75000 19110 75052 19116
rect 74356 18896 74408 18902
rect 74356 18838 74408 18844
rect 74264 18828 74316 18834
rect 74264 18770 74316 18776
rect 74276 18698 74304 18770
rect 74264 18692 74316 18698
rect 74264 18634 74316 18640
rect 73896 18624 73948 18630
rect 73896 18566 73948 18572
rect 73528 18216 73580 18222
rect 73528 18158 73580 18164
rect 73252 17128 73304 17134
rect 73252 17070 73304 17076
rect 73264 16726 73292 17070
rect 73252 16720 73304 16726
rect 73252 16662 73304 16668
rect 73068 16652 73120 16658
rect 73068 16594 73120 16600
rect 73080 13394 73108 16594
rect 73540 14890 73568 18158
rect 73620 18080 73672 18086
rect 73620 18022 73672 18028
rect 73632 16046 73660 18022
rect 73620 16040 73672 16046
rect 73620 15982 73672 15988
rect 73528 14884 73580 14890
rect 73528 14826 73580 14832
rect 73908 14550 73936 18566
rect 74276 17134 74304 18634
rect 74264 17128 74316 17134
rect 74264 17070 74316 17076
rect 73896 14544 73948 14550
rect 73896 14486 73948 14492
rect 74368 14482 74396 18838
rect 75012 18834 75040 19110
rect 75000 18828 75052 18834
rect 75000 18770 75052 18776
rect 75092 18760 75144 18766
rect 75092 18702 75144 18708
rect 75104 17202 75132 18702
rect 75092 17196 75144 17202
rect 75092 17138 75144 17144
rect 75288 16658 75316 19178
rect 75840 18630 75868 20198
rect 81020 20156 81316 20176
rect 81076 20154 81100 20156
rect 81156 20154 81180 20156
rect 81236 20154 81260 20156
rect 81098 20102 81100 20154
rect 81162 20102 81174 20154
rect 81236 20102 81238 20154
rect 81076 20100 81100 20102
rect 81156 20100 81180 20102
rect 81236 20100 81260 20102
rect 81020 20080 81316 20100
rect 111740 20156 112036 20176
rect 111796 20154 111820 20156
rect 111876 20154 111900 20156
rect 111956 20154 111980 20156
rect 111818 20102 111820 20154
rect 111882 20102 111894 20154
rect 111956 20102 111958 20154
rect 111796 20100 111820 20102
rect 111876 20100 111900 20102
rect 111956 20100 111980 20102
rect 111740 20080 112036 20100
rect 121748 20058 121776 117098
rect 124324 116346 124352 117098
rect 127100 116444 127396 116464
rect 127156 116442 127180 116444
rect 127236 116442 127260 116444
rect 127316 116442 127340 116444
rect 127178 116390 127180 116442
rect 127242 116390 127254 116442
rect 127316 116390 127318 116442
rect 127156 116388 127180 116390
rect 127236 116388 127260 116390
rect 127316 116388 127340 116390
rect 127100 116368 127396 116388
rect 128924 116346 128952 117098
rect 124312 116340 124364 116346
rect 124312 116282 124364 116288
rect 128912 116340 128964 116346
rect 128912 116282 128964 116288
rect 127100 115356 127396 115376
rect 127156 115354 127180 115356
rect 127236 115354 127260 115356
rect 127316 115354 127340 115356
rect 127178 115302 127180 115354
rect 127242 115302 127254 115354
rect 127316 115302 127318 115354
rect 127156 115300 127180 115302
rect 127236 115300 127260 115302
rect 127316 115300 127340 115302
rect 127100 115280 127396 115300
rect 127100 114268 127396 114288
rect 127156 114266 127180 114268
rect 127236 114266 127260 114268
rect 127316 114266 127340 114268
rect 127178 114214 127180 114266
rect 127242 114214 127254 114266
rect 127316 114214 127318 114266
rect 127156 114212 127180 114214
rect 127236 114212 127260 114214
rect 127316 114212 127340 114214
rect 127100 114192 127396 114212
rect 127100 113180 127396 113200
rect 127156 113178 127180 113180
rect 127236 113178 127260 113180
rect 127316 113178 127340 113180
rect 127178 113126 127180 113178
rect 127242 113126 127254 113178
rect 127316 113126 127318 113178
rect 127156 113124 127180 113126
rect 127236 113124 127260 113126
rect 127316 113124 127340 113126
rect 127100 113104 127396 113124
rect 127100 112092 127396 112112
rect 127156 112090 127180 112092
rect 127236 112090 127260 112092
rect 127316 112090 127340 112092
rect 127178 112038 127180 112090
rect 127242 112038 127254 112090
rect 127316 112038 127318 112090
rect 127156 112036 127180 112038
rect 127236 112036 127260 112038
rect 127316 112036 127340 112038
rect 127100 112016 127396 112036
rect 127100 111004 127396 111024
rect 127156 111002 127180 111004
rect 127236 111002 127260 111004
rect 127316 111002 127340 111004
rect 127178 110950 127180 111002
rect 127242 110950 127254 111002
rect 127316 110950 127318 111002
rect 127156 110948 127180 110950
rect 127236 110948 127260 110950
rect 127316 110948 127340 110950
rect 127100 110928 127396 110948
rect 127100 109916 127396 109936
rect 127156 109914 127180 109916
rect 127236 109914 127260 109916
rect 127316 109914 127340 109916
rect 127178 109862 127180 109914
rect 127242 109862 127254 109914
rect 127316 109862 127318 109914
rect 127156 109860 127180 109862
rect 127236 109860 127260 109862
rect 127316 109860 127340 109862
rect 127100 109840 127396 109860
rect 127100 108828 127396 108848
rect 127156 108826 127180 108828
rect 127236 108826 127260 108828
rect 127316 108826 127340 108828
rect 127178 108774 127180 108826
rect 127242 108774 127254 108826
rect 127316 108774 127318 108826
rect 127156 108772 127180 108774
rect 127236 108772 127260 108774
rect 127316 108772 127340 108774
rect 127100 108752 127396 108772
rect 127100 107740 127396 107760
rect 127156 107738 127180 107740
rect 127236 107738 127260 107740
rect 127316 107738 127340 107740
rect 127178 107686 127180 107738
rect 127242 107686 127254 107738
rect 127316 107686 127318 107738
rect 127156 107684 127180 107686
rect 127236 107684 127260 107686
rect 127316 107684 127340 107686
rect 127100 107664 127396 107684
rect 127100 106652 127396 106672
rect 127156 106650 127180 106652
rect 127236 106650 127260 106652
rect 127316 106650 127340 106652
rect 127178 106598 127180 106650
rect 127242 106598 127254 106650
rect 127316 106598 127318 106650
rect 127156 106596 127180 106598
rect 127236 106596 127260 106598
rect 127316 106596 127340 106598
rect 127100 106576 127396 106596
rect 127100 105564 127396 105584
rect 127156 105562 127180 105564
rect 127236 105562 127260 105564
rect 127316 105562 127340 105564
rect 127178 105510 127180 105562
rect 127242 105510 127254 105562
rect 127316 105510 127318 105562
rect 127156 105508 127180 105510
rect 127236 105508 127260 105510
rect 127316 105508 127340 105510
rect 127100 105488 127396 105508
rect 127100 104476 127396 104496
rect 127156 104474 127180 104476
rect 127236 104474 127260 104476
rect 127316 104474 127340 104476
rect 127178 104422 127180 104474
rect 127242 104422 127254 104474
rect 127316 104422 127318 104474
rect 127156 104420 127180 104422
rect 127236 104420 127260 104422
rect 127316 104420 127340 104422
rect 127100 104400 127396 104420
rect 127100 103388 127396 103408
rect 127156 103386 127180 103388
rect 127236 103386 127260 103388
rect 127316 103386 127340 103388
rect 127178 103334 127180 103386
rect 127242 103334 127254 103386
rect 127316 103334 127318 103386
rect 127156 103332 127180 103334
rect 127236 103332 127260 103334
rect 127316 103332 127340 103334
rect 127100 103312 127396 103332
rect 127100 102300 127396 102320
rect 127156 102298 127180 102300
rect 127236 102298 127260 102300
rect 127316 102298 127340 102300
rect 127178 102246 127180 102298
rect 127242 102246 127254 102298
rect 127316 102246 127318 102298
rect 127156 102244 127180 102246
rect 127236 102244 127260 102246
rect 127316 102244 127340 102246
rect 127100 102224 127396 102244
rect 127100 101212 127396 101232
rect 127156 101210 127180 101212
rect 127236 101210 127260 101212
rect 127316 101210 127340 101212
rect 127178 101158 127180 101210
rect 127242 101158 127254 101210
rect 127316 101158 127318 101210
rect 127156 101156 127180 101158
rect 127236 101156 127260 101158
rect 127316 101156 127340 101158
rect 127100 101136 127396 101156
rect 127100 100124 127396 100144
rect 127156 100122 127180 100124
rect 127236 100122 127260 100124
rect 127316 100122 127340 100124
rect 127178 100070 127180 100122
rect 127242 100070 127254 100122
rect 127316 100070 127318 100122
rect 127156 100068 127180 100070
rect 127236 100068 127260 100070
rect 127316 100068 127340 100070
rect 127100 100048 127396 100068
rect 127100 99036 127396 99056
rect 127156 99034 127180 99036
rect 127236 99034 127260 99036
rect 127316 99034 127340 99036
rect 127178 98982 127180 99034
rect 127242 98982 127254 99034
rect 127316 98982 127318 99034
rect 127156 98980 127180 98982
rect 127236 98980 127260 98982
rect 127316 98980 127340 98982
rect 127100 98960 127396 98980
rect 127100 97948 127396 97968
rect 127156 97946 127180 97948
rect 127236 97946 127260 97948
rect 127316 97946 127340 97948
rect 127178 97894 127180 97946
rect 127242 97894 127254 97946
rect 127316 97894 127318 97946
rect 127156 97892 127180 97894
rect 127236 97892 127260 97894
rect 127316 97892 127340 97894
rect 127100 97872 127396 97892
rect 127100 96860 127396 96880
rect 127156 96858 127180 96860
rect 127236 96858 127260 96860
rect 127316 96858 127340 96860
rect 127178 96806 127180 96858
rect 127242 96806 127254 96858
rect 127316 96806 127318 96858
rect 127156 96804 127180 96806
rect 127236 96804 127260 96806
rect 127316 96804 127340 96806
rect 127100 96784 127396 96804
rect 127100 95772 127396 95792
rect 127156 95770 127180 95772
rect 127236 95770 127260 95772
rect 127316 95770 127340 95772
rect 127178 95718 127180 95770
rect 127242 95718 127254 95770
rect 127316 95718 127318 95770
rect 127156 95716 127180 95718
rect 127236 95716 127260 95718
rect 127316 95716 127340 95718
rect 127100 95696 127396 95716
rect 127100 94684 127396 94704
rect 127156 94682 127180 94684
rect 127236 94682 127260 94684
rect 127316 94682 127340 94684
rect 127178 94630 127180 94682
rect 127242 94630 127254 94682
rect 127316 94630 127318 94682
rect 127156 94628 127180 94630
rect 127236 94628 127260 94630
rect 127316 94628 127340 94630
rect 127100 94608 127396 94628
rect 127100 93596 127396 93616
rect 127156 93594 127180 93596
rect 127236 93594 127260 93596
rect 127316 93594 127340 93596
rect 127178 93542 127180 93594
rect 127242 93542 127254 93594
rect 127316 93542 127318 93594
rect 127156 93540 127180 93542
rect 127236 93540 127260 93542
rect 127316 93540 127340 93542
rect 127100 93520 127396 93540
rect 127100 92508 127396 92528
rect 127156 92506 127180 92508
rect 127236 92506 127260 92508
rect 127316 92506 127340 92508
rect 127178 92454 127180 92506
rect 127242 92454 127254 92506
rect 127316 92454 127318 92506
rect 127156 92452 127180 92454
rect 127236 92452 127260 92454
rect 127316 92452 127340 92454
rect 127100 92432 127396 92452
rect 127100 91420 127396 91440
rect 127156 91418 127180 91420
rect 127236 91418 127260 91420
rect 127316 91418 127340 91420
rect 127178 91366 127180 91418
rect 127242 91366 127254 91418
rect 127316 91366 127318 91418
rect 127156 91364 127180 91366
rect 127236 91364 127260 91366
rect 127316 91364 127340 91366
rect 127100 91344 127396 91364
rect 127100 90332 127396 90352
rect 127156 90330 127180 90332
rect 127236 90330 127260 90332
rect 127316 90330 127340 90332
rect 127178 90278 127180 90330
rect 127242 90278 127254 90330
rect 127316 90278 127318 90330
rect 127156 90276 127180 90278
rect 127236 90276 127260 90278
rect 127316 90276 127340 90278
rect 127100 90256 127396 90276
rect 127100 89244 127396 89264
rect 127156 89242 127180 89244
rect 127236 89242 127260 89244
rect 127316 89242 127340 89244
rect 127178 89190 127180 89242
rect 127242 89190 127254 89242
rect 127316 89190 127318 89242
rect 127156 89188 127180 89190
rect 127236 89188 127260 89190
rect 127316 89188 127340 89190
rect 127100 89168 127396 89188
rect 127100 88156 127396 88176
rect 127156 88154 127180 88156
rect 127236 88154 127260 88156
rect 127316 88154 127340 88156
rect 127178 88102 127180 88154
rect 127242 88102 127254 88154
rect 127316 88102 127318 88154
rect 127156 88100 127180 88102
rect 127236 88100 127260 88102
rect 127316 88100 127340 88102
rect 127100 88080 127396 88100
rect 127100 87068 127396 87088
rect 127156 87066 127180 87068
rect 127236 87066 127260 87068
rect 127316 87066 127340 87068
rect 127178 87014 127180 87066
rect 127242 87014 127254 87066
rect 127316 87014 127318 87066
rect 127156 87012 127180 87014
rect 127236 87012 127260 87014
rect 127316 87012 127340 87014
rect 127100 86992 127396 87012
rect 127100 85980 127396 86000
rect 127156 85978 127180 85980
rect 127236 85978 127260 85980
rect 127316 85978 127340 85980
rect 127178 85926 127180 85978
rect 127242 85926 127254 85978
rect 127316 85926 127318 85978
rect 127156 85924 127180 85926
rect 127236 85924 127260 85926
rect 127316 85924 127340 85926
rect 127100 85904 127396 85924
rect 127100 84892 127396 84912
rect 127156 84890 127180 84892
rect 127236 84890 127260 84892
rect 127316 84890 127340 84892
rect 127178 84838 127180 84890
rect 127242 84838 127254 84890
rect 127316 84838 127318 84890
rect 127156 84836 127180 84838
rect 127236 84836 127260 84838
rect 127316 84836 127340 84838
rect 127100 84816 127396 84836
rect 127100 83804 127396 83824
rect 127156 83802 127180 83804
rect 127236 83802 127260 83804
rect 127316 83802 127340 83804
rect 127178 83750 127180 83802
rect 127242 83750 127254 83802
rect 127316 83750 127318 83802
rect 127156 83748 127180 83750
rect 127236 83748 127260 83750
rect 127316 83748 127340 83750
rect 127100 83728 127396 83748
rect 127100 82716 127396 82736
rect 127156 82714 127180 82716
rect 127236 82714 127260 82716
rect 127316 82714 127340 82716
rect 127178 82662 127180 82714
rect 127242 82662 127254 82714
rect 127316 82662 127318 82714
rect 127156 82660 127180 82662
rect 127236 82660 127260 82662
rect 127316 82660 127340 82662
rect 127100 82640 127396 82660
rect 127100 81628 127396 81648
rect 127156 81626 127180 81628
rect 127236 81626 127260 81628
rect 127316 81626 127340 81628
rect 127178 81574 127180 81626
rect 127242 81574 127254 81626
rect 127316 81574 127318 81626
rect 127156 81572 127180 81574
rect 127236 81572 127260 81574
rect 127316 81572 127340 81574
rect 127100 81552 127396 81572
rect 127100 80540 127396 80560
rect 127156 80538 127180 80540
rect 127236 80538 127260 80540
rect 127316 80538 127340 80540
rect 127178 80486 127180 80538
rect 127242 80486 127254 80538
rect 127316 80486 127318 80538
rect 127156 80484 127180 80486
rect 127236 80484 127260 80486
rect 127316 80484 127340 80486
rect 127100 80464 127396 80484
rect 127100 79452 127396 79472
rect 127156 79450 127180 79452
rect 127236 79450 127260 79452
rect 127316 79450 127340 79452
rect 127178 79398 127180 79450
rect 127242 79398 127254 79450
rect 127316 79398 127318 79450
rect 127156 79396 127180 79398
rect 127236 79396 127260 79398
rect 127316 79396 127340 79398
rect 127100 79376 127396 79396
rect 127100 78364 127396 78384
rect 127156 78362 127180 78364
rect 127236 78362 127260 78364
rect 127316 78362 127340 78364
rect 127178 78310 127180 78362
rect 127242 78310 127254 78362
rect 127316 78310 127318 78362
rect 127156 78308 127180 78310
rect 127236 78308 127260 78310
rect 127316 78308 127340 78310
rect 127100 78288 127396 78308
rect 127100 77276 127396 77296
rect 127156 77274 127180 77276
rect 127236 77274 127260 77276
rect 127316 77274 127340 77276
rect 127178 77222 127180 77274
rect 127242 77222 127254 77274
rect 127316 77222 127318 77274
rect 127156 77220 127180 77222
rect 127236 77220 127260 77222
rect 127316 77220 127340 77222
rect 127100 77200 127396 77220
rect 127100 76188 127396 76208
rect 127156 76186 127180 76188
rect 127236 76186 127260 76188
rect 127316 76186 127340 76188
rect 127178 76134 127180 76186
rect 127242 76134 127254 76186
rect 127316 76134 127318 76186
rect 127156 76132 127180 76134
rect 127236 76132 127260 76134
rect 127316 76132 127340 76134
rect 127100 76112 127396 76132
rect 127100 75100 127396 75120
rect 127156 75098 127180 75100
rect 127236 75098 127260 75100
rect 127316 75098 127340 75100
rect 127178 75046 127180 75098
rect 127242 75046 127254 75098
rect 127316 75046 127318 75098
rect 127156 75044 127180 75046
rect 127236 75044 127260 75046
rect 127316 75044 127340 75046
rect 127100 75024 127396 75044
rect 127100 74012 127396 74032
rect 127156 74010 127180 74012
rect 127236 74010 127260 74012
rect 127316 74010 127340 74012
rect 127178 73958 127180 74010
rect 127242 73958 127254 74010
rect 127316 73958 127318 74010
rect 127156 73956 127180 73958
rect 127236 73956 127260 73958
rect 127316 73956 127340 73958
rect 127100 73936 127396 73956
rect 127100 72924 127396 72944
rect 127156 72922 127180 72924
rect 127236 72922 127260 72924
rect 127316 72922 127340 72924
rect 127178 72870 127180 72922
rect 127242 72870 127254 72922
rect 127316 72870 127318 72922
rect 127156 72868 127180 72870
rect 127236 72868 127260 72870
rect 127316 72868 127340 72870
rect 127100 72848 127396 72868
rect 127100 71836 127396 71856
rect 127156 71834 127180 71836
rect 127236 71834 127260 71836
rect 127316 71834 127340 71836
rect 127178 71782 127180 71834
rect 127242 71782 127254 71834
rect 127316 71782 127318 71834
rect 127156 71780 127180 71782
rect 127236 71780 127260 71782
rect 127316 71780 127340 71782
rect 127100 71760 127396 71780
rect 127100 70748 127396 70768
rect 127156 70746 127180 70748
rect 127236 70746 127260 70748
rect 127316 70746 127340 70748
rect 127178 70694 127180 70746
rect 127242 70694 127254 70746
rect 127316 70694 127318 70746
rect 127156 70692 127180 70694
rect 127236 70692 127260 70694
rect 127316 70692 127340 70694
rect 127100 70672 127396 70692
rect 127100 69660 127396 69680
rect 127156 69658 127180 69660
rect 127236 69658 127260 69660
rect 127316 69658 127340 69660
rect 127178 69606 127180 69658
rect 127242 69606 127254 69658
rect 127316 69606 127318 69658
rect 127156 69604 127180 69606
rect 127236 69604 127260 69606
rect 127316 69604 127340 69606
rect 127100 69584 127396 69604
rect 127100 68572 127396 68592
rect 127156 68570 127180 68572
rect 127236 68570 127260 68572
rect 127316 68570 127340 68572
rect 127178 68518 127180 68570
rect 127242 68518 127254 68570
rect 127316 68518 127318 68570
rect 127156 68516 127180 68518
rect 127236 68516 127260 68518
rect 127316 68516 127340 68518
rect 127100 68496 127396 68516
rect 127100 67484 127396 67504
rect 127156 67482 127180 67484
rect 127236 67482 127260 67484
rect 127316 67482 127340 67484
rect 127178 67430 127180 67482
rect 127242 67430 127254 67482
rect 127316 67430 127318 67482
rect 127156 67428 127180 67430
rect 127236 67428 127260 67430
rect 127316 67428 127340 67430
rect 127100 67408 127396 67428
rect 127100 66396 127396 66416
rect 127156 66394 127180 66396
rect 127236 66394 127260 66396
rect 127316 66394 127340 66396
rect 127178 66342 127180 66394
rect 127242 66342 127254 66394
rect 127316 66342 127318 66394
rect 127156 66340 127180 66342
rect 127236 66340 127260 66342
rect 127316 66340 127340 66342
rect 127100 66320 127396 66340
rect 127100 65308 127396 65328
rect 127156 65306 127180 65308
rect 127236 65306 127260 65308
rect 127316 65306 127340 65308
rect 127178 65254 127180 65306
rect 127242 65254 127254 65306
rect 127316 65254 127318 65306
rect 127156 65252 127180 65254
rect 127236 65252 127260 65254
rect 127316 65252 127340 65254
rect 127100 65232 127396 65252
rect 127100 64220 127396 64240
rect 127156 64218 127180 64220
rect 127236 64218 127260 64220
rect 127316 64218 127340 64220
rect 127178 64166 127180 64218
rect 127242 64166 127254 64218
rect 127316 64166 127318 64218
rect 127156 64164 127180 64166
rect 127236 64164 127260 64166
rect 127316 64164 127340 64166
rect 127100 64144 127396 64164
rect 127100 63132 127396 63152
rect 127156 63130 127180 63132
rect 127236 63130 127260 63132
rect 127316 63130 127340 63132
rect 127178 63078 127180 63130
rect 127242 63078 127254 63130
rect 127316 63078 127318 63130
rect 127156 63076 127180 63078
rect 127236 63076 127260 63078
rect 127316 63076 127340 63078
rect 127100 63056 127396 63076
rect 127100 62044 127396 62064
rect 127156 62042 127180 62044
rect 127236 62042 127260 62044
rect 127316 62042 127340 62044
rect 127178 61990 127180 62042
rect 127242 61990 127254 62042
rect 127316 61990 127318 62042
rect 127156 61988 127180 61990
rect 127236 61988 127260 61990
rect 127316 61988 127340 61990
rect 127100 61968 127396 61988
rect 127100 60956 127396 60976
rect 127156 60954 127180 60956
rect 127236 60954 127260 60956
rect 127316 60954 127340 60956
rect 127178 60902 127180 60954
rect 127242 60902 127254 60954
rect 127316 60902 127318 60954
rect 127156 60900 127180 60902
rect 127236 60900 127260 60902
rect 127316 60900 127340 60902
rect 127100 60880 127396 60900
rect 127100 59868 127396 59888
rect 127156 59866 127180 59868
rect 127236 59866 127260 59868
rect 127316 59866 127340 59868
rect 127178 59814 127180 59866
rect 127242 59814 127254 59866
rect 127316 59814 127318 59866
rect 127156 59812 127180 59814
rect 127236 59812 127260 59814
rect 127316 59812 127340 59814
rect 127100 59792 127396 59812
rect 127100 58780 127396 58800
rect 127156 58778 127180 58780
rect 127236 58778 127260 58780
rect 127316 58778 127340 58780
rect 127178 58726 127180 58778
rect 127242 58726 127254 58778
rect 127316 58726 127318 58778
rect 127156 58724 127180 58726
rect 127236 58724 127260 58726
rect 127316 58724 127340 58726
rect 127100 58704 127396 58724
rect 127100 57692 127396 57712
rect 127156 57690 127180 57692
rect 127236 57690 127260 57692
rect 127316 57690 127340 57692
rect 127178 57638 127180 57690
rect 127242 57638 127254 57690
rect 127316 57638 127318 57690
rect 127156 57636 127180 57638
rect 127236 57636 127260 57638
rect 127316 57636 127340 57638
rect 127100 57616 127396 57636
rect 127100 56604 127396 56624
rect 127156 56602 127180 56604
rect 127236 56602 127260 56604
rect 127316 56602 127340 56604
rect 127178 56550 127180 56602
rect 127242 56550 127254 56602
rect 127316 56550 127318 56602
rect 127156 56548 127180 56550
rect 127236 56548 127260 56550
rect 127316 56548 127340 56550
rect 127100 56528 127396 56548
rect 127100 55516 127396 55536
rect 127156 55514 127180 55516
rect 127236 55514 127260 55516
rect 127316 55514 127340 55516
rect 127178 55462 127180 55514
rect 127242 55462 127254 55514
rect 127316 55462 127318 55514
rect 127156 55460 127180 55462
rect 127236 55460 127260 55462
rect 127316 55460 127340 55462
rect 127100 55440 127396 55460
rect 127100 54428 127396 54448
rect 127156 54426 127180 54428
rect 127236 54426 127260 54428
rect 127316 54426 127340 54428
rect 127178 54374 127180 54426
rect 127242 54374 127254 54426
rect 127316 54374 127318 54426
rect 127156 54372 127180 54374
rect 127236 54372 127260 54374
rect 127316 54372 127340 54374
rect 127100 54352 127396 54372
rect 127100 53340 127396 53360
rect 127156 53338 127180 53340
rect 127236 53338 127260 53340
rect 127316 53338 127340 53340
rect 127178 53286 127180 53338
rect 127242 53286 127254 53338
rect 127316 53286 127318 53338
rect 127156 53284 127180 53286
rect 127236 53284 127260 53286
rect 127316 53284 127340 53286
rect 127100 53264 127396 53284
rect 127100 52252 127396 52272
rect 127156 52250 127180 52252
rect 127236 52250 127260 52252
rect 127316 52250 127340 52252
rect 127178 52198 127180 52250
rect 127242 52198 127254 52250
rect 127316 52198 127318 52250
rect 127156 52196 127180 52198
rect 127236 52196 127260 52198
rect 127316 52196 127340 52198
rect 127100 52176 127396 52196
rect 127100 51164 127396 51184
rect 127156 51162 127180 51164
rect 127236 51162 127260 51164
rect 127316 51162 127340 51164
rect 127178 51110 127180 51162
rect 127242 51110 127254 51162
rect 127316 51110 127318 51162
rect 127156 51108 127180 51110
rect 127236 51108 127260 51110
rect 127316 51108 127340 51110
rect 127100 51088 127396 51108
rect 127100 50076 127396 50096
rect 127156 50074 127180 50076
rect 127236 50074 127260 50076
rect 127316 50074 127340 50076
rect 127178 50022 127180 50074
rect 127242 50022 127254 50074
rect 127316 50022 127318 50074
rect 127156 50020 127180 50022
rect 127236 50020 127260 50022
rect 127316 50020 127340 50022
rect 127100 50000 127396 50020
rect 127100 48988 127396 49008
rect 127156 48986 127180 48988
rect 127236 48986 127260 48988
rect 127316 48986 127340 48988
rect 127178 48934 127180 48986
rect 127242 48934 127254 48986
rect 127316 48934 127318 48986
rect 127156 48932 127180 48934
rect 127236 48932 127260 48934
rect 127316 48932 127340 48934
rect 127100 48912 127396 48932
rect 127100 47900 127396 47920
rect 127156 47898 127180 47900
rect 127236 47898 127260 47900
rect 127316 47898 127340 47900
rect 127178 47846 127180 47898
rect 127242 47846 127254 47898
rect 127316 47846 127318 47898
rect 127156 47844 127180 47846
rect 127236 47844 127260 47846
rect 127316 47844 127340 47846
rect 127100 47824 127396 47844
rect 127100 46812 127396 46832
rect 127156 46810 127180 46812
rect 127236 46810 127260 46812
rect 127316 46810 127340 46812
rect 127178 46758 127180 46810
rect 127242 46758 127254 46810
rect 127316 46758 127318 46810
rect 127156 46756 127180 46758
rect 127236 46756 127260 46758
rect 127316 46756 127340 46758
rect 127100 46736 127396 46756
rect 127100 45724 127396 45744
rect 127156 45722 127180 45724
rect 127236 45722 127260 45724
rect 127316 45722 127340 45724
rect 127178 45670 127180 45722
rect 127242 45670 127254 45722
rect 127316 45670 127318 45722
rect 127156 45668 127180 45670
rect 127236 45668 127260 45670
rect 127316 45668 127340 45670
rect 127100 45648 127396 45668
rect 127100 44636 127396 44656
rect 127156 44634 127180 44636
rect 127236 44634 127260 44636
rect 127316 44634 127340 44636
rect 127178 44582 127180 44634
rect 127242 44582 127254 44634
rect 127316 44582 127318 44634
rect 127156 44580 127180 44582
rect 127236 44580 127260 44582
rect 127316 44580 127340 44582
rect 127100 44560 127396 44580
rect 127100 43548 127396 43568
rect 127156 43546 127180 43548
rect 127236 43546 127260 43548
rect 127316 43546 127340 43548
rect 127178 43494 127180 43546
rect 127242 43494 127254 43546
rect 127316 43494 127318 43546
rect 127156 43492 127180 43494
rect 127236 43492 127260 43494
rect 127316 43492 127340 43494
rect 127100 43472 127396 43492
rect 127100 42460 127396 42480
rect 127156 42458 127180 42460
rect 127236 42458 127260 42460
rect 127316 42458 127340 42460
rect 127178 42406 127180 42458
rect 127242 42406 127254 42458
rect 127316 42406 127318 42458
rect 127156 42404 127180 42406
rect 127236 42404 127260 42406
rect 127316 42404 127340 42406
rect 127100 42384 127396 42404
rect 127100 41372 127396 41392
rect 127156 41370 127180 41372
rect 127236 41370 127260 41372
rect 127316 41370 127340 41372
rect 127178 41318 127180 41370
rect 127242 41318 127254 41370
rect 127316 41318 127318 41370
rect 127156 41316 127180 41318
rect 127236 41316 127260 41318
rect 127316 41316 127340 41318
rect 127100 41296 127396 41316
rect 127100 40284 127396 40304
rect 127156 40282 127180 40284
rect 127236 40282 127260 40284
rect 127316 40282 127340 40284
rect 127178 40230 127180 40282
rect 127242 40230 127254 40282
rect 127316 40230 127318 40282
rect 127156 40228 127180 40230
rect 127236 40228 127260 40230
rect 127316 40228 127340 40230
rect 127100 40208 127396 40228
rect 127100 39196 127396 39216
rect 127156 39194 127180 39196
rect 127236 39194 127260 39196
rect 127316 39194 127340 39196
rect 127178 39142 127180 39194
rect 127242 39142 127254 39194
rect 127316 39142 127318 39194
rect 127156 39140 127180 39142
rect 127236 39140 127260 39142
rect 127316 39140 127340 39142
rect 127100 39120 127396 39140
rect 127100 38108 127396 38128
rect 127156 38106 127180 38108
rect 127236 38106 127260 38108
rect 127316 38106 127340 38108
rect 127178 38054 127180 38106
rect 127242 38054 127254 38106
rect 127316 38054 127318 38106
rect 127156 38052 127180 38054
rect 127236 38052 127260 38054
rect 127316 38052 127340 38054
rect 127100 38032 127396 38052
rect 127100 37020 127396 37040
rect 127156 37018 127180 37020
rect 127236 37018 127260 37020
rect 127316 37018 127340 37020
rect 127178 36966 127180 37018
rect 127242 36966 127254 37018
rect 127316 36966 127318 37018
rect 127156 36964 127180 36966
rect 127236 36964 127260 36966
rect 127316 36964 127340 36966
rect 127100 36944 127396 36964
rect 127100 35932 127396 35952
rect 127156 35930 127180 35932
rect 127236 35930 127260 35932
rect 127316 35930 127340 35932
rect 127178 35878 127180 35930
rect 127242 35878 127254 35930
rect 127316 35878 127318 35930
rect 127156 35876 127180 35878
rect 127236 35876 127260 35878
rect 127316 35876 127340 35878
rect 127100 35856 127396 35876
rect 127100 34844 127396 34864
rect 127156 34842 127180 34844
rect 127236 34842 127260 34844
rect 127316 34842 127340 34844
rect 127178 34790 127180 34842
rect 127242 34790 127254 34842
rect 127316 34790 127318 34842
rect 127156 34788 127180 34790
rect 127236 34788 127260 34790
rect 127316 34788 127340 34790
rect 127100 34768 127396 34788
rect 127100 33756 127396 33776
rect 127156 33754 127180 33756
rect 127236 33754 127260 33756
rect 127316 33754 127340 33756
rect 127178 33702 127180 33754
rect 127242 33702 127254 33754
rect 127316 33702 127318 33754
rect 127156 33700 127180 33702
rect 127236 33700 127260 33702
rect 127316 33700 127340 33702
rect 127100 33680 127396 33700
rect 127100 32668 127396 32688
rect 127156 32666 127180 32668
rect 127236 32666 127260 32668
rect 127316 32666 127340 32668
rect 127178 32614 127180 32666
rect 127242 32614 127254 32666
rect 127316 32614 127318 32666
rect 127156 32612 127180 32614
rect 127236 32612 127260 32614
rect 127316 32612 127340 32614
rect 127100 32592 127396 32612
rect 127100 31580 127396 31600
rect 127156 31578 127180 31580
rect 127236 31578 127260 31580
rect 127316 31578 127340 31580
rect 127178 31526 127180 31578
rect 127242 31526 127254 31578
rect 127316 31526 127318 31578
rect 127156 31524 127180 31526
rect 127236 31524 127260 31526
rect 127316 31524 127340 31526
rect 127100 31504 127396 31524
rect 127100 30492 127396 30512
rect 127156 30490 127180 30492
rect 127236 30490 127260 30492
rect 127316 30490 127340 30492
rect 127178 30438 127180 30490
rect 127242 30438 127254 30490
rect 127316 30438 127318 30490
rect 127156 30436 127180 30438
rect 127236 30436 127260 30438
rect 127316 30436 127340 30438
rect 127100 30416 127396 30436
rect 127100 29404 127396 29424
rect 127156 29402 127180 29404
rect 127236 29402 127260 29404
rect 127316 29402 127340 29404
rect 127178 29350 127180 29402
rect 127242 29350 127254 29402
rect 127316 29350 127318 29402
rect 127156 29348 127180 29350
rect 127236 29348 127260 29350
rect 127316 29348 127340 29350
rect 127100 29328 127396 29348
rect 127100 28316 127396 28336
rect 127156 28314 127180 28316
rect 127236 28314 127260 28316
rect 127316 28314 127340 28316
rect 127178 28262 127180 28314
rect 127242 28262 127254 28314
rect 127316 28262 127318 28314
rect 127156 28260 127180 28262
rect 127236 28260 127260 28262
rect 127316 28260 127340 28262
rect 127100 28240 127396 28260
rect 127100 27228 127396 27248
rect 127156 27226 127180 27228
rect 127236 27226 127260 27228
rect 127316 27226 127340 27228
rect 127178 27174 127180 27226
rect 127242 27174 127254 27226
rect 127316 27174 127318 27226
rect 127156 27172 127180 27174
rect 127236 27172 127260 27174
rect 127316 27172 127340 27174
rect 127100 27152 127396 27172
rect 127100 26140 127396 26160
rect 127156 26138 127180 26140
rect 127236 26138 127260 26140
rect 127316 26138 127340 26140
rect 127178 26086 127180 26138
rect 127242 26086 127254 26138
rect 127316 26086 127318 26138
rect 127156 26084 127180 26086
rect 127236 26084 127260 26086
rect 127316 26084 127340 26086
rect 127100 26064 127396 26084
rect 127100 25052 127396 25072
rect 127156 25050 127180 25052
rect 127236 25050 127260 25052
rect 127316 25050 127340 25052
rect 127178 24998 127180 25050
rect 127242 24998 127254 25050
rect 127316 24998 127318 25050
rect 127156 24996 127180 24998
rect 127236 24996 127260 24998
rect 127316 24996 127340 24998
rect 127100 24976 127396 24996
rect 127100 23964 127396 23984
rect 127156 23962 127180 23964
rect 127236 23962 127260 23964
rect 127316 23962 127340 23964
rect 127178 23910 127180 23962
rect 127242 23910 127254 23962
rect 127316 23910 127318 23962
rect 127156 23908 127180 23910
rect 127236 23908 127260 23910
rect 127316 23908 127340 23910
rect 127100 23888 127396 23908
rect 127100 22876 127396 22896
rect 127156 22874 127180 22876
rect 127236 22874 127260 22876
rect 127316 22874 127340 22876
rect 127178 22822 127180 22874
rect 127242 22822 127254 22874
rect 127316 22822 127318 22874
rect 127156 22820 127180 22822
rect 127236 22820 127260 22822
rect 127316 22820 127340 22822
rect 127100 22800 127396 22820
rect 127100 21788 127396 21808
rect 127156 21786 127180 21788
rect 127236 21786 127260 21788
rect 127316 21786 127340 21788
rect 127178 21734 127180 21786
rect 127242 21734 127254 21786
rect 127316 21734 127318 21786
rect 127156 21732 127180 21734
rect 127236 21732 127260 21734
rect 127316 21732 127340 21734
rect 127100 21712 127396 21732
rect 127100 20700 127396 20720
rect 127156 20698 127180 20700
rect 127236 20698 127260 20700
rect 127316 20698 127340 20700
rect 127178 20646 127180 20698
rect 127242 20646 127254 20698
rect 127316 20646 127318 20698
rect 127156 20644 127180 20646
rect 127236 20644 127260 20646
rect 127316 20644 127340 20646
rect 127100 20624 127396 20644
rect 121736 20052 121788 20058
rect 121736 19994 121788 20000
rect 130764 19990 130792 117098
rect 133524 116346 133552 117098
rect 133512 116340 133564 116346
rect 133512 116282 133564 116288
rect 130752 19984 130804 19990
rect 130752 19926 130804 19932
rect 96380 19612 96676 19632
rect 96436 19610 96460 19612
rect 96516 19610 96540 19612
rect 96596 19610 96620 19612
rect 96458 19558 96460 19610
rect 96522 19558 96534 19610
rect 96596 19558 96598 19610
rect 96436 19556 96460 19558
rect 96516 19556 96540 19558
rect 96596 19556 96620 19558
rect 96380 19536 96676 19556
rect 127100 19612 127396 19632
rect 127156 19610 127180 19612
rect 127236 19610 127260 19612
rect 127316 19610 127340 19612
rect 127178 19558 127180 19610
rect 127242 19558 127254 19610
rect 127316 19558 127318 19610
rect 127156 19556 127180 19558
rect 127236 19556 127260 19558
rect 127316 19556 127340 19558
rect 127100 19536 127396 19556
rect 135456 19514 135484 117098
rect 138032 116346 138060 117098
rect 138020 116340 138072 116346
rect 138020 116282 138072 116288
rect 135444 19508 135496 19514
rect 135444 19450 135496 19456
rect 140424 19174 140452 117098
rect 142460 116988 142756 117008
rect 142516 116986 142540 116988
rect 142596 116986 142620 116988
rect 142676 116986 142700 116988
rect 142538 116934 142540 116986
rect 142602 116934 142614 116986
rect 142676 116934 142678 116986
rect 142516 116932 142540 116934
rect 142596 116932 142620 116934
rect 142676 116932 142700 116934
rect 142460 116912 142756 116932
rect 143184 116346 143212 117098
rect 143172 116340 143224 116346
rect 143172 116282 143224 116288
rect 142460 115900 142756 115920
rect 142516 115898 142540 115900
rect 142596 115898 142620 115900
rect 142676 115898 142700 115900
rect 142538 115846 142540 115898
rect 142602 115846 142614 115898
rect 142676 115846 142678 115898
rect 142516 115844 142540 115846
rect 142596 115844 142620 115846
rect 142676 115844 142700 115846
rect 142460 115824 142756 115844
rect 142460 114812 142756 114832
rect 142516 114810 142540 114812
rect 142596 114810 142620 114812
rect 142676 114810 142700 114812
rect 142538 114758 142540 114810
rect 142602 114758 142614 114810
rect 142676 114758 142678 114810
rect 142516 114756 142540 114758
rect 142596 114756 142620 114758
rect 142676 114756 142700 114758
rect 142460 114736 142756 114756
rect 142460 113724 142756 113744
rect 142516 113722 142540 113724
rect 142596 113722 142620 113724
rect 142676 113722 142700 113724
rect 142538 113670 142540 113722
rect 142602 113670 142614 113722
rect 142676 113670 142678 113722
rect 142516 113668 142540 113670
rect 142596 113668 142620 113670
rect 142676 113668 142700 113670
rect 142460 113648 142756 113668
rect 142460 112636 142756 112656
rect 142516 112634 142540 112636
rect 142596 112634 142620 112636
rect 142676 112634 142700 112636
rect 142538 112582 142540 112634
rect 142602 112582 142614 112634
rect 142676 112582 142678 112634
rect 142516 112580 142540 112582
rect 142596 112580 142620 112582
rect 142676 112580 142700 112582
rect 142460 112560 142756 112580
rect 142460 111548 142756 111568
rect 142516 111546 142540 111548
rect 142596 111546 142620 111548
rect 142676 111546 142700 111548
rect 142538 111494 142540 111546
rect 142602 111494 142614 111546
rect 142676 111494 142678 111546
rect 142516 111492 142540 111494
rect 142596 111492 142620 111494
rect 142676 111492 142700 111494
rect 142460 111472 142756 111492
rect 142460 110460 142756 110480
rect 142516 110458 142540 110460
rect 142596 110458 142620 110460
rect 142676 110458 142700 110460
rect 142538 110406 142540 110458
rect 142602 110406 142614 110458
rect 142676 110406 142678 110458
rect 142516 110404 142540 110406
rect 142596 110404 142620 110406
rect 142676 110404 142700 110406
rect 142460 110384 142756 110404
rect 142460 109372 142756 109392
rect 142516 109370 142540 109372
rect 142596 109370 142620 109372
rect 142676 109370 142700 109372
rect 142538 109318 142540 109370
rect 142602 109318 142614 109370
rect 142676 109318 142678 109370
rect 142516 109316 142540 109318
rect 142596 109316 142620 109318
rect 142676 109316 142700 109318
rect 142460 109296 142756 109316
rect 142460 108284 142756 108304
rect 142516 108282 142540 108284
rect 142596 108282 142620 108284
rect 142676 108282 142700 108284
rect 142538 108230 142540 108282
rect 142602 108230 142614 108282
rect 142676 108230 142678 108282
rect 142516 108228 142540 108230
rect 142596 108228 142620 108230
rect 142676 108228 142700 108230
rect 142460 108208 142756 108228
rect 142460 107196 142756 107216
rect 142516 107194 142540 107196
rect 142596 107194 142620 107196
rect 142676 107194 142700 107196
rect 142538 107142 142540 107194
rect 142602 107142 142614 107194
rect 142676 107142 142678 107194
rect 142516 107140 142540 107142
rect 142596 107140 142620 107142
rect 142676 107140 142700 107142
rect 142460 107120 142756 107140
rect 142460 106108 142756 106128
rect 142516 106106 142540 106108
rect 142596 106106 142620 106108
rect 142676 106106 142700 106108
rect 142538 106054 142540 106106
rect 142602 106054 142614 106106
rect 142676 106054 142678 106106
rect 142516 106052 142540 106054
rect 142596 106052 142620 106054
rect 142676 106052 142700 106054
rect 142460 106032 142756 106052
rect 142460 105020 142756 105040
rect 142516 105018 142540 105020
rect 142596 105018 142620 105020
rect 142676 105018 142700 105020
rect 142538 104966 142540 105018
rect 142602 104966 142614 105018
rect 142676 104966 142678 105018
rect 142516 104964 142540 104966
rect 142596 104964 142620 104966
rect 142676 104964 142700 104966
rect 142460 104944 142756 104964
rect 142460 103932 142756 103952
rect 142516 103930 142540 103932
rect 142596 103930 142620 103932
rect 142676 103930 142700 103932
rect 142538 103878 142540 103930
rect 142602 103878 142614 103930
rect 142676 103878 142678 103930
rect 142516 103876 142540 103878
rect 142596 103876 142620 103878
rect 142676 103876 142700 103878
rect 142460 103856 142756 103876
rect 142460 102844 142756 102864
rect 142516 102842 142540 102844
rect 142596 102842 142620 102844
rect 142676 102842 142700 102844
rect 142538 102790 142540 102842
rect 142602 102790 142614 102842
rect 142676 102790 142678 102842
rect 142516 102788 142540 102790
rect 142596 102788 142620 102790
rect 142676 102788 142700 102790
rect 142460 102768 142756 102788
rect 142460 101756 142756 101776
rect 142516 101754 142540 101756
rect 142596 101754 142620 101756
rect 142676 101754 142700 101756
rect 142538 101702 142540 101754
rect 142602 101702 142614 101754
rect 142676 101702 142678 101754
rect 142516 101700 142540 101702
rect 142596 101700 142620 101702
rect 142676 101700 142700 101702
rect 142460 101680 142756 101700
rect 142460 100668 142756 100688
rect 142516 100666 142540 100668
rect 142596 100666 142620 100668
rect 142676 100666 142700 100668
rect 142538 100614 142540 100666
rect 142602 100614 142614 100666
rect 142676 100614 142678 100666
rect 142516 100612 142540 100614
rect 142596 100612 142620 100614
rect 142676 100612 142700 100614
rect 142460 100592 142756 100612
rect 142460 99580 142756 99600
rect 142516 99578 142540 99580
rect 142596 99578 142620 99580
rect 142676 99578 142700 99580
rect 142538 99526 142540 99578
rect 142602 99526 142614 99578
rect 142676 99526 142678 99578
rect 142516 99524 142540 99526
rect 142596 99524 142620 99526
rect 142676 99524 142700 99526
rect 142460 99504 142756 99524
rect 142460 98492 142756 98512
rect 142516 98490 142540 98492
rect 142596 98490 142620 98492
rect 142676 98490 142700 98492
rect 142538 98438 142540 98490
rect 142602 98438 142614 98490
rect 142676 98438 142678 98490
rect 142516 98436 142540 98438
rect 142596 98436 142620 98438
rect 142676 98436 142700 98438
rect 142460 98416 142756 98436
rect 142460 97404 142756 97424
rect 142516 97402 142540 97404
rect 142596 97402 142620 97404
rect 142676 97402 142700 97404
rect 142538 97350 142540 97402
rect 142602 97350 142614 97402
rect 142676 97350 142678 97402
rect 142516 97348 142540 97350
rect 142596 97348 142620 97350
rect 142676 97348 142700 97350
rect 142460 97328 142756 97348
rect 142460 96316 142756 96336
rect 142516 96314 142540 96316
rect 142596 96314 142620 96316
rect 142676 96314 142700 96316
rect 142538 96262 142540 96314
rect 142602 96262 142614 96314
rect 142676 96262 142678 96314
rect 142516 96260 142540 96262
rect 142596 96260 142620 96262
rect 142676 96260 142700 96262
rect 142460 96240 142756 96260
rect 142460 95228 142756 95248
rect 142516 95226 142540 95228
rect 142596 95226 142620 95228
rect 142676 95226 142700 95228
rect 142538 95174 142540 95226
rect 142602 95174 142614 95226
rect 142676 95174 142678 95226
rect 142516 95172 142540 95174
rect 142596 95172 142620 95174
rect 142676 95172 142700 95174
rect 142460 95152 142756 95172
rect 142460 94140 142756 94160
rect 142516 94138 142540 94140
rect 142596 94138 142620 94140
rect 142676 94138 142700 94140
rect 142538 94086 142540 94138
rect 142602 94086 142614 94138
rect 142676 94086 142678 94138
rect 142516 94084 142540 94086
rect 142596 94084 142620 94086
rect 142676 94084 142700 94086
rect 142460 94064 142756 94084
rect 142460 93052 142756 93072
rect 142516 93050 142540 93052
rect 142596 93050 142620 93052
rect 142676 93050 142700 93052
rect 142538 92998 142540 93050
rect 142602 92998 142614 93050
rect 142676 92998 142678 93050
rect 142516 92996 142540 92998
rect 142596 92996 142620 92998
rect 142676 92996 142700 92998
rect 142460 92976 142756 92996
rect 142460 91964 142756 91984
rect 142516 91962 142540 91964
rect 142596 91962 142620 91964
rect 142676 91962 142700 91964
rect 142538 91910 142540 91962
rect 142602 91910 142614 91962
rect 142676 91910 142678 91962
rect 142516 91908 142540 91910
rect 142596 91908 142620 91910
rect 142676 91908 142700 91910
rect 142460 91888 142756 91908
rect 142460 90876 142756 90896
rect 142516 90874 142540 90876
rect 142596 90874 142620 90876
rect 142676 90874 142700 90876
rect 142538 90822 142540 90874
rect 142602 90822 142614 90874
rect 142676 90822 142678 90874
rect 142516 90820 142540 90822
rect 142596 90820 142620 90822
rect 142676 90820 142700 90822
rect 142460 90800 142756 90820
rect 142460 89788 142756 89808
rect 142516 89786 142540 89788
rect 142596 89786 142620 89788
rect 142676 89786 142700 89788
rect 142538 89734 142540 89786
rect 142602 89734 142614 89786
rect 142676 89734 142678 89786
rect 142516 89732 142540 89734
rect 142596 89732 142620 89734
rect 142676 89732 142700 89734
rect 142460 89712 142756 89732
rect 142460 88700 142756 88720
rect 142516 88698 142540 88700
rect 142596 88698 142620 88700
rect 142676 88698 142700 88700
rect 142538 88646 142540 88698
rect 142602 88646 142614 88698
rect 142676 88646 142678 88698
rect 142516 88644 142540 88646
rect 142596 88644 142620 88646
rect 142676 88644 142700 88646
rect 142460 88624 142756 88644
rect 142460 87612 142756 87632
rect 142516 87610 142540 87612
rect 142596 87610 142620 87612
rect 142676 87610 142700 87612
rect 142538 87558 142540 87610
rect 142602 87558 142614 87610
rect 142676 87558 142678 87610
rect 142516 87556 142540 87558
rect 142596 87556 142620 87558
rect 142676 87556 142700 87558
rect 142460 87536 142756 87556
rect 142460 86524 142756 86544
rect 142516 86522 142540 86524
rect 142596 86522 142620 86524
rect 142676 86522 142700 86524
rect 142538 86470 142540 86522
rect 142602 86470 142614 86522
rect 142676 86470 142678 86522
rect 142516 86468 142540 86470
rect 142596 86468 142620 86470
rect 142676 86468 142700 86470
rect 142460 86448 142756 86468
rect 142460 85436 142756 85456
rect 142516 85434 142540 85436
rect 142596 85434 142620 85436
rect 142676 85434 142700 85436
rect 142538 85382 142540 85434
rect 142602 85382 142614 85434
rect 142676 85382 142678 85434
rect 142516 85380 142540 85382
rect 142596 85380 142620 85382
rect 142676 85380 142700 85382
rect 142460 85360 142756 85380
rect 142460 84348 142756 84368
rect 142516 84346 142540 84348
rect 142596 84346 142620 84348
rect 142676 84346 142700 84348
rect 142538 84294 142540 84346
rect 142602 84294 142614 84346
rect 142676 84294 142678 84346
rect 142516 84292 142540 84294
rect 142596 84292 142620 84294
rect 142676 84292 142700 84294
rect 142460 84272 142756 84292
rect 142460 83260 142756 83280
rect 142516 83258 142540 83260
rect 142596 83258 142620 83260
rect 142676 83258 142700 83260
rect 142538 83206 142540 83258
rect 142602 83206 142614 83258
rect 142676 83206 142678 83258
rect 142516 83204 142540 83206
rect 142596 83204 142620 83206
rect 142676 83204 142700 83206
rect 142460 83184 142756 83204
rect 142460 82172 142756 82192
rect 142516 82170 142540 82172
rect 142596 82170 142620 82172
rect 142676 82170 142700 82172
rect 142538 82118 142540 82170
rect 142602 82118 142614 82170
rect 142676 82118 142678 82170
rect 142516 82116 142540 82118
rect 142596 82116 142620 82118
rect 142676 82116 142700 82118
rect 142460 82096 142756 82116
rect 142460 81084 142756 81104
rect 142516 81082 142540 81084
rect 142596 81082 142620 81084
rect 142676 81082 142700 81084
rect 142538 81030 142540 81082
rect 142602 81030 142614 81082
rect 142676 81030 142678 81082
rect 142516 81028 142540 81030
rect 142596 81028 142620 81030
rect 142676 81028 142700 81030
rect 142460 81008 142756 81028
rect 142460 79996 142756 80016
rect 142516 79994 142540 79996
rect 142596 79994 142620 79996
rect 142676 79994 142700 79996
rect 142538 79942 142540 79994
rect 142602 79942 142614 79994
rect 142676 79942 142678 79994
rect 142516 79940 142540 79942
rect 142596 79940 142620 79942
rect 142676 79940 142700 79942
rect 142460 79920 142756 79940
rect 142460 78908 142756 78928
rect 142516 78906 142540 78908
rect 142596 78906 142620 78908
rect 142676 78906 142700 78908
rect 142538 78854 142540 78906
rect 142602 78854 142614 78906
rect 142676 78854 142678 78906
rect 142516 78852 142540 78854
rect 142596 78852 142620 78854
rect 142676 78852 142700 78854
rect 142460 78832 142756 78852
rect 142460 77820 142756 77840
rect 142516 77818 142540 77820
rect 142596 77818 142620 77820
rect 142676 77818 142700 77820
rect 142538 77766 142540 77818
rect 142602 77766 142614 77818
rect 142676 77766 142678 77818
rect 142516 77764 142540 77766
rect 142596 77764 142620 77766
rect 142676 77764 142700 77766
rect 142460 77744 142756 77764
rect 142460 76732 142756 76752
rect 142516 76730 142540 76732
rect 142596 76730 142620 76732
rect 142676 76730 142700 76732
rect 142538 76678 142540 76730
rect 142602 76678 142614 76730
rect 142676 76678 142678 76730
rect 142516 76676 142540 76678
rect 142596 76676 142620 76678
rect 142676 76676 142700 76678
rect 142460 76656 142756 76676
rect 142460 75644 142756 75664
rect 142516 75642 142540 75644
rect 142596 75642 142620 75644
rect 142676 75642 142700 75644
rect 142538 75590 142540 75642
rect 142602 75590 142614 75642
rect 142676 75590 142678 75642
rect 142516 75588 142540 75590
rect 142596 75588 142620 75590
rect 142676 75588 142700 75590
rect 142460 75568 142756 75588
rect 142460 74556 142756 74576
rect 142516 74554 142540 74556
rect 142596 74554 142620 74556
rect 142676 74554 142700 74556
rect 142538 74502 142540 74554
rect 142602 74502 142614 74554
rect 142676 74502 142678 74554
rect 142516 74500 142540 74502
rect 142596 74500 142620 74502
rect 142676 74500 142700 74502
rect 142460 74480 142756 74500
rect 142460 73468 142756 73488
rect 142516 73466 142540 73468
rect 142596 73466 142620 73468
rect 142676 73466 142700 73468
rect 142538 73414 142540 73466
rect 142602 73414 142614 73466
rect 142676 73414 142678 73466
rect 142516 73412 142540 73414
rect 142596 73412 142620 73414
rect 142676 73412 142700 73414
rect 142460 73392 142756 73412
rect 142460 72380 142756 72400
rect 142516 72378 142540 72380
rect 142596 72378 142620 72380
rect 142676 72378 142700 72380
rect 142538 72326 142540 72378
rect 142602 72326 142614 72378
rect 142676 72326 142678 72378
rect 142516 72324 142540 72326
rect 142596 72324 142620 72326
rect 142676 72324 142700 72326
rect 142460 72304 142756 72324
rect 142460 71292 142756 71312
rect 142516 71290 142540 71292
rect 142596 71290 142620 71292
rect 142676 71290 142700 71292
rect 142538 71238 142540 71290
rect 142602 71238 142614 71290
rect 142676 71238 142678 71290
rect 142516 71236 142540 71238
rect 142596 71236 142620 71238
rect 142676 71236 142700 71238
rect 142460 71216 142756 71236
rect 142460 70204 142756 70224
rect 142516 70202 142540 70204
rect 142596 70202 142620 70204
rect 142676 70202 142700 70204
rect 142538 70150 142540 70202
rect 142602 70150 142614 70202
rect 142676 70150 142678 70202
rect 142516 70148 142540 70150
rect 142596 70148 142620 70150
rect 142676 70148 142700 70150
rect 142460 70128 142756 70148
rect 142460 69116 142756 69136
rect 142516 69114 142540 69116
rect 142596 69114 142620 69116
rect 142676 69114 142700 69116
rect 142538 69062 142540 69114
rect 142602 69062 142614 69114
rect 142676 69062 142678 69114
rect 142516 69060 142540 69062
rect 142596 69060 142620 69062
rect 142676 69060 142700 69062
rect 142460 69040 142756 69060
rect 142460 68028 142756 68048
rect 142516 68026 142540 68028
rect 142596 68026 142620 68028
rect 142676 68026 142700 68028
rect 142538 67974 142540 68026
rect 142602 67974 142614 68026
rect 142676 67974 142678 68026
rect 142516 67972 142540 67974
rect 142596 67972 142620 67974
rect 142676 67972 142700 67974
rect 142460 67952 142756 67972
rect 142460 66940 142756 66960
rect 142516 66938 142540 66940
rect 142596 66938 142620 66940
rect 142676 66938 142700 66940
rect 142538 66886 142540 66938
rect 142602 66886 142614 66938
rect 142676 66886 142678 66938
rect 142516 66884 142540 66886
rect 142596 66884 142620 66886
rect 142676 66884 142700 66886
rect 142460 66864 142756 66884
rect 142460 65852 142756 65872
rect 142516 65850 142540 65852
rect 142596 65850 142620 65852
rect 142676 65850 142700 65852
rect 142538 65798 142540 65850
rect 142602 65798 142614 65850
rect 142676 65798 142678 65850
rect 142516 65796 142540 65798
rect 142596 65796 142620 65798
rect 142676 65796 142700 65798
rect 142460 65776 142756 65796
rect 142460 64764 142756 64784
rect 142516 64762 142540 64764
rect 142596 64762 142620 64764
rect 142676 64762 142700 64764
rect 142538 64710 142540 64762
rect 142602 64710 142614 64762
rect 142676 64710 142678 64762
rect 142516 64708 142540 64710
rect 142596 64708 142620 64710
rect 142676 64708 142700 64710
rect 142460 64688 142756 64708
rect 142460 63676 142756 63696
rect 142516 63674 142540 63676
rect 142596 63674 142620 63676
rect 142676 63674 142700 63676
rect 142538 63622 142540 63674
rect 142602 63622 142614 63674
rect 142676 63622 142678 63674
rect 142516 63620 142540 63622
rect 142596 63620 142620 63622
rect 142676 63620 142700 63622
rect 142460 63600 142756 63620
rect 142460 62588 142756 62608
rect 142516 62586 142540 62588
rect 142596 62586 142620 62588
rect 142676 62586 142700 62588
rect 142538 62534 142540 62586
rect 142602 62534 142614 62586
rect 142676 62534 142678 62586
rect 142516 62532 142540 62534
rect 142596 62532 142620 62534
rect 142676 62532 142700 62534
rect 142460 62512 142756 62532
rect 142460 61500 142756 61520
rect 142516 61498 142540 61500
rect 142596 61498 142620 61500
rect 142676 61498 142700 61500
rect 142538 61446 142540 61498
rect 142602 61446 142614 61498
rect 142676 61446 142678 61498
rect 142516 61444 142540 61446
rect 142596 61444 142620 61446
rect 142676 61444 142700 61446
rect 142460 61424 142756 61444
rect 142460 60412 142756 60432
rect 142516 60410 142540 60412
rect 142596 60410 142620 60412
rect 142676 60410 142700 60412
rect 142538 60358 142540 60410
rect 142602 60358 142614 60410
rect 142676 60358 142678 60410
rect 142516 60356 142540 60358
rect 142596 60356 142620 60358
rect 142676 60356 142700 60358
rect 142460 60336 142756 60356
rect 142460 59324 142756 59344
rect 142516 59322 142540 59324
rect 142596 59322 142620 59324
rect 142676 59322 142700 59324
rect 142538 59270 142540 59322
rect 142602 59270 142614 59322
rect 142676 59270 142678 59322
rect 142516 59268 142540 59270
rect 142596 59268 142620 59270
rect 142676 59268 142700 59270
rect 142460 59248 142756 59268
rect 142460 58236 142756 58256
rect 142516 58234 142540 58236
rect 142596 58234 142620 58236
rect 142676 58234 142700 58236
rect 142538 58182 142540 58234
rect 142602 58182 142614 58234
rect 142676 58182 142678 58234
rect 142516 58180 142540 58182
rect 142596 58180 142620 58182
rect 142676 58180 142700 58182
rect 142460 58160 142756 58180
rect 142460 57148 142756 57168
rect 142516 57146 142540 57148
rect 142596 57146 142620 57148
rect 142676 57146 142700 57148
rect 142538 57094 142540 57146
rect 142602 57094 142614 57146
rect 142676 57094 142678 57146
rect 142516 57092 142540 57094
rect 142596 57092 142620 57094
rect 142676 57092 142700 57094
rect 142460 57072 142756 57092
rect 142460 56060 142756 56080
rect 142516 56058 142540 56060
rect 142596 56058 142620 56060
rect 142676 56058 142700 56060
rect 142538 56006 142540 56058
rect 142602 56006 142614 56058
rect 142676 56006 142678 56058
rect 142516 56004 142540 56006
rect 142596 56004 142620 56006
rect 142676 56004 142700 56006
rect 142460 55984 142756 56004
rect 142460 54972 142756 54992
rect 142516 54970 142540 54972
rect 142596 54970 142620 54972
rect 142676 54970 142700 54972
rect 142538 54918 142540 54970
rect 142602 54918 142614 54970
rect 142676 54918 142678 54970
rect 142516 54916 142540 54918
rect 142596 54916 142620 54918
rect 142676 54916 142700 54918
rect 142460 54896 142756 54916
rect 142460 53884 142756 53904
rect 142516 53882 142540 53884
rect 142596 53882 142620 53884
rect 142676 53882 142700 53884
rect 142538 53830 142540 53882
rect 142602 53830 142614 53882
rect 142676 53830 142678 53882
rect 142516 53828 142540 53830
rect 142596 53828 142620 53830
rect 142676 53828 142700 53830
rect 142460 53808 142756 53828
rect 142460 52796 142756 52816
rect 142516 52794 142540 52796
rect 142596 52794 142620 52796
rect 142676 52794 142700 52796
rect 142538 52742 142540 52794
rect 142602 52742 142614 52794
rect 142676 52742 142678 52794
rect 142516 52740 142540 52742
rect 142596 52740 142620 52742
rect 142676 52740 142700 52742
rect 142460 52720 142756 52740
rect 142460 51708 142756 51728
rect 142516 51706 142540 51708
rect 142596 51706 142620 51708
rect 142676 51706 142700 51708
rect 142538 51654 142540 51706
rect 142602 51654 142614 51706
rect 142676 51654 142678 51706
rect 142516 51652 142540 51654
rect 142596 51652 142620 51654
rect 142676 51652 142700 51654
rect 142460 51632 142756 51652
rect 142460 50620 142756 50640
rect 142516 50618 142540 50620
rect 142596 50618 142620 50620
rect 142676 50618 142700 50620
rect 142538 50566 142540 50618
rect 142602 50566 142614 50618
rect 142676 50566 142678 50618
rect 142516 50564 142540 50566
rect 142596 50564 142620 50566
rect 142676 50564 142700 50566
rect 142460 50544 142756 50564
rect 142460 49532 142756 49552
rect 142516 49530 142540 49532
rect 142596 49530 142620 49532
rect 142676 49530 142700 49532
rect 142538 49478 142540 49530
rect 142602 49478 142614 49530
rect 142676 49478 142678 49530
rect 142516 49476 142540 49478
rect 142596 49476 142620 49478
rect 142676 49476 142700 49478
rect 142460 49456 142756 49476
rect 142460 48444 142756 48464
rect 142516 48442 142540 48444
rect 142596 48442 142620 48444
rect 142676 48442 142700 48444
rect 142538 48390 142540 48442
rect 142602 48390 142614 48442
rect 142676 48390 142678 48442
rect 142516 48388 142540 48390
rect 142596 48388 142620 48390
rect 142676 48388 142700 48390
rect 142460 48368 142756 48388
rect 142460 47356 142756 47376
rect 142516 47354 142540 47356
rect 142596 47354 142620 47356
rect 142676 47354 142700 47356
rect 142538 47302 142540 47354
rect 142602 47302 142614 47354
rect 142676 47302 142678 47354
rect 142516 47300 142540 47302
rect 142596 47300 142620 47302
rect 142676 47300 142700 47302
rect 142460 47280 142756 47300
rect 142460 46268 142756 46288
rect 142516 46266 142540 46268
rect 142596 46266 142620 46268
rect 142676 46266 142700 46268
rect 142538 46214 142540 46266
rect 142602 46214 142614 46266
rect 142676 46214 142678 46266
rect 142516 46212 142540 46214
rect 142596 46212 142620 46214
rect 142676 46212 142700 46214
rect 142460 46192 142756 46212
rect 142460 45180 142756 45200
rect 142516 45178 142540 45180
rect 142596 45178 142620 45180
rect 142676 45178 142700 45180
rect 142538 45126 142540 45178
rect 142602 45126 142614 45178
rect 142676 45126 142678 45178
rect 142516 45124 142540 45126
rect 142596 45124 142620 45126
rect 142676 45124 142700 45126
rect 142460 45104 142756 45124
rect 142460 44092 142756 44112
rect 142516 44090 142540 44092
rect 142596 44090 142620 44092
rect 142676 44090 142700 44092
rect 142538 44038 142540 44090
rect 142602 44038 142614 44090
rect 142676 44038 142678 44090
rect 142516 44036 142540 44038
rect 142596 44036 142620 44038
rect 142676 44036 142700 44038
rect 142460 44016 142756 44036
rect 142460 43004 142756 43024
rect 142516 43002 142540 43004
rect 142596 43002 142620 43004
rect 142676 43002 142700 43004
rect 142538 42950 142540 43002
rect 142602 42950 142614 43002
rect 142676 42950 142678 43002
rect 142516 42948 142540 42950
rect 142596 42948 142620 42950
rect 142676 42948 142700 42950
rect 142460 42928 142756 42948
rect 142460 41916 142756 41936
rect 142516 41914 142540 41916
rect 142596 41914 142620 41916
rect 142676 41914 142700 41916
rect 142538 41862 142540 41914
rect 142602 41862 142614 41914
rect 142676 41862 142678 41914
rect 142516 41860 142540 41862
rect 142596 41860 142620 41862
rect 142676 41860 142700 41862
rect 142460 41840 142756 41860
rect 142460 40828 142756 40848
rect 142516 40826 142540 40828
rect 142596 40826 142620 40828
rect 142676 40826 142700 40828
rect 142538 40774 142540 40826
rect 142602 40774 142614 40826
rect 142676 40774 142678 40826
rect 142516 40772 142540 40774
rect 142596 40772 142620 40774
rect 142676 40772 142700 40774
rect 142460 40752 142756 40772
rect 142460 39740 142756 39760
rect 142516 39738 142540 39740
rect 142596 39738 142620 39740
rect 142676 39738 142700 39740
rect 142538 39686 142540 39738
rect 142602 39686 142614 39738
rect 142676 39686 142678 39738
rect 142516 39684 142540 39686
rect 142596 39684 142620 39686
rect 142676 39684 142700 39686
rect 142460 39664 142756 39684
rect 142460 38652 142756 38672
rect 142516 38650 142540 38652
rect 142596 38650 142620 38652
rect 142676 38650 142700 38652
rect 142538 38598 142540 38650
rect 142602 38598 142614 38650
rect 142676 38598 142678 38650
rect 142516 38596 142540 38598
rect 142596 38596 142620 38598
rect 142676 38596 142700 38598
rect 142460 38576 142756 38596
rect 142460 37564 142756 37584
rect 142516 37562 142540 37564
rect 142596 37562 142620 37564
rect 142676 37562 142700 37564
rect 142538 37510 142540 37562
rect 142602 37510 142614 37562
rect 142676 37510 142678 37562
rect 142516 37508 142540 37510
rect 142596 37508 142620 37510
rect 142676 37508 142700 37510
rect 142460 37488 142756 37508
rect 142460 36476 142756 36496
rect 142516 36474 142540 36476
rect 142596 36474 142620 36476
rect 142676 36474 142700 36476
rect 142538 36422 142540 36474
rect 142602 36422 142614 36474
rect 142676 36422 142678 36474
rect 142516 36420 142540 36422
rect 142596 36420 142620 36422
rect 142676 36420 142700 36422
rect 142460 36400 142756 36420
rect 142460 35388 142756 35408
rect 142516 35386 142540 35388
rect 142596 35386 142620 35388
rect 142676 35386 142700 35388
rect 142538 35334 142540 35386
rect 142602 35334 142614 35386
rect 142676 35334 142678 35386
rect 142516 35332 142540 35334
rect 142596 35332 142620 35334
rect 142676 35332 142700 35334
rect 142460 35312 142756 35332
rect 142460 34300 142756 34320
rect 142516 34298 142540 34300
rect 142596 34298 142620 34300
rect 142676 34298 142700 34300
rect 142538 34246 142540 34298
rect 142602 34246 142614 34298
rect 142676 34246 142678 34298
rect 142516 34244 142540 34246
rect 142596 34244 142620 34246
rect 142676 34244 142700 34246
rect 142460 34224 142756 34244
rect 142460 33212 142756 33232
rect 142516 33210 142540 33212
rect 142596 33210 142620 33212
rect 142676 33210 142700 33212
rect 142538 33158 142540 33210
rect 142602 33158 142614 33210
rect 142676 33158 142678 33210
rect 142516 33156 142540 33158
rect 142596 33156 142620 33158
rect 142676 33156 142700 33158
rect 142460 33136 142756 33156
rect 142460 32124 142756 32144
rect 142516 32122 142540 32124
rect 142596 32122 142620 32124
rect 142676 32122 142700 32124
rect 142538 32070 142540 32122
rect 142602 32070 142614 32122
rect 142676 32070 142678 32122
rect 142516 32068 142540 32070
rect 142596 32068 142620 32070
rect 142676 32068 142700 32070
rect 142460 32048 142756 32068
rect 142460 31036 142756 31056
rect 142516 31034 142540 31036
rect 142596 31034 142620 31036
rect 142676 31034 142700 31036
rect 142538 30982 142540 31034
rect 142602 30982 142614 31034
rect 142676 30982 142678 31034
rect 142516 30980 142540 30982
rect 142596 30980 142620 30982
rect 142676 30980 142700 30982
rect 142460 30960 142756 30980
rect 142460 29948 142756 29968
rect 142516 29946 142540 29948
rect 142596 29946 142620 29948
rect 142676 29946 142700 29948
rect 142538 29894 142540 29946
rect 142602 29894 142614 29946
rect 142676 29894 142678 29946
rect 142516 29892 142540 29894
rect 142596 29892 142620 29894
rect 142676 29892 142700 29894
rect 142460 29872 142756 29892
rect 142460 28860 142756 28880
rect 142516 28858 142540 28860
rect 142596 28858 142620 28860
rect 142676 28858 142700 28860
rect 142538 28806 142540 28858
rect 142602 28806 142614 28858
rect 142676 28806 142678 28858
rect 142516 28804 142540 28806
rect 142596 28804 142620 28806
rect 142676 28804 142700 28806
rect 142460 28784 142756 28804
rect 142460 27772 142756 27792
rect 142516 27770 142540 27772
rect 142596 27770 142620 27772
rect 142676 27770 142700 27772
rect 142538 27718 142540 27770
rect 142602 27718 142614 27770
rect 142676 27718 142678 27770
rect 142516 27716 142540 27718
rect 142596 27716 142620 27718
rect 142676 27716 142700 27718
rect 142460 27696 142756 27716
rect 142460 26684 142756 26704
rect 142516 26682 142540 26684
rect 142596 26682 142620 26684
rect 142676 26682 142700 26684
rect 142538 26630 142540 26682
rect 142602 26630 142614 26682
rect 142676 26630 142678 26682
rect 142516 26628 142540 26630
rect 142596 26628 142620 26630
rect 142676 26628 142700 26630
rect 142460 26608 142756 26628
rect 142460 25596 142756 25616
rect 142516 25594 142540 25596
rect 142596 25594 142620 25596
rect 142676 25594 142700 25596
rect 142538 25542 142540 25594
rect 142602 25542 142614 25594
rect 142676 25542 142678 25594
rect 142516 25540 142540 25542
rect 142596 25540 142620 25542
rect 142676 25540 142700 25542
rect 142460 25520 142756 25540
rect 142460 24508 142756 24528
rect 142516 24506 142540 24508
rect 142596 24506 142620 24508
rect 142676 24506 142700 24508
rect 142538 24454 142540 24506
rect 142602 24454 142614 24506
rect 142676 24454 142678 24506
rect 142516 24452 142540 24454
rect 142596 24452 142620 24454
rect 142676 24452 142700 24454
rect 142460 24432 142756 24452
rect 142460 23420 142756 23440
rect 142516 23418 142540 23420
rect 142596 23418 142620 23420
rect 142676 23418 142700 23420
rect 142538 23366 142540 23418
rect 142602 23366 142614 23418
rect 142676 23366 142678 23418
rect 142516 23364 142540 23366
rect 142596 23364 142620 23366
rect 142676 23364 142700 23366
rect 142460 23344 142756 23364
rect 142460 22332 142756 22352
rect 142516 22330 142540 22332
rect 142596 22330 142620 22332
rect 142676 22330 142700 22332
rect 142538 22278 142540 22330
rect 142602 22278 142614 22330
rect 142676 22278 142678 22330
rect 142516 22276 142540 22278
rect 142596 22276 142620 22278
rect 142676 22276 142700 22278
rect 142460 22256 142756 22276
rect 142460 21244 142756 21264
rect 142516 21242 142540 21244
rect 142596 21242 142620 21244
rect 142676 21242 142700 21244
rect 142538 21190 142540 21242
rect 142602 21190 142614 21242
rect 142676 21190 142678 21242
rect 142516 21188 142540 21190
rect 142596 21188 142620 21190
rect 142676 21188 142700 21190
rect 142460 21168 142756 21188
rect 142460 20156 142756 20176
rect 142516 20154 142540 20156
rect 142596 20154 142620 20156
rect 142676 20154 142700 20156
rect 142538 20102 142540 20154
rect 142602 20102 142614 20154
rect 142676 20102 142678 20154
rect 142516 20100 142540 20102
rect 142596 20100 142620 20102
rect 142676 20100 142700 20102
rect 142460 20080 142756 20100
rect 140412 19168 140464 19174
rect 140412 19110 140464 19116
rect 81020 19068 81316 19088
rect 81076 19066 81100 19068
rect 81156 19066 81180 19068
rect 81236 19066 81260 19068
rect 81098 19014 81100 19066
rect 81162 19014 81174 19066
rect 81236 19014 81238 19066
rect 81076 19012 81100 19014
rect 81156 19012 81180 19014
rect 81236 19012 81260 19014
rect 81020 18992 81316 19012
rect 111740 19068 112036 19088
rect 111796 19066 111820 19068
rect 111876 19066 111900 19068
rect 111956 19066 111980 19068
rect 111818 19014 111820 19066
rect 111882 19014 111894 19066
rect 111956 19014 111958 19066
rect 111796 19012 111820 19014
rect 111876 19012 111900 19014
rect 111956 19012 111980 19014
rect 111740 18992 112036 19012
rect 142460 19068 142756 19088
rect 142516 19066 142540 19068
rect 142596 19066 142620 19068
rect 142676 19066 142700 19068
rect 142538 19014 142540 19066
rect 142602 19014 142614 19066
rect 142676 19014 142678 19066
rect 142516 19012 142540 19014
rect 142596 19012 142620 19014
rect 142676 19012 142700 19014
rect 142460 18992 142756 19012
rect 144564 18834 144592 117098
rect 146772 116346 146800 117098
rect 146760 116340 146812 116346
rect 146760 116282 146812 116288
rect 149532 20398 149560 117098
rect 150912 116346 150940 117098
rect 154132 116346 154160 117098
rect 154868 116346 154896 117098
rect 158812 116748 158864 116754
rect 158812 116690 158864 116696
rect 157820 116444 158116 116464
rect 157876 116442 157900 116444
rect 157956 116442 157980 116444
rect 158036 116442 158060 116444
rect 157898 116390 157900 116442
rect 157962 116390 157974 116442
rect 158036 116390 158038 116442
rect 157876 116388 157900 116390
rect 157956 116388 157980 116390
rect 158036 116388 158060 116390
rect 157820 116368 158116 116388
rect 150900 116340 150952 116346
rect 150900 116282 150952 116288
rect 154120 116340 154172 116346
rect 154120 116282 154172 116288
rect 154856 116340 154908 116346
rect 154856 116282 154908 116288
rect 158824 116142 158852 116690
rect 159100 116346 159128 117098
rect 162044 116890 162072 117098
rect 162124 117088 162176 117094
rect 162124 117030 162176 117036
rect 162032 116884 162084 116890
rect 162032 116826 162084 116832
rect 162136 116346 162164 117030
rect 164344 116346 164372 117098
rect 168208 116346 168236 117098
rect 159088 116340 159140 116346
rect 159088 116282 159140 116288
rect 162124 116340 162176 116346
rect 162124 116282 162176 116288
rect 164332 116340 164384 116346
rect 164332 116282 164384 116288
rect 168196 116340 168248 116346
rect 168196 116282 168248 116288
rect 171244 116142 171272 117098
rect 172900 116346 172928 117098
rect 173180 116988 173476 117008
rect 173236 116986 173260 116988
rect 173316 116986 173340 116988
rect 173396 116986 173420 116988
rect 173258 116934 173260 116986
rect 173322 116934 173334 116986
rect 173396 116934 173398 116986
rect 173236 116932 173260 116934
rect 173316 116932 173340 116934
rect 173396 116932 173420 116934
rect 173180 116912 173476 116932
rect 176028 116346 176056 117098
rect 176948 116346 176976 117098
rect 177580 117088 177632 117094
rect 177580 117030 177632 117036
rect 177592 116346 177620 117030
rect 172888 116340 172940 116346
rect 172888 116282 172940 116288
rect 176016 116340 176068 116346
rect 176016 116282 176068 116288
rect 176936 116340 176988 116346
rect 176936 116282 176988 116288
rect 177580 116340 177632 116346
rect 177580 116282 177632 116288
rect 158812 116136 158864 116142
rect 158812 116078 158864 116084
rect 171232 116136 171284 116142
rect 171232 116078 171284 116084
rect 173180 115900 173476 115920
rect 173236 115898 173260 115900
rect 173316 115898 173340 115900
rect 173396 115898 173420 115900
rect 173258 115846 173260 115898
rect 173322 115846 173334 115898
rect 173396 115846 173398 115898
rect 173236 115844 173260 115846
rect 173316 115844 173340 115846
rect 173396 115844 173420 115846
rect 173180 115824 173476 115844
rect 157820 115356 158116 115376
rect 157876 115354 157900 115356
rect 157956 115354 157980 115356
rect 158036 115354 158060 115356
rect 157898 115302 157900 115354
rect 157962 115302 157974 115354
rect 158036 115302 158038 115354
rect 157876 115300 157900 115302
rect 157956 115300 157980 115302
rect 158036 115300 158060 115302
rect 157820 115280 158116 115300
rect 173180 114812 173476 114832
rect 173236 114810 173260 114812
rect 173316 114810 173340 114812
rect 173396 114810 173420 114812
rect 173258 114758 173260 114810
rect 173322 114758 173334 114810
rect 173396 114758 173398 114810
rect 173236 114756 173260 114758
rect 173316 114756 173340 114758
rect 173396 114756 173420 114758
rect 173180 114736 173476 114756
rect 157820 114268 158116 114288
rect 157876 114266 157900 114268
rect 157956 114266 157980 114268
rect 158036 114266 158060 114268
rect 157898 114214 157900 114266
rect 157962 114214 157974 114266
rect 158036 114214 158038 114266
rect 157876 114212 157900 114214
rect 157956 114212 157980 114214
rect 158036 114212 158060 114214
rect 157820 114192 158116 114212
rect 173180 113724 173476 113744
rect 173236 113722 173260 113724
rect 173316 113722 173340 113724
rect 173396 113722 173420 113724
rect 173258 113670 173260 113722
rect 173322 113670 173334 113722
rect 173396 113670 173398 113722
rect 173236 113668 173260 113670
rect 173316 113668 173340 113670
rect 173396 113668 173420 113670
rect 173180 113648 173476 113668
rect 157820 113180 158116 113200
rect 157876 113178 157900 113180
rect 157956 113178 157980 113180
rect 158036 113178 158060 113180
rect 157898 113126 157900 113178
rect 157962 113126 157974 113178
rect 158036 113126 158038 113178
rect 157876 113124 157900 113126
rect 157956 113124 157980 113126
rect 158036 113124 158060 113126
rect 157820 113104 158116 113124
rect 173180 112636 173476 112656
rect 173236 112634 173260 112636
rect 173316 112634 173340 112636
rect 173396 112634 173420 112636
rect 173258 112582 173260 112634
rect 173322 112582 173334 112634
rect 173396 112582 173398 112634
rect 173236 112580 173260 112582
rect 173316 112580 173340 112582
rect 173396 112580 173420 112582
rect 173180 112560 173476 112580
rect 157820 112092 158116 112112
rect 157876 112090 157900 112092
rect 157956 112090 157980 112092
rect 158036 112090 158060 112092
rect 157898 112038 157900 112090
rect 157962 112038 157974 112090
rect 158036 112038 158038 112090
rect 157876 112036 157900 112038
rect 157956 112036 157980 112038
rect 158036 112036 158060 112038
rect 157820 112016 158116 112036
rect 173180 111548 173476 111568
rect 173236 111546 173260 111548
rect 173316 111546 173340 111548
rect 173396 111546 173420 111548
rect 173258 111494 173260 111546
rect 173322 111494 173334 111546
rect 173396 111494 173398 111546
rect 173236 111492 173260 111494
rect 173316 111492 173340 111494
rect 173396 111492 173420 111494
rect 173180 111472 173476 111492
rect 157820 111004 158116 111024
rect 157876 111002 157900 111004
rect 157956 111002 157980 111004
rect 158036 111002 158060 111004
rect 157898 110950 157900 111002
rect 157962 110950 157974 111002
rect 158036 110950 158038 111002
rect 157876 110948 157900 110950
rect 157956 110948 157980 110950
rect 158036 110948 158060 110950
rect 157820 110928 158116 110948
rect 173180 110460 173476 110480
rect 173236 110458 173260 110460
rect 173316 110458 173340 110460
rect 173396 110458 173420 110460
rect 173258 110406 173260 110458
rect 173322 110406 173334 110458
rect 173396 110406 173398 110458
rect 173236 110404 173260 110406
rect 173316 110404 173340 110406
rect 173396 110404 173420 110406
rect 173180 110384 173476 110404
rect 157820 109916 158116 109936
rect 157876 109914 157900 109916
rect 157956 109914 157980 109916
rect 158036 109914 158060 109916
rect 157898 109862 157900 109914
rect 157962 109862 157974 109914
rect 158036 109862 158038 109914
rect 157876 109860 157900 109862
rect 157956 109860 157980 109862
rect 158036 109860 158060 109862
rect 157820 109840 158116 109860
rect 173180 109372 173476 109392
rect 173236 109370 173260 109372
rect 173316 109370 173340 109372
rect 173396 109370 173420 109372
rect 173258 109318 173260 109370
rect 173322 109318 173334 109370
rect 173396 109318 173398 109370
rect 173236 109316 173260 109318
rect 173316 109316 173340 109318
rect 173396 109316 173420 109318
rect 173180 109296 173476 109316
rect 157820 108828 158116 108848
rect 157876 108826 157900 108828
rect 157956 108826 157980 108828
rect 158036 108826 158060 108828
rect 157898 108774 157900 108826
rect 157962 108774 157974 108826
rect 158036 108774 158038 108826
rect 157876 108772 157900 108774
rect 157956 108772 157980 108774
rect 158036 108772 158060 108774
rect 157820 108752 158116 108772
rect 173180 108284 173476 108304
rect 173236 108282 173260 108284
rect 173316 108282 173340 108284
rect 173396 108282 173420 108284
rect 173258 108230 173260 108282
rect 173322 108230 173334 108282
rect 173396 108230 173398 108282
rect 173236 108228 173260 108230
rect 173316 108228 173340 108230
rect 173396 108228 173420 108230
rect 173180 108208 173476 108228
rect 157820 107740 158116 107760
rect 157876 107738 157900 107740
rect 157956 107738 157980 107740
rect 158036 107738 158060 107740
rect 157898 107686 157900 107738
rect 157962 107686 157974 107738
rect 158036 107686 158038 107738
rect 157876 107684 157900 107686
rect 157956 107684 157980 107686
rect 158036 107684 158060 107686
rect 157820 107664 158116 107684
rect 173180 107196 173476 107216
rect 173236 107194 173260 107196
rect 173316 107194 173340 107196
rect 173396 107194 173420 107196
rect 173258 107142 173260 107194
rect 173322 107142 173334 107194
rect 173396 107142 173398 107194
rect 173236 107140 173260 107142
rect 173316 107140 173340 107142
rect 173396 107140 173420 107142
rect 173180 107120 173476 107140
rect 157820 106652 158116 106672
rect 157876 106650 157900 106652
rect 157956 106650 157980 106652
rect 158036 106650 158060 106652
rect 157898 106598 157900 106650
rect 157962 106598 157974 106650
rect 158036 106598 158038 106650
rect 157876 106596 157900 106598
rect 157956 106596 157980 106598
rect 158036 106596 158060 106598
rect 157820 106576 158116 106596
rect 173180 106108 173476 106128
rect 173236 106106 173260 106108
rect 173316 106106 173340 106108
rect 173396 106106 173420 106108
rect 173258 106054 173260 106106
rect 173322 106054 173334 106106
rect 173396 106054 173398 106106
rect 173236 106052 173260 106054
rect 173316 106052 173340 106054
rect 173396 106052 173420 106054
rect 173180 106032 173476 106052
rect 157820 105564 158116 105584
rect 157876 105562 157900 105564
rect 157956 105562 157980 105564
rect 158036 105562 158060 105564
rect 157898 105510 157900 105562
rect 157962 105510 157974 105562
rect 158036 105510 158038 105562
rect 157876 105508 157900 105510
rect 157956 105508 157980 105510
rect 158036 105508 158060 105510
rect 157820 105488 158116 105508
rect 173180 105020 173476 105040
rect 173236 105018 173260 105020
rect 173316 105018 173340 105020
rect 173396 105018 173420 105020
rect 173258 104966 173260 105018
rect 173322 104966 173334 105018
rect 173396 104966 173398 105018
rect 173236 104964 173260 104966
rect 173316 104964 173340 104966
rect 173396 104964 173420 104966
rect 173180 104944 173476 104964
rect 157820 104476 158116 104496
rect 157876 104474 157900 104476
rect 157956 104474 157980 104476
rect 158036 104474 158060 104476
rect 157898 104422 157900 104474
rect 157962 104422 157974 104474
rect 158036 104422 158038 104474
rect 157876 104420 157900 104422
rect 157956 104420 157980 104422
rect 158036 104420 158060 104422
rect 157820 104400 158116 104420
rect 173180 103932 173476 103952
rect 173236 103930 173260 103932
rect 173316 103930 173340 103932
rect 173396 103930 173420 103932
rect 173258 103878 173260 103930
rect 173322 103878 173334 103930
rect 173396 103878 173398 103930
rect 173236 103876 173260 103878
rect 173316 103876 173340 103878
rect 173396 103876 173420 103878
rect 173180 103856 173476 103876
rect 157820 103388 158116 103408
rect 157876 103386 157900 103388
rect 157956 103386 157980 103388
rect 158036 103386 158060 103388
rect 157898 103334 157900 103386
rect 157962 103334 157974 103386
rect 158036 103334 158038 103386
rect 157876 103332 157900 103334
rect 157956 103332 157980 103334
rect 158036 103332 158060 103334
rect 157820 103312 158116 103332
rect 173180 102844 173476 102864
rect 173236 102842 173260 102844
rect 173316 102842 173340 102844
rect 173396 102842 173420 102844
rect 173258 102790 173260 102842
rect 173322 102790 173334 102842
rect 173396 102790 173398 102842
rect 173236 102788 173260 102790
rect 173316 102788 173340 102790
rect 173396 102788 173420 102790
rect 173180 102768 173476 102788
rect 157820 102300 158116 102320
rect 157876 102298 157900 102300
rect 157956 102298 157980 102300
rect 158036 102298 158060 102300
rect 157898 102246 157900 102298
rect 157962 102246 157974 102298
rect 158036 102246 158038 102298
rect 157876 102244 157900 102246
rect 157956 102244 157980 102246
rect 158036 102244 158060 102246
rect 157820 102224 158116 102244
rect 173180 101756 173476 101776
rect 173236 101754 173260 101756
rect 173316 101754 173340 101756
rect 173396 101754 173420 101756
rect 173258 101702 173260 101754
rect 173322 101702 173334 101754
rect 173396 101702 173398 101754
rect 173236 101700 173260 101702
rect 173316 101700 173340 101702
rect 173396 101700 173420 101702
rect 173180 101680 173476 101700
rect 157820 101212 158116 101232
rect 157876 101210 157900 101212
rect 157956 101210 157980 101212
rect 158036 101210 158060 101212
rect 157898 101158 157900 101210
rect 157962 101158 157974 101210
rect 158036 101158 158038 101210
rect 157876 101156 157900 101158
rect 157956 101156 157980 101158
rect 158036 101156 158060 101158
rect 157820 101136 158116 101156
rect 173180 100668 173476 100688
rect 173236 100666 173260 100668
rect 173316 100666 173340 100668
rect 173396 100666 173420 100668
rect 173258 100614 173260 100666
rect 173322 100614 173334 100666
rect 173396 100614 173398 100666
rect 173236 100612 173260 100614
rect 173316 100612 173340 100614
rect 173396 100612 173420 100614
rect 173180 100592 173476 100612
rect 157820 100124 158116 100144
rect 157876 100122 157900 100124
rect 157956 100122 157980 100124
rect 158036 100122 158060 100124
rect 157898 100070 157900 100122
rect 157962 100070 157974 100122
rect 158036 100070 158038 100122
rect 157876 100068 157900 100070
rect 157956 100068 157980 100070
rect 158036 100068 158060 100070
rect 157820 100048 158116 100068
rect 173180 99580 173476 99600
rect 173236 99578 173260 99580
rect 173316 99578 173340 99580
rect 173396 99578 173420 99580
rect 173258 99526 173260 99578
rect 173322 99526 173334 99578
rect 173396 99526 173398 99578
rect 173236 99524 173260 99526
rect 173316 99524 173340 99526
rect 173396 99524 173420 99526
rect 173180 99504 173476 99524
rect 157820 99036 158116 99056
rect 157876 99034 157900 99036
rect 157956 99034 157980 99036
rect 158036 99034 158060 99036
rect 157898 98982 157900 99034
rect 157962 98982 157974 99034
rect 158036 98982 158038 99034
rect 157876 98980 157900 98982
rect 157956 98980 157980 98982
rect 158036 98980 158060 98982
rect 157820 98960 158116 98980
rect 173180 98492 173476 98512
rect 173236 98490 173260 98492
rect 173316 98490 173340 98492
rect 173396 98490 173420 98492
rect 173258 98438 173260 98490
rect 173322 98438 173334 98490
rect 173396 98438 173398 98490
rect 173236 98436 173260 98438
rect 173316 98436 173340 98438
rect 173396 98436 173420 98438
rect 173180 98416 173476 98436
rect 157820 97948 158116 97968
rect 157876 97946 157900 97948
rect 157956 97946 157980 97948
rect 158036 97946 158060 97948
rect 157898 97894 157900 97946
rect 157962 97894 157974 97946
rect 158036 97894 158038 97946
rect 157876 97892 157900 97894
rect 157956 97892 157980 97894
rect 158036 97892 158060 97894
rect 157820 97872 158116 97892
rect 173180 97404 173476 97424
rect 173236 97402 173260 97404
rect 173316 97402 173340 97404
rect 173396 97402 173420 97404
rect 173258 97350 173260 97402
rect 173322 97350 173334 97402
rect 173396 97350 173398 97402
rect 173236 97348 173260 97350
rect 173316 97348 173340 97350
rect 173396 97348 173420 97350
rect 173180 97328 173476 97348
rect 157820 96860 158116 96880
rect 157876 96858 157900 96860
rect 157956 96858 157980 96860
rect 158036 96858 158060 96860
rect 157898 96806 157900 96858
rect 157962 96806 157974 96858
rect 158036 96806 158038 96858
rect 157876 96804 157900 96806
rect 157956 96804 157980 96806
rect 158036 96804 158060 96806
rect 157820 96784 158116 96804
rect 173180 96316 173476 96336
rect 173236 96314 173260 96316
rect 173316 96314 173340 96316
rect 173396 96314 173420 96316
rect 173258 96262 173260 96314
rect 173322 96262 173334 96314
rect 173396 96262 173398 96314
rect 173236 96260 173260 96262
rect 173316 96260 173340 96262
rect 173396 96260 173420 96262
rect 173180 96240 173476 96260
rect 157820 95772 158116 95792
rect 157876 95770 157900 95772
rect 157956 95770 157980 95772
rect 158036 95770 158060 95772
rect 157898 95718 157900 95770
rect 157962 95718 157974 95770
rect 158036 95718 158038 95770
rect 157876 95716 157900 95718
rect 157956 95716 157980 95718
rect 158036 95716 158060 95718
rect 157820 95696 158116 95716
rect 173180 95228 173476 95248
rect 173236 95226 173260 95228
rect 173316 95226 173340 95228
rect 173396 95226 173420 95228
rect 173258 95174 173260 95226
rect 173322 95174 173334 95226
rect 173396 95174 173398 95226
rect 173236 95172 173260 95174
rect 173316 95172 173340 95174
rect 173396 95172 173420 95174
rect 173180 95152 173476 95172
rect 157820 94684 158116 94704
rect 157876 94682 157900 94684
rect 157956 94682 157980 94684
rect 158036 94682 158060 94684
rect 157898 94630 157900 94682
rect 157962 94630 157974 94682
rect 158036 94630 158038 94682
rect 157876 94628 157900 94630
rect 157956 94628 157980 94630
rect 158036 94628 158060 94630
rect 157820 94608 158116 94628
rect 173180 94140 173476 94160
rect 173236 94138 173260 94140
rect 173316 94138 173340 94140
rect 173396 94138 173420 94140
rect 173258 94086 173260 94138
rect 173322 94086 173334 94138
rect 173396 94086 173398 94138
rect 173236 94084 173260 94086
rect 173316 94084 173340 94086
rect 173396 94084 173420 94086
rect 173180 94064 173476 94084
rect 157820 93596 158116 93616
rect 157876 93594 157900 93596
rect 157956 93594 157980 93596
rect 158036 93594 158060 93596
rect 157898 93542 157900 93594
rect 157962 93542 157974 93594
rect 158036 93542 158038 93594
rect 157876 93540 157900 93542
rect 157956 93540 157980 93542
rect 158036 93540 158060 93542
rect 157820 93520 158116 93540
rect 173180 93052 173476 93072
rect 173236 93050 173260 93052
rect 173316 93050 173340 93052
rect 173396 93050 173420 93052
rect 173258 92998 173260 93050
rect 173322 92998 173334 93050
rect 173396 92998 173398 93050
rect 173236 92996 173260 92998
rect 173316 92996 173340 92998
rect 173396 92996 173420 92998
rect 173180 92976 173476 92996
rect 157820 92508 158116 92528
rect 157876 92506 157900 92508
rect 157956 92506 157980 92508
rect 158036 92506 158060 92508
rect 157898 92454 157900 92506
rect 157962 92454 157974 92506
rect 158036 92454 158038 92506
rect 157876 92452 157900 92454
rect 157956 92452 157980 92454
rect 158036 92452 158060 92454
rect 157820 92432 158116 92452
rect 173180 91964 173476 91984
rect 173236 91962 173260 91964
rect 173316 91962 173340 91964
rect 173396 91962 173420 91964
rect 173258 91910 173260 91962
rect 173322 91910 173334 91962
rect 173396 91910 173398 91962
rect 173236 91908 173260 91910
rect 173316 91908 173340 91910
rect 173396 91908 173420 91910
rect 173180 91888 173476 91908
rect 157820 91420 158116 91440
rect 157876 91418 157900 91420
rect 157956 91418 157980 91420
rect 158036 91418 158060 91420
rect 157898 91366 157900 91418
rect 157962 91366 157974 91418
rect 158036 91366 158038 91418
rect 157876 91364 157900 91366
rect 157956 91364 157980 91366
rect 158036 91364 158060 91366
rect 157820 91344 158116 91364
rect 173180 90876 173476 90896
rect 173236 90874 173260 90876
rect 173316 90874 173340 90876
rect 173396 90874 173420 90876
rect 173258 90822 173260 90874
rect 173322 90822 173334 90874
rect 173396 90822 173398 90874
rect 173236 90820 173260 90822
rect 173316 90820 173340 90822
rect 173396 90820 173420 90822
rect 173180 90800 173476 90820
rect 157820 90332 158116 90352
rect 157876 90330 157900 90332
rect 157956 90330 157980 90332
rect 158036 90330 158060 90332
rect 157898 90278 157900 90330
rect 157962 90278 157974 90330
rect 158036 90278 158038 90330
rect 157876 90276 157900 90278
rect 157956 90276 157980 90278
rect 158036 90276 158060 90278
rect 157820 90256 158116 90276
rect 173180 89788 173476 89808
rect 173236 89786 173260 89788
rect 173316 89786 173340 89788
rect 173396 89786 173420 89788
rect 173258 89734 173260 89786
rect 173322 89734 173334 89786
rect 173396 89734 173398 89786
rect 173236 89732 173260 89734
rect 173316 89732 173340 89734
rect 173396 89732 173420 89734
rect 173180 89712 173476 89732
rect 157820 89244 158116 89264
rect 157876 89242 157900 89244
rect 157956 89242 157980 89244
rect 158036 89242 158060 89244
rect 157898 89190 157900 89242
rect 157962 89190 157974 89242
rect 158036 89190 158038 89242
rect 157876 89188 157900 89190
rect 157956 89188 157980 89190
rect 158036 89188 158060 89190
rect 157820 89168 158116 89188
rect 173180 88700 173476 88720
rect 173236 88698 173260 88700
rect 173316 88698 173340 88700
rect 173396 88698 173420 88700
rect 173258 88646 173260 88698
rect 173322 88646 173334 88698
rect 173396 88646 173398 88698
rect 173236 88644 173260 88646
rect 173316 88644 173340 88646
rect 173396 88644 173420 88646
rect 173180 88624 173476 88644
rect 157820 88156 158116 88176
rect 157876 88154 157900 88156
rect 157956 88154 157980 88156
rect 158036 88154 158060 88156
rect 157898 88102 157900 88154
rect 157962 88102 157974 88154
rect 158036 88102 158038 88154
rect 157876 88100 157900 88102
rect 157956 88100 157980 88102
rect 158036 88100 158060 88102
rect 157820 88080 158116 88100
rect 173180 87612 173476 87632
rect 173236 87610 173260 87612
rect 173316 87610 173340 87612
rect 173396 87610 173420 87612
rect 173258 87558 173260 87610
rect 173322 87558 173334 87610
rect 173396 87558 173398 87610
rect 173236 87556 173260 87558
rect 173316 87556 173340 87558
rect 173396 87556 173420 87558
rect 173180 87536 173476 87556
rect 157820 87068 158116 87088
rect 157876 87066 157900 87068
rect 157956 87066 157980 87068
rect 158036 87066 158060 87068
rect 157898 87014 157900 87066
rect 157962 87014 157974 87066
rect 158036 87014 158038 87066
rect 157876 87012 157900 87014
rect 157956 87012 157980 87014
rect 158036 87012 158060 87014
rect 157820 86992 158116 87012
rect 173180 86524 173476 86544
rect 173236 86522 173260 86524
rect 173316 86522 173340 86524
rect 173396 86522 173420 86524
rect 173258 86470 173260 86522
rect 173322 86470 173334 86522
rect 173396 86470 173398 86522
rect 173236 86468 173260 86470
rect 173316 86468 173340 86470
rect 173396 86468 173420 86470
rect 173180 86448 173476 86468
rect 157820 85980 158116 86000
rect 157876 85978 157900 85980
rect 157956 85978 157980 85980
rect 158036 85978 158060 85980
rect 157898 85926 157900 85978
rect 157962 85926 157974 85978
rect 158036 85926 158038 85978
rect 157876 85924 157900 85926
rect 157956 85924 157980 85926
rect 158036 85924 158060 85926
rect 157820 85904 158116 85924
rect 173180 85436 173476 85456
rect 173236 85434 173260 85436
rect 173316 85434 173340 85436
rect 173396 85434 173420 85436
rect 173258 85382 173260 85434
rect 173322 85382 173334 85434
rect 173396 85382 173398 85434
rect 173236 85380 173260 85382
rect 173316 85380 173340 85382
rect 173396 85380 173420 85382
rect 173180 85360 173476 85380
rect 157820 84892 158116 84912
rect 157876 84890 157900 84892
rect 157956 84890 157980 84892
rect 158036 84890 158060 84892
rect 157898 84838 157900 84890
rect 157962 84838 157974 84890
rect 158036 84838 158038 84890
rect 157876 84836 157900 84838
rect 157956 84836 157980 84838
rect 158036 84836 158060 84838
rect 157820 84816 158116 84836
rect 173180 84348 173476 84368
rect 173236 84346 173260 84348
rect 173316 84346 173340 84348
rect 173396 84346 173420 84348
rect 173258 84294 173260 84346
rect 173322 84294 173334 84346
rect 173396 84294 173398 84346
rect 173236 84292 173260 84294
rect 173316 84292 173340 84294
rect 173396 84292 173420 84294
rect 173180 84272 173476 84292
rect 157820 83804 158116 83824
rect 157876 83802 157900 83804
rect 157956 83802 157980 83804
rect 158036 83802 158060 83804
rect 157898 83750 157900 83802
rect 157962 83750 157974 83802
rect 158036 83750 158038 83802
rect 157876 83748 157900 83750
rect 157956 83748 157980 83750
rect 158036 83748 158060 83750
rect 157820 83728 158116 83748
rect 173180 83260 173476 83280
rect 173236 83258 173260 83260
rect 173316 83258 173340 83260
rect 173396 83258 173420 83260
rect 173258 83206 173260 83258
rect 173322 83206 173334 83258
rect 173396 83206 173398 83258
rect 173236 83204 173260 83206
rect 173316 83204 173340 83206
rect 173396 83204 173420 83206
rect 173180 83184 173476 83204
rect 157820 82716 158116 82736
rect 157876 82714 157900 82716
rect 157956 82714 157980 82716
rect 158036 82714 158060 82716
rect 157898 82662 157900 82714
rect 157962 82662 157974 82714
rect 158036 82662 158038 82714
rect 157876 82660 157900 82662
rect 157956 82660 157980 82662
rect 158036 82660 158060 82662
rect 157820 82640 158116 82660
rect 173180 82172 173476 82192
rect 173236 82170 173260 82172
rect 173316 82170 173340 82172
rect 173396 82170 173420 82172
rect 173258 82118 173260 82170
rect 173322 82118 173334 82170
rect 173396 82118 173398 82170
rect 173236 82116 173260 82118
rect 173316 82116 173340 82118
rect 173396 82116 173420 82118
rect 173180 82096 173476 82116
rect 157820 81628 158116 81648
rect 157876 81626 157900 81628
rect 157956 81626 157980 81628
rect 158036 81626 158060 81628
rect 157898 81574 157900 81626
rect 157962 81574 157974 81626
rect 158036 81574 158038 81626
rect 157876 81572 157900 81574
rect 157956 81572 157980 81574
rect 158036 81572 158060 81574
rect 157820 81552 158116 81572
rect 173180 81084 173476 81104
rect 173236 81082 173260 81084
rect 173316 81082 173340 81084
rect 173396 81082 173420 81084
rect 173258 81030 173260 81082
rect 173322 81030 173334 81082
rect 173396 81030 173398 81082
rect 173236 81028 173260 81030
rect 173316 81028 173340 81030
rect 173396 81028 173420 81030
rect 173180 81008 173476 81028
rect 157820 80540 158116 80560
rect 157876 80538 157900 80540
rect 157956 80538 157980 80540
rect 158036 80538 158060 80540
rect 157898 80486 157900 80538
rect 157962 80486 157974 80538
rect 158036 80486 158038 80538
rect 157876 80484 157900 80486
rect 157956 80484 157980 80486
rect 158036 80484 158060 80486
rect 157820 80464 158116 80484
rect 173180 79996 173476 80016
rect 173236 79994 173260 79996
rect 173316 79994 173340 79996
rect 173396 79994 173420 79996
rect 173258 79942 173260 79994
rect 173322 79942 173334 79994
rect 173396 79942 173398 79994
rect 173236 79940 173260 79942
rect 173316 79940 173340 79942
rect 173396 79940 173420 79942
rect 173180 79920 173476 79940
rect 157820 79452 158116 79472
rect 157876 79450 157900 79452
rect 157956 79450 157980 79452
rect 158036 79450 158060 79452
rect 157898 79398 157900 79450
rect 157962 79398 157974 79450
rect 158036 79398 158038 79450
rect 157876 79396 157900 79398
rect 157956 79396 157980 79398
rect 158036 79396 158060 79398
rect 157820 79376 158116 79396
rect 173180 78908 173476 78928
rect 173236 78906 173260 78908
rect 173316 78906 173340 78908
rect 173396 78906 173420 78908
rect 173258 78854 173260 78906
rect 173322 78854 173334 78906
rect 173396 78854 173398 78906
rect 173236 78852 173260 78854
rect 173316 78852 173340 78854
rect 173396 78852 173420 78854
rect 173180 78832 173476 78852
rect 157820 78364 158116 78384
rect 157876 78362 157900 78364
rect 157956 78362 157980 78364
rect 158036 78362 158060 78364
rect 157898 78310 157900 78362
rect 157962 78310 157974 78362
rect 158036 78310 158038 78362
rect 157876 78308 157900 78310
rect 157956 78308 157980 78310
rect 158036 78308 158060 78310
rect 157820 78288 158116 78308
rect 173180 77820 173476 77840
rect 173236 77818 173260 77820
rect 173316 77818 173340 77820
rect 173396 77818 173420 77820
rect 173258 77766 173260 77818
rect 173322 77766 173334 77818
rect 173396 77766 173398 77818
rect 173236 77764 173260 77766
rect 173316 77764 173340 77766
rect 173396 77764 173420 77766
rect 173180 77744 173476 77764
rect 157820 77276 158116 77296
rect 157876 77274 157900 77276
rect 157956 77274 157980 77276
rect 158036 77274 158060 77276
rect 157898 77222 157900 77274
rect 157962 77222 157974 77274
rect 158036 77222 158038 77274
rect 157876 77220 157900 77222
rect 157956 77220 157980 77222
rect 158036 77220 158060 77222
rect 157820 77200 158116 77220
rect 173180 76732 173476 76752
rect 173236 76730 173260 76732
rect 173316 76730 173340 76732
rect 173396 76730 173420 76732
rect 173258 76678 173260 76730
rect 173322 76678 173334 76730
rect 173396 76678 173398 76730
rect 173236 76676 173260 76678
rect 173316 76676 173340 76678
rect 173396 76676 173420 76678
rect 173180 76656 173476 76676
rect 157820 76188 158116 76208
rect 157876 76186 157900 76188
rect 157956 76186 157980 76188
rect 158036 76186 158060 76188
rect 157898 76134 157900 76186
rect 157962 76134 157974 76186
rect 158036 76134 158038 76186
rect 157876 76132 157900 76134
rect 157956 76132 157980 76134
rect 158036 76132 158060 76134
rect 157820 76112 158116 76132
rect 173180 75644 173476 75664
rect 173236 75642 173260 75644
rect 173316 75642 173340 75644
rect 173396 75642 173420 75644
rect 173258 75590 173260 75642
rect 173322 75590 173334 75642
rect 173396 75590 173398 75642
rect 173236 75588 173260 75590
rect 173316 75588 173340 75590
rect 173396 75588 173420 75590
rect 173180 75568 173476 75588
rect 157820 75100 158116 75120
rect 157876 75098 157900 75100
rect 157956 75098 157980 75100
rect 158036 75098 158060 75100
rect 157898 75046 157900 75098
rect 157962 75046 157974 75098
rect 158036 75046 158038 75098
rect 157876 75044 157900 75046
rect 157956 75044 157980 75046
rect 158036 75044 158060 75046
rect 157820 75024 158116 75044
rect 173180 74556 173476 74576
rect 173236 74554 173260 74556
rect 173316 74554 173340 74556
rect 173396 74554 173420 74556
rect 173258 74502 173260 74554
rect 173322 74502 173334 74554
rect 173396 74502 173398 74554
rect 173236 74500 173260 74502
rect 173316 74500 173340 74502
rect 173396 74500 173420 74502
rect 173180 74480 173476 74500
rect 157820 74012 158116 74032
rect 157876 74010 157900 74012
rect 157956 74010 157980 74012
rect 158036 74010 158060 74012
rect 157898 73958 157900 74010
rect 157962 73958 157974 74010
rect 158036 73958 158038 74010
rect 157876 73956 157900 73958
rect 157956 73956 157980 73958
rect 158036 73956 158060 73958
rect 157820 73936 158116 73956
rect 173180 73468 173476 73488
rect 173236 73466 173260 73468
rect 173316 73466 173340 73468
rect 173396 73466 173420 73468
rect 173258 73414 173260 73466
rect 173322 73414 173334 73466
rect 173396 73414 173398 73466
rect 173236 73412 173260 73414
rect 173316 73412 173340 73414
rect 173396 73412 173420 73414
rect 173180 73392 173476 73412
rect 157820 72924 158116 72944
rect 157876 72922 157900 72924
rect 157956 72922 157980 72924
rect 158036 72922 158060 72924
rect 157898 72870 157900 72922
rect 157962 72870 157974 72922
rect 158036 72870 158038 72922
rect 157876 72868 157900 72870
rect 157956 72868 157980 72870
rect 158036 72868 158060 72870
rect 157820 72848 158116 72868
rect 173180 72380 173476 72400
rect 173236 72378 173260 72380
rect 173316 72378 173340 72380
rect 173396 72378 173420 72380
rect 173258 72326 173260 72378
rect 173322 72326 173334 72378
rect 173396 72326 173398 72378
rect 173236 72324 173260 72326
rect 173316 72324 173340 72326
rect 173396 72324 173420 72326
rect 173180 72304 173476 72324
rect 157820 71836 158116 71856
rect 157876 71834 157900 71836
rect 157956 71834 157980 71836
rect 158036 71834 158060 71836
rect 157898 71782 157900 71834
rect 157962 71782 157974 71834
rect 158036 71782 158038 71834
rect 157876 71780 157900 71782
rect 157956 71780 157980 71782
rect 158036 71780 158060 71782
rect 157820 71760 158116 71780
rect 173180 71292 173476 71312
rect 173236 71290 173260 71292
rect 173316 71290 173340 71292
rect 173396 71290 173420 71292
rect 173258 71238 173260 71290
rect 173322 71238 173334 71290
rect 173396 71238 173398 71290
rect 173236 71236 173260 71238
rect 173316 71236 173340 71238
rect 173396 71236 173420 71238
rect 173180 71216 173476 71236
rect 157820 70748 158116 70768
rect 157876 70746 157900 70748
rect 157956 70746 157980 70748
rect 158036 70746 158060 70748
rect 157898 70694 157900 70746
rect 157962 70694 157974 70746
rect 158036 70694 158038 70746
rect 157876 70692 157900 70694
rect 157956 70692 157980 70694
rect 158036 70692 158060 70694
rect 157820 70672 158116 70692
rect 173180 70204 173476 70224
rect 173236 70202 173260 70204
rect 173316 70202 173340 70204
rect 173396 70202 173420 70204
rect 173258 70150 173260 70202
rect 173322 70150 173334 70202
rect 173396 70150 173398 70202
rect 173236 70148 173260 70150
rect 173316 70148 173340 70150
rect 173396 70148 173420 70150
rect 173180 70128 173476 70148
rect 157820 69660 158116 69680
rect 157876 69658 157900 69660
rect 157956 69658 157980 69660
rect 158036 69658 158060 69660
rect 157898 69606 157900 69658
rect 157962 69606 157974 69658
rect 158036 69606 158038 69658
rect 157876 69604 157900 69606
rect 157956 69604 157980 69606
rect 158036 69604 158060 69606
rect 157820 69584 158116 69604
rect 173180 69116 173476 69136
rect 173236 69114 173260 69116
rect 173316 69114 173340 69116
rect 173396 69114 173420 69116
rect 173258 69062 173260 69114
rect 173322 69062 173334 69114
rect 173396 69062 173398 69114
rect 173236 69060 173260 69062
rect 173316 69060 173340 69062
rect 173396 69060 173420 69062
rect 173180 69040 173476 69060
rect 157820 68572 158116 68592
rect 157876 68570 157900 68572
rect 157956 68570 157980 68572
rect 158036 68570 158060 68572
rect 157898 68518 157900 68570
rect 157962 68518 157974 68570
rect 158036 68518 158038 68570
rect 157876 68516 157900 68518
rect 157956 68516 157980 68518
rect 158036 68516 158060 68518
rect 157820 68496 158116 68516
rect 173180 68028 173476 68048
rect 173236 68026 173260 68028
rect 173316 68026 173340 68028
rect 173396 68026 173420 68028
rect 173258 67974 173260 68026
rect 173322 67974 173334 68026
rect 173396 67974 173398 68026
rect 173236 67972 173260 67974
rect 173316 67972 173340 67974
rect 173396 67972 173420 67974
rect 173180 67952 173476 67972
rect 157820 67484 158116 67504
rect 157876 67482 157900 67484
rect 157956 67482 157980 67484
rect 158036 67482 158060 67484
rect 157898 67430 157900 67482
rect 157962 67430 157974 67482
rect 158036 67430 158038 67482
rect 157876 67428 157900 67430
rect 157956 67428 157980 67430
rect 158036 67428 158060 67430
rect 157820 67408 158116 67428
rect 173180 66940 173476 66960
rect 173236 66938 173260 66940
rect 173316 66938 173340 66940
rect 173396 66938 173420 66940
rect 173258 66886 173260 66938
rect 173322 66886 173334 66938
rect 173396 66886 173398 66938
rect 173236 66884 173260 66886
rect 173316 66884 173340 66886
rect 173396 66884 173420 66886
rect 173180 66864 173476 66884
rect 157820 66396 158116 66416
rect 157876 66394 157900 66396
rect 157956 66394 157980 66396
rect 158036 66394 158060 66396
rect 157898 66342 157900 66394
rect 157962 66342 157974 66394
rect 158036 66342 158038 66394
rect 157876 66340 157900 66342
rect 157956 66340 157980 66342
rect 158036 66340 158060 66342
rect 157820 66320 158116 66340
rect 173180 65852 173476 65872
rect 173236 65850 173260 65852
rect 173316 65850 173340 65852
rect 173396 65850 173420 65852
rect 173258 65798 173260 65850
rect 173322 65798 173334 65850
rect 173396 65798 173398 65850
rect 173236 65796 173260 65798
rect 173316 65796 173340 65798
rect 173396 65796 173420 65798
rect 173180 65776 173476 65796
rect 157820 65308 158116 65328
rect 157876 65306 157900 65308
rect 157956 65306 157980 65308
rect 158036 65306 158060 65308
rect 157898 65254 157900 65306
rect 157962 65254 157974 65306
rect 158036 65254 158038 65306
rect 157876 65252 157900 65254
rect 157956 65252 157980 65254
rect 158036 65252 158060 65254
rect 157820 65232 158116 65252
rect 173180 64764 173476 64784
rect 173236 64762 173260 64764
rect 173316 64762 173340 64764
rect 173396 64762 173420 64764
rect 173258 64710 173260 64762
rect 173322 64710 173334 64762
rect 173396 64710 173398 64762
rect 173236 64708 173260 64710
rect 173316 64708 173340 64710
rect 173396 64708 173420 64710
rect 173180 64688 173476 64708
rect 157820 64220 158116 64240
rect 157876 64218 157900 64220
rect 157956 64218 157980 64220
rect 158036 64218 158060 64220
rect 157898 64166 157900 64218
rect 157962 64166 157974 64218
rect 158036 64166 158038 64218
rect 157876 64164 157900 64166
rect 157956 64164 157980 64166
rect 158036 64164 158060 64166
rect 157820 64144 158116 64164
rect 173180 63676 173476 63696
rect 173236 63674 173260 63676
rect 173316 63674 173340 63676
rect 173396 63674 173420 63676
rect 173258 63622 173260 63674
rect 173322 63622 173334 63674
rect 173396 63622 173398 63674
rect 173236 63620 173260 63622
rect 173316 63620 173340 63622
rect 173396 63620 173420 63622
rect 173180 63600 173476 63620
rect 157820 63132 158116 63152
rect 157876 63130 157900 63132
rect 157956 63130 157980 63132
rect 158036 63130 158060 63132
rect 157898 63078 157900 63130
rect 157962 63078 157974 63130
rect 158036 63078 158038 63130
rect 157876 63076 157900 63078
rect 157956 63076 157980 63078
rect 158036 63076 158060 63078
rect 157820 63056 158116 63076
rect 173180 62588 173476 62608
rect 173236 62586 173260 62588
rect 173316 62586 173340 62588
rect 173396 62586 173420 62588
rect 173258 62534 173260 62586
rect 173322 62534 173334 62586
rect 173396 62534 173398 62586
rect 173236 62532 173260 62534
rect 173316 62532 173340 62534
rect 173396 62532 173420 62534
rect 173180 62512 173476 62532
rect 157820 62044 158116 62064
rect 157876 62042 157900 62044
rect 157956 62042 157980 62044
rect 158036 62042 158060 62044
rect 157898 61990 157900 62042
rect 157962 61990 157974 62042
rect 158036 61990 158038 62042
rect 157876 61988 157900 61990
rect 157956 61988 157980 61990
rect 158036 61988 158060 61990
rect 157820 61968 158116 61988
rect 173180 61500 173476 61520
rect 173236 61498 173260 61500
rect 173316 61498 173340 61500
rect 173396 61498 173420 61500
rect 173258 61446 173260 61498
rect 173322 61446 173334 61498
rect 173396 61446 173398 61498
rect 173236 61444 173260 61446
rect 173316 61444 173340 61446
rect 173396 61444 173420 61446
rect 173180 61424 173476 61444
rect 157820 60956 158116 60976
rect 157876 60954 157900 60956
rect 157956 60954 157980 60956
rect 158036 60954 158060 60956
rect 157898 60902 157900 60954
rect 157962 60902 157974 60954
rect 158036 60902 158038 60954
rect 157876 60900 157900 60902
rect 157956 60900 157980 60902
rect 158036 60900 158060 60902
rect 157820 60880 158116 60900
rect 173180 60412 173476 60432
rect 173236 60410 173260 60412
rect 173316 60410 173340 60412
rect 173396 60410 173420 60412
rect 173258 60358 173260 60410
rect 173322 60358 173334 60410
rect 173396 60358 173398 60410
rect 173236 60356 173260 60358
rect 173316 60356 173340 60358
rect 173396 60356 173420 60358
rect 173180 60336 173476 60356
rect 176936 60172 176988 60178
rect 176936 60114 176988 60120
rect 157820 59868 158116 59888
rect 157876 59866 157900 59868
rect 157956 59866 157980 59868
rect 158036 59866 158060 59868
rect 157898 59814 157900 59866
rect 157962 59814 157974 59866
rect 158036 59814 158038 59866
rect 157876 59812 157900 59814
rect 157956 59812 157980 59814
rect 158036 59812 158060 59814
rect 157820 59792 158116 59812
rect 176948 59770 176976 60114
rect 178130 60072 178186 60081
rect 178130 60007 178132 60016
rect 178184 60007 178186 60016
rect 178132 59978 178184 59984
rect 176936 59764 176988 59770
rect 176936 59706 176988 59712
rect 173180 59324 173476 59344
rect 173236 59322 173260 59324
rect 173316 59322 173340 59324
rect 173396 59322 173420 59324
rect 173258 59270 173260 59322
rect 173322 59270 173334 59322
rect 173396 59270 173398 59322
rect 173236 59268 173260 59270
rect 173316 59268 173340 59270
rect 173396 59268 173420 59270
rect 173180 59248 173476 59268
rect 157820 58780 158116 58800
rect 157876 58778 157900 58780
rect 157956 58778 157980 58780
rect 158036 58778 158060 58780
rect 157898 58726 157900 58778
rect 157962 58726 157974 58778
rect 158036 58726 158038 58778
rect 157876 58724 157900 58726
rect 157956 58724 157980 58726
rect 158036 58724 158060 58726
rect 157820 58704 158116 58724
rect 173180 58236 173476 58256
rect 173236 58234 173260 58236
rect 173316 58234 173340 58236
rect 173396 58234 173420 58236
rect 173258 58182 173260 58234
rect 173322 58182 173334 58234
rect 173396 58182 173398 58234
rect 173236 58180 173260 58182
rect 173316 58180 173340 58182
rect 173396 58180 173420 58182
rect 173180 58160 173476 58180
rect 157820 57692 158116 57712
rect 157876 57690 157900 57692
rect 157956 57690 157980 57692
rect 158036 57690 158060 57692
rect 157898 57638 157900 57690
rect 157962 57638 157974 57690
rect 158036 57638 158038 57690
rect 157876 57636 157900 57638
rect 157956 57636 157980 57638
rect 158036 57636 158060 57638
rect 157820 57616 158116 57636
rect 173180 57148 173476 57168
rect 173236 57146 173260 57148
rect 173316 57146 173340 57148
rect 173396 57146 173420 57148
rect 173258 57094 173260 57146
rect 173322 57094 173334 57146
rect 173396 57094 173398 57146
rect 173236 57092 173260 57094
rect 173316 57092 173340 57094
rect 173396 57092 173420 57094
rect 173180 57072 173476 57092
rect 157820 56604 158116 56624
rect 157876 56602 157900 56604
rect 157956 56602 157980 56604
rect 158036 56602 158060 56604
rect 157898 56550 157900 56602
rect 157962 56550 157974 56602
rect 158036 56550 158038 56602
rect 157876 56548 157900 56550
rect 157956 56548 157980 56550
rect 158036 56548 158060 56550
rect 157820 56528 158116 56548
rect 173180 56060 173476 56080
rect 173236 56058 173260 56060
rect 173316 56058 173340 56060
rect 173396 56058 173420 56060
rect 173258 56006 173260 56058
rect 173322 56006 173334 56058
rect 173396 56006 173398 56058
rect 173236 56004 173260 56006
rect 173316 56004 173340 56006
rect 173396 56004 173420 56006
rect 173180 55984 173476 56004
rect 157820 55516 158116 55536
rect 157876 55514 157900 55516
rect 157956 55514 157980 55516
rect 158036 55514 158060 55516
rect 157898 55462 157900 55514
rect 157962 55462 157974 55514
rect 158036 55462 158038 55514
rect 157876 55460 157900 55462
rect 157956 55460 157980 55462
rect 158036 55460 158060 55462
rect 157820 55440 158116 55460
rect 173180 54972 173476 54992
rect 173236 54970 173260 54972
rect 173316 54970 173340 54972
rect 173396 54970 173420 54972
rect 173258 54918 173260 54970
rect 173322 54918 173334 54970
rect 173396 54918 173398 54970
rect 173236 54916 173260 54918
rect 173316 54916 173340 54918
rect 173396 54916 173420 54918
rect 173180 54896 173476 54916
rect 157820 54428 158116 54448
rect 157876 54426 157900 54428
rect 157956 54426 157980 54428
rect 158036 54426 158060 54428
rect 157898 54374 157900 54426
rect 157962 54374 157974 54426
rect 158036 54374 158038 54426
rect 157876 54372 157900 54374
rect 157956 54372 157980 54374
rect 158036 54372 158060 54374
rect 157820 54352 158116 54372
rect 173180 53884 173476 53904
rect 173236 53882 173260 53884
rect 173316 53882 173340 53884
rect 173396 53882 173420 53884
rect 173258 53830 173260 53882
rect 173322 53830 173334 53882
rect 173396 53830 173398 53882
rect 173236 53828 173260 53830
rect 173316 53828 173340 53830
rect 173396 53828 173420 53830
rect 173180 53808 173476 53828
rect 157820 53340 158116 53360
rect 157876 53338 157900 53340
rect 157956 53338 157980 53340
rect 158036 53338 158060 53340
rect 157898 53286 157900 53338
rect 157962 53286 157974 53338
rect 158036 53286 158038 53338
rect 157876 53284 157900 53286
rect 157956 53284 157980 53286
rect 158036 53284 158060 53286
rect 157820 53264 158116 53284
rect 173180 52796 173476 52816
rect 173236 52794 173260 52796
rect 173316 52794 173340 52796
rect 173396 52794 173420 52796
rect 173258 52742 173260 52794
rect 173322 52742 173334 52794
rect 173396 52742 173398 52794
rect 173236 52740 173260 52742
rect 173316 52740 173340 52742
rect 173396 52740 173420 52742
rect 173180 52720 173476 52740
rect 157820 52252 158116 52272
rect 157876 52250 157900 52252
rect 157956 52250 157980 52252
rect 158036 52250 158060 52252
rect 157898 52198 157900 52250
rect 157962 52198 157974 52250
rect 158036 52198 158038 52250
rect 157876 52196 157900 52198
rect 157956 52196 157980 52198
rect 158036 52196 158060 52198
rect 157820 52176 158116 52196
rect 173180 51708 173476 51728
rect 173236 51706 173260 51708
rect 173316 51706 173340 51708
rect 173396 51706 173420 51708
rect 173258 51654 173260 51706
rect 173322 51654 173334 51706
rect 173396 51654 173398 51706
rect 173236 51652 173260 51654
rect 173316 51652 173340 51654
rect 173396 51652 173420 51654
rect 173180 51632 173476 51652
rect 157820 51164 158116 51184
rect 157876 51162 157900 51164
rect 157956 51162 157980 51164
rect 158036 51162 158060 51164
rect 157898 51110 157900 51162
rect 157962 51110 157974 51162
rect 158036 51110 158038 51162
rect 157876 51108 157900 51110
rect 157956 51108 157980 51110
rect 158036 51108 158060 51110
rect 157820 51088 158116 51108
rect 173180 50620 173476 50640
rect 173236 50618 173260 50620
rect 173316 50618 173340 50620
rect 173396 50618 173420 50620
rect 173258 50566 173260 50618
rect 173322 50566 173334 50618
rect 173396 50566 173398 50618
rect 173236 50564 173260 50566
rect 173316 50564 173340 50566
rect 173396 50564 173420 50566
rect 173180 50544 173476 50564
rect 157820 50076 158116 50096
rect 157876 50074 157900 50076
rect 157956 50074 157980 50076
rect 158036 50074 158060 50076
rect 157898 50022 157900 50074
rect 157962 50022 157974 50074
rect 158036 50022 158038 50074
rect 157876 50020 157900 50022
rect 157956 50020 157980 50022
rect 158036 50020 158060 50022
rect 157820 50000 158116 50020
rect 173180 49532 173476 49552
rect 173236 49530 173260 49532
rect 173316 49530 173340 49532
rect 173396 49530 173420 49532
rect 173258 49478 173260 49530
rect 173322 49478 173334 49530
rect 173396 49478 173398 49530
rect 173236 49476 173260 49478
rect 173316 49476 173340 49478
rect 173396 49476 173420 49478
rect 173180 49456 173476 49476
rect 157820 48988 158116 49008
rect 157876 48986 157900 48988
rect 157956 48986 157980 48988
rect 158036 48986 158060 48988
rect 157898 48934 157900 48986
rect 157962 48934 157974 48986
rect 158036 48934 158038 48986
rect 157876 48932 157900 48934
rect 157956 48932 157980 48934
rect 158036 48932 158060 48934
rect 157820 48912 158116 48932
rect 173180 48444 173476 48464
rect 173236 48442 173260 48444
rect 173316 48442 173340 48444
rect 173396 48442 173420 48444
rect 173258 48390 173260 48442
rect 173322 48390 173334 48442
rect 173396 48390 173398 48442
rect 173236 48388 173260 48390
rect 173316 48388 173340 48390
rect 173396 48388 173420 48390
rect 173180 48368 173476 48388
rect 157820 47900 158116 47920
rect 157876 47898 157900 47900
rect 157956 47898 157980 47900
rect 158036 47898 158060 47900
rect 157898 47846 157900 47898
rect 157962 47846 157974 47898
rect 158036 47846 158038 47898
rect 157876 47844 157900 47846
rect 157956 47844 157980 47846
rect 158036 47844 158060 47846
rect 157820 47824 158116 47844
rect 173180 47356 173476 47376
rect 173236 47354 173260 47356
rect 173316 47354 173340 47356
rect 173396 47354 173420 47356
rect 173258 47302 173260 47354
rect 173322 47302 173334 47354
rect 173396 47302 173398 47354
rect 173236 47300 173260 47302
rect 173316 47300 173340 47302
rect 173396 47300 173420 47302
rect 173180 47280 173476 47300
rect 157820 46812 158116 46832
rect 157876 46810 157900 46812
rect 157956 46810 157980 46812
rect 158036 46810 158060 46812
rect 157898 46758 157900 46810
rect 157962 46758 157974 46810
rect 158036 46758 158038 46810
rect 157876 46756 157900 46758
rect 157956 46756 157980 46758
rect 158036 46756 158060 46758
rect 157820 46736 158116 46756
rect 173180 46268 173476 46288
rect 173236 46266 173260 46268
rect 173316 46266 173340 46268
rect 173396 46266 173420 46268
rect 173258 46214 173260 46266
rect 173322 46214 173334 46266
rect 173396 46214 173398 46266
rect 173236 46212 173260 46214
rect 173316 46212 173340 46214
rect 173396 46212 173420 46214
rect 173180 46192 173476 46212
rect 157820 45724 158116 45744
rect 157876 45722 157900 45724
rect 157956 45722 157980 45724
rect 158036 45722 158060 45724
rect 157898 45670 157900 45722
rect 157962 45670 157974 45722
rect 158036 45670 158038 45722
rect 157876 45668 157900 45670
rect 157956 45668 157980 45670
rect 158036 45668 158060 45670
rect 157820 45648 158116 45668
rect 173180 45180 173476 45200
rect 173236 45178 173260 45180
rect 173316 45178 173340 45180
rect 173396 45178 173420 45180
rect 173258 45126 173260 45178
rect 173322 45126 173334 45178
rect 173396 45126 173398 45178
rect 173236 45124 173260 45126
rect 173316 45124 173340 45126
rect 173396 45124 173420 45126
rect 173180 45104 173476 45124
rect 157820 44636 158116 44656
rect 157876 44634 157900 44636
rect 157956 44634 157980 44636
rect 158036 44634 158060 44636
rect 157898 44582 157900 44634
rect 157962 44582 157974 44634
rect 158036 44582 158038 44634
rect 157876 44580 157900 44582
rect 157956 44580 157980 44582
rect 158036 44580 158060 44582
rect 157820 44560 158116 44580
rect 173180 44092 173476 44112
rect 173236 44090 173260 44092
rect 173316 44090 173340 44092
rect 173396 44090 173420 44092
rect 173258 44038 173260 44090
rect 173322 44038 173334 44090
rect 173396 44038 173398 44090
rect 173236 44036 173260 44038
rect 173316 44036 173340 44038
rect 173396 44036 173420 44038
rect 173180 44016 173476 44036
rect 157820 43548 158116 43568
rect 157876 43546 157900 43548
rect 157956 43546 157980 43548
rect 158036 43546 158060 43548
rect 157898 43494 157900 43546
rect 157962 43494 157974 43546
rect 158036 43494 158038 43546
rect 157876 43492 157900 43494
rect 157956 43492 157980 43494
rect 158036 43492 158060 43494
rect 157820 43472 158116 43492
rect 173180 43004 173476 43024
rect 173236 43002 173260 43004
rect 173316 43002 173340 43004
rect 173396 43002 173420 43004
rect 173258 42950 173260 43002
rect 173322 42950 173334 43002
rect 173396 42950 173398 43002
rect 173236 42948 173260 42950
rect 173316 42948 173340 42950
rect 173396 42948 173420 42950
rect 173180 42928 173476 42948
rect 157820 42460 158116 42480
rect 157876 42458 157900 42460
rect 157956 42458 157980 42460
rect 158036 42458 158060 42460
rect 157898 42406 157900 42458
rect 157962 42406 157974 42458
rect 158036 42406 158038 42458
rect 157876 42404 157900 42406
rect 157956 42404 157980 42406
rect 158036 42404 158060 42406
rect 157820 42384 158116 42404
rect 173180 41916 173476 41936
rect 173236 41914 173260 41916
rect 173316 41914 173340 41916
rect 173396 41914 173420 41916
rect 173258 41862 173260 41914
rect 173322 41862 173334 41914
rect 173396 41862 173398 41914
rect 173236 41860 173260 41862
rect 173316 41860 173340 41862
rect 173396 41860 173420 41862
rect 173180 41840 173476 41860
rect 157820 41372 158116 41392
rect 157876 41370 157900 41372
rect 157956 41370 157980 41372
rect 158036 41370 158060 41372
rect 157898 41318 157900 41370
rect 157962 41318 157974 41370
rect 158036 41318 158038 41370
rect 157876 41316 157900 41318
rect 157956 41316 157980 41318
rect 158036 41316 158060 41318
rect 157820 41296 158116 41316
rect 173180 40828 173476 40848
rect 173236 40826 173260 40828
rect 173316 40826 173340 40828
rect 173396 40826 173420 40828
rect 173258 40774 173260 40826
rect 173322 40774 173334 40826
rect 173396 40774 173398 40826
rect 173236 40772 173260 40774
rect 173316 40772 173340 40774
rect 173396 40772 173420 40774
rect 173180 40752 173476 40772
rect 157820 40284 158116 40304
rect 157876 40282 157900 40284
rect 157956 40282 157980 40284
rect 158036 40282 158060 40284
rect 157898 40230 157900 40282
rect 157962 40230 157974 40282
rect 158036 40230 158038 40282
rect 157876 40228 157900 40230
rect 157956 40228 157980 40230
rect 158036 40228 158060 40230
rect 157820 40208 158116 40228
rect 173180 39740 173476 39760
rect 173236 39738 173260 39740
rect 173316 39738 173340 39740
rect 173396 39738 173420 39740
rect 173258 39686 173260 39738
rect 173322 39686 173334 39738
rect 173396 39686 173398 39738
rect 173236 39684 173260 39686
rect 173316 39684 173340 39686
rect 173396 39684 173420 39686
rect 173180 39664 173476 39684
rect 157820 39196 158116 39216
rect 157876 39194 157900 39196
rect 157956 39194 157980 39196
rect 158036 39194 158060 39196
rect 157898 39142 157900 39194
rect 157962 39142 157974 39194
rect 158036 39142 158038 39194
rect 157876 39140 157900 39142
rect 157956 39140 157980 39142
rect 158036 39140 158060 39142
rect 157820 39120 158116 39140
rect 173180 38652 173476 38672
rect 173236 38650 173260 38652
rect 173316 38650 173340 38652
rect 173396 38650 173420 38652
rect 173258 38598 173260 38650
rect 173322 38598 173334 38650
rect 173396 38598 173398 38650
rect 173236 38596 173260 38598
rect 173316 38596 173340 38598
rect 173396 38596 173420 38598
rect 173180 38576 173476 38596
rect 157820 38108 158116 38128
rect 157876 38106 157900 38108
rect 157956 38106 157980 38108
rect 158036 38106 158060 38108
rect 157898 38054 157900 38106
rect 157962 38054 157974 38106
rect 158036 38054 158038 38106
rect 157876 38052 157900 38054
rect 157956 38052 157980 38054
rect 158036 38052 158060 38054
rect 157820 38032 158116 38052
rect 173180 37564 173476 37584
rect 173236 37562 173260 37564
rect 173316 37562 173340 37564
rect 173396 37562 173420 37564
rect 173258 37510 173260 37562
rect 173322 37510 173334 37562
rect 173396 37510 173398 37562
rect 173236 37508 173260 37510
rect 173316 37508 173340 37510
rect 173396 37508 173420 37510
rect 173180 37488 173476 37508
rect 157820 37020 158116 37040
rect 157876 37018 157900 37020
rect 157956 37018 157980 37020
rect 158036 37018 158060 37020
rect 157898 36966 157900 37018
rect 157962 36966 157974 37018
rect 158036 36966 158038 37018
rect 157876 36964 157900 36966
rect 157956 36964 157980 36966
rect 158036 36964 158060 36966
rect 157820 36944 158116 36964
rect 173180 36476 173476 36496
rect 173236 36474 173260 36476
rect 173316 36474 173340 36476
rect 173396 36474 173420 36476
rect 173258 36422 173260 36474
rect 173322 36422 173334 36474
rect 173396 36422 173398 36474
rect 173236 36420 173260 36422
rect 173316 36420 173340 36422
rect 173396 36420 173420 36422
rect 173180 36400 173476 36420
rect 157820 35932 158116 35952
rect 157876 35930 157900 35932
rect 157956 35930 157980 35932
rect 158036 35930 158060 35932
rect 157898 35878 157900 35930
rect 157962 35878 157974 35930
rect 158036 35878 158038 35930
rect 157876 35876 157900 35878
rect 157956 35876 157980 35878
rect 158036 35876 158060 35878
rect 157820 35856 158116 35876
rect 173180 35388 173476 35408
rect 173236 35386 173260 35388
rect 173316 35386 173340 35388
rect 173396 35386 173420 35388
rect 173258 35334 173260 35386
rect 173322 35334 173334 35386
rect 173396 35334 173398 35386
rect 173236 35332 173260 35334
rect 173316 35332 173340 35334
rect 173396 35332 173420 35334
rect 173180 35312 173476 35332
rect 157820 34844 158116 34864
rect 157876 34842 157900 34844
rect 157956 34842 157980 34844
rect 158036 34842 158060 34844
rect 157898 34790 157900 34842
rect 157962 34790 157974 34842
rect 158036 34790 158038 34842
rect 157876 34788 157900 34790
rect 157956 34788 157980 34790
rect 158036 34788 158060 34790
rect 157820 34768 158116 34788
rect 173180 34300 173476 34320
rect 173236 34298 173260 34300
rect 173316 34298 173340 34300
rect 173396 34298 173420 34300
rect 173258 34246 173260 34298
rect 173322 34246 173334 34298
rect 173396 34246 173398 34298
rect 173236 34244 173260 34246
rect 173316 34244 173340 34246
rect 173396 34244 173420 34246
rect 173180 34224 173476 34244
rect 157820 33756 158116 33776
rect 157876 33754 157900 33756
rect 157956 33754 157980 33756
rect 158036 33754 158060 33756
rect 157898 33702 157900 33754
rect 157962 33702 157974 33754
rect 158036 33702 158038 33754
rect 157876 33700 157900 33702
rect 157956 33700 157980 33702
rect 158036 33700 158060 33702
rect 157820 33680 158116 33700
rect 173180 33212 173476 33232
rect 173236 33210 173260 33212
rect 173316 33210 173340 33212
rect 173396 33210 173420 33212
rect 173258 33158 173260 33210
rect 173322 33158 173334 33210
rect 173396 33158 173398 33210
rect 173236 33156 173260 33158
rect 173316 33156 173340 33158
rect 173396 33156 173420 33158
rect 173180 33136 173476 33156
rect 157820 32668 158116 32688
rect 157876 32666 157900 32668
rect 157956 32666 157980 32668
rect 158036 32666 158060 32668
rect 157898 32614 157900 32666
rect 157962 32614 157974 32666
rect 158036 32614 158038 32666
rect 157876 32612 157900 32614
rect 157956 32612 157980 32614
rect 158036 32612 158060 32614
rect 157820 32592 158116 32612
rect 173180 32124 173476 32144
rect 173236 32122 173260 32124
rect 173316 32122 173340 32124
rect 173396 32122 173420 32124
rect 173258 32070 173260 32122
rect 173322 32070 173334 32122
rect 173396 32070 173398 32122
rect 173236 32068 173260 32070
rect 173316 32068 173340 32070
rect 173396 32068 173420 32070
rect 173180 32048 173476 32068
rect 157820 31580 158116 31600
rect 157876 31578 157900 31580
rect 157956 31578 157980 31580
rect 158036 31578 158060 31580
rect 157898 31526 157900 31578
rect 157962 31526 157974 31578
rect 158036 31526 158038 31578
rect 157876 31524 157900 31526
rect 157956 31524 157980 31526
rect 158036 31524 158060 31526
rect 157820 31504 158116 31524
rect 173180 31036 173476 31056
rect 173236 31034 173260 31036
rect 173316 31034 173340 31036
rect 173396 31034 173420 31036
rect 173258 30982 173260 31034
rect 173322 30982 173334 31034
rect 173396 30982 173398 31034
rect 173236 30980 173260 30982
rect 173316 30980 173340 30982
rect 173396 30980 173420 30982
rect 173180 30960 173476 30980
rect 157820 30492 158116 30512
rect 157876 30490 157900 30492
rect 157956 30490 157980 30492
rect 158036 30490 158060 30492
rect 157898 30438 157900 30490
rect 157962 30438 157974 30490
rect 158036 30438 158038 30490
rect 157876 30436 157900 30438
rect 157956 30436 157980 30438
rect 158036 30436 158060 30438
rect 157820 30416 158116 30436
rect 173180 29948 173476 29968
rect 173236 29946 173260 29948
rect 173316 29946 173340 29948
rect 173396 29946 173420 29948
rect 173258 29894 173260 29946
rect 173322 29894 173334 29946
rect 173396 29894 173398 29946
rect 173236 29892 173260 29894
rect 173316 29892 173340 29894
rect 173396 29892 173420 29894
rect 173180 29872 173476 29892
rect 157820 29404 158116 29424
rect 157876 29402 157900 29404
rect 157956 29402 157980 29404
rect 158036 29402 158060 29404
rect 157898 29350 157900 29402
rect 157962 29350 157974 29402
rect 158036 29350 158038 29402
rect 157876 29348 157900 29350
rect 157956 29348 157980 29350
rect 158036 29348 158060 29350
rect 157820 29328 158116 29348
rect 173180 28860 173476 28880
rect 173236 28858 173260 28860
rect 173316 28858 173340 28860
rect 173396 28858 173420 28860
rect 173258 28806 173260 28858
rect 173322 28806 173334 28858
rect 173396 28806 173398 28858
rect 173236 28804 173260 28806
rect 173316 28804 173340 28806
rect 173396 28804 173420 28806
rect 173180 28784 173476 28804
rect 157820 28316 158116 28336
rect 157876 28314 157900 28316
rect 157956 28314 157980 28316
rect 158036 28314 158060 28316
rect 157898 28262 157900 28314
rect 157962 28262 157974 28314
rect 158036 28262 158038 28314
rect 157876 28260 157900 28262
rect 157956 28260 157980 28262
rect 158036 28260 158060 28262
rect 157820 28240 158116 28260
rect 173180 27772 173476 27792
rect 173236 27770 173260 27772
rect 173316 27770 173340 27772
rect 173396 27770 173420 27772
rect 173258 27718 173260 27770
rect 173322 27718 173334 27770
rect 173396 27718 173398 27770
rect 173236 27716 173260 27718
rect 173316 27716 173340 27718
rect 173396 27716 173420 27718
rect 173180 27696 173476 27716
rect 157820 27228 158116 27248
rect 157876 27226 157900 27228
rect 157956 27226 157980 27228
rect 158036 27226 158060 27228
rect 157898 27174 157900 27226
rect 157962 27174 157974 27226
rect 158036 27174 158038 27226
rect 157876 27172 157900 27174
rect 157956 27172 157980 27174
rect 158036 27172 158060 27174
rect 157820 27152 158116 27172
rect 173180 26684 173476 26704
rect 173236 26682 173260 26684
rect 173316 26682 173340 26684
rect 173396 26682 173420 26684
rect 173258 26630 173260 26682
rect 173322 26630 173334 26682
rect 173396 26630 173398 26682
rect 173236 26628 173260 26630
rect 173316 26628 173340 26630
rect 173396 26628 173420 26630
rect 173180 26608 173476 26628
rect 157820 26140 158116 26160
rect 157876 26138 157900 26140
rect 157956 26138 157980 26140
rect 158036 26138 158060 26140
rect 157898 26086 157900 26138
rect 157962 26086 157974 26138
rect 158036 26086 158038 26138
rect 157876 26084 157900 26086
rect 157956 26084 157980 26086
rect 158036 26084 158060 26086
rect 157820 26064 158116 26084
rect 173180 25596 173476 25616
rect 173236 25594 173260 25596
rect 173316 25594 173340 25596
rect 173396 25594 173420 25596
rect 173258 25542 173260 25594
rect 173322 25542 173334 25594
rect 173396 25542 173398 25594
rect 173236 25540 173260 25542
rect 173316 25540 173340 25542
rect 173396 25540 173420 25542
rect 173180 25520 173476 25540
rect 157820 25052 158116 25072
rect 157876 25050 157900 25052
rect 157956 25050 157980 25052
rect 158036 25050 158060 25052
rect 157898 24998 157900 25050
rect 157962 24998 157974 25050
rect 158036 24998 158038 25050
rect 157876 24996 157900 24998
rect 157956 24996 157980 24998
rect 158036 24996 158060 24998
rect 157820 24976 158116 24996
rect 173180 24508 173476 24528
rect 173236 24506 173260 24508
rect 173316 24506 173340 24508
rect 173396 24506 173420 24508
rect 173258 24454 173260 24506
rect 173322 24454 173334 24506
rect 173396 24454 173398 24506
rect 173236 24452 173260 24454
rect 173316 24452 173340 24454
rect 173396 24452 173420 24454
rect 173180 24432 173476 24452
rect 157820 23964 158116 23984
rect 157876 23962 157900 23964
rect 157956 23962 157980 23964
rect 158036 23962 158060 23964
rect 157898 23910 157900 23962
rect 157962 23910 157974 23962
rect 158036 23910 158038 23962
rect 157876 23908 157900 23910
rect 157956 23908 157980 23910
rect 158036 23908 158060 23910
rect 157820 23888 158116 23908
rect 173180 23420 173476 23440
rect 173236 23418 173260 23420
rect 173316 23418 173340 23420
rect 173396 23418 173420 23420
rect 173258 23366 173260 23418
rect 173322 23366 173334 23418
rect 173396 23366 173398 23418
rect 173236 23364 173260 23366
rect 173316 23364 173340 23366
rect 173396 23364 173420 23366
rect 173180 23344 173476 23364
rect 157820 22876 158116 22896
rect 157876 22874 157900 22876
rect 157956 22874 157980 22876
rect 158036 22874 158060 22876
rect 157898 22822 157900 22874
rect 157962 22822 157974 22874
rect 158036 22822 158038 22874
rect 157876 22820 157900 22822
rect 157956 22820 157980 22822
rect 158036 22820 158060 22822
rect 157820 22800 158116 22820
rect 173180 22332 173476 22352
rect 173236 22330 173260 22332
rect 173316 22330 173340 22332
rect 173396 22330 173420 22332
rect 173258 22278 173260 22330
rect 173322 22278 173334 22330
rect 173396 22278 173398 22330
rect 173236 22276 173260 22278
rect 173316 22276 173340 22278
rect 173396 22276 173420 22278
rect 173180 22256 173476 22276
rect 157820 21788 158116 21808
rect 157876 21786 157900 21788
rect 157956 21786 157980 21788
rect 158036 21786 158060 21788
rect 157898 21734 157900 21786
rect 157962 21734 157974 21786
rect 158036 21734 158038 21786
rect 157876 21732 157900 21734
rect 157956 21732 157980 21734
rect 158036 21732 158060 21734
rect 157820 21712 158116 21732
rect 173180 21244 173476 21264
rect 173236 21242 173260 21244
rect 173316 21242 173340 21244
rect 173396 21242 173420 21244
rect 173258 21190 173260 21242
rect 173322 21190 173334 21242
rect 173396 21190 173398 21242
rect 173236 21188 173260 21190
rect 173316 21188 173340 21190
rect 173396 21188 173420 21190
rect 173180 21168 173476 21188
rect 157820 20700 158116 20720
rect 157876 20698 157900 20700
rect 157956 20698 157980 20700
rect 158036 20698 158060 20700
rect 157898 20646 157900 20698
rect 157962 20646 157974 20698
rect 158036 20646 158038 20698
rect 157876 20644 157900 20646
rect 157956 20644 157980 20646
rect 158036 20644 158060 20646
rect 157820 20624 158116 20644
rect 149520 20392 149572 20398
rect 149520 20334 149572 20340
rect 173180 20156 173476 20176
rect 173236 20154 173260 20156
rect 173316 20154 173340 20156
rect 173396 20154 173420 20156
rect 173258 20102 173260 20154
rect 173322 20102 173334 20154
rect 173396 20102 173398 20154
rect 173236 20100 173260 20102
rect 173316 20100 173340 20102
rect 173396 20100 173420 20102
rect 173180 20080 173476 20100
rect 157820 19612 158116 19632
rect 157876 19610 157900 19612
rect 157956 19610 157980 19612
rect 158036 19610 158060 19612
rect 157898 19558 157900 19610
rect 157962 19558 157974 19610
rect 158036 19558 158038 19610
rect 157876 19556 157900 19558
rect 157956 19556 157980 19558
rect 158036 19556 158060 19558
rect 157820 19536 158116 19556
rect 173180 19068 173476 19088
rect 173236 19066 173260 19068
rect 173316 19066 173340 19068
rect 173396 19066 173420 19068
rect 173258 19014 173260 19066
rect 173322 19014 173334 19066
rect 173396 19014 173398 19066
rect 173236 19012 173260 19014
rect 173316 19012 173340 19014
rect 173396 19012 173420 19014
rect 173180 18992 173476 19012
rect 144552 18828 144604 18834
rect 144552 18770 144604 18776
rect 75828 18624 75880 18630
rect 75828 18566 75880 18572
rect 96380 18524 96676 18544
rect 96436 18522 96460 18524
rect 96516 18522 96540 18524
rect 96596 18522 96620 18524
rect 96458 18470 96460 18522
rect 96522 18470 96534 18522
rect 96596 18470 96598 18522
rect 96436 18468 96460 18470
rect 96516 18468 96540 18470
rect 96596 18468 96620 18470
rect 96380 18448 96676 18468
rect 127100 18524 127396 18544
rect 127156 18522 127180 18524
rect 127236 18522 127260 18524
rect 127316 18522 127340 18524
rect 127178 18470 127180 18522
rect 127242 18470 127254 18522
rect 127316 18470 127318 18522
rect 127156 18468 127180 18470
rect 127236 18468 127260 18470
rect 127316 18468 127340 18470
rect 127100 18448 127396 18468
rect 157820 18524 158116 18544
rect 157876 18522 157900 18524
rect 157956 18522 157980 18524
rect 158036 18522 158060 18524
rect 157898 18470 157900 18522
rect 157962 18470 157974 18522
rect 158036 18470 158038 18522
rect 157876 18468 157900 18470
rect 157956 18468 157980 18470
rect 158036 18468 158060 18470
rect 157820 18448 158116 18468
rect 81020 17980 81316 18000
rect 81076 17978 81100 17980
rect 81156 17978 81180 17980
rect 81236 17978 81260 17980
rect 81098 17926 81100 17978
rect 81162 17926 81174 17978
rect 81236 17926 81238 17978
rect 81076 17924 81100 17926
rect 81156 17924 81180 17926
rect 81236 17924 81260 17926
rect 81020 17904 81316 17924
rect 111740 17980 112036 18000
rect 111796 17978 111820 17980
rect 111876 17978 111900 17980
rect 111956 17978 111980 17980
rect 111818 17926 111820 17978
rect 111882 17926 111894 17978
rect 111956 17926 111958 17978
rect 111796 17924 111820 17926
rect 111876 17924 111900 17926
rect 111956 17924 111980 17926
rect 111740 17904 112036 17924
rect 142460 17980 142756 18000
rect 142516 17978 142540 17980
rect 142596 17978 142620 17980
rect 142676 17978 142700 17980
rect 142538 17926 142540 17978
rect 142602 17926 142614 17978
rect 142676 17926 142678 17978
rect 142516 17924 142540 17926
rect 142596 17924 142620 17926
rect 142676 17924 142700 17926
rect 142460 17904 142756 17924
rect 173180 17980 173476 18000
rect 173236 17978 173260 17980
rect 173316 17978 173340 17980
rect 173396 17978 173420 17980
rect 173258 17926 173260 17978
rect 173322 17926 173334 17978
rect 173396 17926 173398 17978
rect 173236 17924 173260 17926
rect 173316 17924 173340 17926
rect 173396 17924 173420 17926
rect 173180 17904 173476 17924
rect 96380 17436 96676 17456
rect 96436 17434 96460 17436
rect 96516 17434 96540 17436
rect 96596 17434 96620 17436
rect 96458 17382 96460 17434
rect 96522 17382 96534 17434
rect 96596 17382 96598 17434
rect 96436 17380 96460 17382
rect 96516 17380 96540 17382
rect 96596 17380 96620 17382
rect 96380 17360 96676 17380
rect 127100 17436 127396 17456
rect 127156 17434 127180 17436
rect 127236 17434 127260 17436
rect 127316 17434 127340 17436
rect 127178 17382 127180 17434
rect 127242 17382 127254 17434
rect 127316 17382 127318 17434
rect 127156 17380 127180 17382
rect 127236 17380 127260 17382
rect 127316 17380 127340 17382
rect 127100 17360 127396 17380
rect 157820 17436 158116 17456
rect 157876 17434 157900 17436
rect 157956 17434 157980 17436
rect 158036 17434 158060 17436
rect 157898 17382 157900 17434
rect 157962 17382 157974 17434
rect 158036 17382 158038 17434
rect 157876 17380 157900 17382
rect 157956 17380 157980 17382
rect 158036 17380 158060 17382
rect 157820 17360 158116 17380
rect 81020 16892 81316 16912
rect 81076 16890 81100 16892
rect 81156 16890 81180 16892
rect 81236 16890 81260 16892
rect 81098 16838 81100 16890
rect 81162 16838 81174 16890
rect 81236 16838 81238 16890
rect 81076 16836 81100 16838
rect 81156 16836 81180 16838
rect 81236 16836 81260 16838
rect 81020 16816 81316 16836
rect 111740 16892 112036 16912
rect 111796 16890 111820 16892
rect 111876 16890 111900 16892
rect 111956 16890 111980 16892
rect 111818 16838 111820 16890
rect 111882 16838 111894 16890
rect 111956 16838 111958 16890
rect 111796 16836 111820 16838
rect 111876 16836 111900 16838
rect 111956 16836 111980 16838
rect 111740 16816 112036 16836
rect 142460 16892 142756 16912
rect 142516 16890 142540 16892
rect 142596 16890 142620 16892
rect 142676 16890 142700 16892
rect 142538 16838 142540 16890
rect 142602 16838 142614 16890
rect 142676 16838 142678 16890
rect 142516 16836 142540 16838
rect 142596 16836 142620 16838
rect 142676 16836 142700 16838
rect 142460 16816 142756 16836
rect 173180 16892 173476 16912
rect 173236 16890 173260 16892
rect 173316 16890 173340 16892
rect 173396 16890 173420 16892
rect 173258 16838 173260 16890
rect 173322 16838 173334 16890
rect 173396 16838 173398 16890
rect 173236 16836 173260 16838
rect 173316 16836 173340 16838
rect 173396 16836 173420 16838
rect 173180 16816 173476 16836
rect 75276 16652 75328 16658
rect 75276 16594 75328 16600
rect 96380 16348 96676 16368
rect 96436 16346 96460 16348
rect 96516 16346 96540 16348
rect 96596 16346 96620 16348
rect 96458 16294 96460 16346
rect 96522 16294 96534 16346
rect 96596 16294 96598 16346
rect 96436 16292 96460 16294
rect 96516 16292 96540 16294
rect 96596 16292 96620 16294
rect 96380 16272 96676 16292
rect 127100 16348 127396 16368
rect 127156 16346 127180 16348
rect 127236 16346 127260 16348
rect 127316 16346 127340 16348
rect 127178 16294 127180 16346
rect 127242 16294 127254 16346
rect 127316 16294 127318 16346
rect 127156 16292 127180 16294
rect 127236 16292 127260 16294
rect 127316 16292 127340 16294
rect 127100 16272 127396 16292
rect 157820 16348 158116 16368
rect 157876 16346 157900 16348
rect 157956 16346 157980 16348
rect 158036 16346 158060 16348
rect 157898 16294 157900 16346
rect 157962 16294 157974 16346
rect 158036 16294 158038 16346
rect 157876 16292 157900 16294
rect 157956 16292 157980 16294
rect 158036 16292 158060 16294
rect 157820 16272 158116 16292
rect 81020 15804 81316 15824
rect 81076 15802 81100 15804
rect 81156 15802 81180 15804
rect 81236 15802 81260 15804
rect 81098 15750 81100 15802
rect 81162 15750 81174 15802
rect 81236 15750 81238 15802
rect 81076 15748 81100 15750
rect 81156 15748 81180 15750
rect 81236 15748 81260 15750
rect 81020 15728 81316 15748
rect 111740 15804 112036 15824
rect 111796 15802 111820 15804
rect 111876 15802 111900 15804
rect 111956 15802 111980 15804
rect 111818 15750 111820 15802
rect 111882 15750 111894 15802
rect 111956 15750 111958 15802
rect 111796 15748 111820 15750
rect 111876 15748 111900 15750
rect 111956 15748 111980 15750
rect 111740 15728 112036 15748
rect 142460 15804 142756 15824
rect 142516 15802 142540 15804
rect 142596 15802 142620 15804
rect 142676 15802 142700 15804
rect 142538 15750 142540 15802
rect 142602 15750 142614 15802
rect 142676 15750 142678 15802
rect 142516 15748 142540 15750
rect 142596 15748 142620 15750
rect 142676 15748 142700 15750
rect 142460 15728 142756 15748
rect 173180 15804 173476 15824
rect 173236 15802 173260 15804
rect 173316 15802 173340 15804
rect 173396 15802 173420 15804
rect 173258 15750 173260 15802
rect 173322 15750 173334 15802
rect 173396 15750 173398 15802
rect 173236 15748 173260 15750
rect 173316 15748 173340 15750
rect 173396 15748 173420 15750
rect 173180 15728 173476 15748
rect 96380 15260 96676 15280
rect 96436 15258 96460 15260
rect 96516 15258 96540 15260
rect 96596 15258 96620 15260
rect 96458 15206 96460 15258
rect 96522 15206 96534 15258
rect 96596 15206 96598 15258
rect 96436 15204 96460 15206
rect 96516 15204 96540 15206
rect 96596 15204 96620 15206
rect 96380 15184 96676 15204
rect 127100 15260 127396 15280
rect 127156 15258 127180 15260
rect 127236 15258 127260 15260
rect 127316 15258 127340 15260
rect 127178 15206 127180 15258
rect 127242 15206 127254 15258
rect 127316 15206 127318 15258
rect 127156 15204 127180 15206
rect 127236 15204 127260 15206
rect 127316 15204 127340 15206
rect 127100 15184 127396 15204
rect 157820 15260 158116 15280
rect 157876 15258 157900 15260
rect 157956 15258 157980 15260
rect 158036 15258 158060 15260
rect 157898 15206 157900 15258
rect 157962 15206 157974 15258
rect 158036 15206 158038 15258
rect 157876 15204 157900 15206
rect 157956 15204 157980 15206
rect 158036 15204 158060 15206
rect 157820 15184 158116 15204
rect 81020 14716 81316 14736
rect 81076 14714 81100 14716
rect 81156 14714 81180 14716
rect 81236 14714 81260 14716
rect 81098 14662 81100 14714
rect 81162 14662 81174 14714
rect 81236 14662 81238 14714
rect 81076 14660 81100 14662
rect 81156 14660 81180 14662
rect 81236 14660 81260 14662
rect 81020 14640 81316 14660
rect 111740 14716 112036 14736
rect 111796 14714 111820 14716
rect 111876 14714 111900 14716
rect 111956 14714 111980 14716
rect 111818 14662 111820 14714
rect 111882 14662 111894 14714
rect 111956 14662 111958 14714
rect 111796 14660 111820 14662
rect 111876 14660 111900 14662
rect 111956 14660 111980 14662
rect 111740 14640 112036 14660
rect 142460 14716 142756 14736
rect 142516 14714 142540 14716
rect 142596 14714 142620 14716
rect 142676 14714 142700 14716
rect 142538 14662 142540 14714
rect 142602 14662 142614 14714
rect 142676 14662 142678 14714
rect 142516 14660 142540 14662
rect 142596 14660 142620 14662
rect 142676 14660 142700 14662
rect 142460 14640 142756 14660
rect 173180 14716 173476 14736
rect 173236 14714 173260 14716
rect 173316 14714 173340 14716
rect 173396 14714 173420 14716
rect 173258 14662 173260 14714
rect 173322 14662 173334 14714
rect 173396 14662 173398 14714
rect 173236 14660 173260 14662
rect 173316 14660 173340 14662
rect 173396 14660 173420 14662
rect 173180 14640 173476 14660
rect 74356 14476 74408 14482
rect 74356 14418 74408 14424
rect 101312 14340 101364 14346
rect 101312 14282 101364 14288
rect 96380 14172 96676 14192
rect 96436 14170 96460 14172
rect 96516 14170 96540 14172
rect 96596 14170 96620 14172
rect 96458 14118 96460 14170
rect 96522 14118 96534 14170
rect 96596 14118 96598 14170
rect 96436 14116 96460 14118
rect 96516 14116 96540 14118
rect 96596 14116 96620 14118
rect 96380 14096 96676 14116
rect 81020 13628 81316 13648
rect 81076 13626 81100 13628
rect 81156 13626 81180 13628
rect 81236 13626 81260 13628
rect 81098 13574 81100 13626
rect 81162 13574 81174 13626
rect 81236 13574 81238 13626
rect 81076 13572 81100 13574
rect 81156 13572 81180 13574
rect 81236 13572 81260 13574
rect 81020 13552 81316 13572
rect 73068 13388 73120 13394
rect 73068 13330 73120 13336
rect 73896 13320 73948 13326
rect 73896 13262 73948 13268
rect 72976 12776 73028 12782
rect 72976 12718 73028 12724
rect 71136 11348 71188 11354
rect 71136 11290 71188 11296
rect 72516 9648 72568 9654
rect 72516 9590 72568 9596
rect 71320 8288 71372 8294
rect 71320 8230 71372 8236
rect 70952 6928 71004 6934
rect 70952 6870 71004 6876
rect 70676 6860 70728 6866
rect 70676 6802 70728 6808
rect 71332 6254 71360 8230
rect 71320 6248 71372 6254
rect 70308 6190 70360 6196
rect 70398 6216 70454 6225
rect 71320 6190 71372 6196
rect 70398 6151 70454 6160
rect 71136 6112 71188 6118
rect 71136 6054 71188 6060
rect 70216 5704 70268 5710
rect 70216 5646 70268 5652
rect 70032 3392 70084 3398
rect 70032 3334 70084 3340
rect 69940 3188 69992 3194
rect 69940 3130 69992 3136
rect 70032 3120 70084 3126
rect 70030 3088 70032 3097
rect 70084 3088 70086 3097
rect 70030 3023 70086 3032
rect 70228 2922 70256 5646
rect 70584 4684 70636 4690
rect 70584 4626 70636 4632
rect 70400 3936 70452 3942
rect 70400 3878 70452 3884
rect 70412 3126 70440 3878
rect 70492 3392 70544 3398
rect 70492 3334 70544 3340
rect 70308 3120 70360 3126
rect 70308 3062 70360 3068
rect 70400 3120 70452 3126
rect 70400 3062 70452 3068
rect 70216 2916 70268 2922
rect 70216 2858 70268 2864
rect 69940 2508 69992 2514
rect 69940 2450 69992 2456
rect 69952 1306 69980 2450
rect 70216 2304 70268 2310
rect 70216 2246 70268 2252
rect 69860 1278 69980 1306
rect 69572 1148 69624 1154
rect 69572 1090 69624 1096
rect 69860 800 69888 1278
rect 70228 800 70256 2246
rect 70320 1358 70348 3062
rect 70504 2961 70532 3334
rect 70490 2952 70546 2961
rect 70490 2887 70546 2896
rect 70308 1352 70360 1358
rect 70308 1294 70360 1300
rect 70596 800 70624 4626
rect 71044 4140 71096 4146
rect 71044 4082 71096 4088
rect 70952 4072 71004 4078
rect 70952 4014 71004 4020
rect 70860 4004 70912 4010
rect 70860 3946 70912 3952
rect 70676 3732 70728 3738
rect 70676 3674 70728 3680
rect 70768 3732 70820 3738
rect 70768 3674 70820 3680
rect 70688 3233 70716 3674
rect 70674 3224 70730 3233
rect 70674 3159 70730 3168
rect 70780 3058 70808 3674
rect 70872 3602 70900 3946
rect 70860 3596 70912 3602
rect 70860 3538 70912 3544
rect 70768 3052 70820 3058
rect 70768 2994 70820 3000
rect 70964 800 70992 4014
rect 71056 3942 71084 4082
rect 71044 3936 71096 3942
rect 71044 3878 71096 3884
rect 71148 2650 71176 6054
rect 72056 5840 72108 5846
rect 72056 5782 72108 5788
rect 72068 5370 72096 5782
rect 72056 5364 72108 5370
rect 72056 5306 72108 5312
rect 71964 5092 72016 5098
rect 71964 5034 72016 5040
rect 71780 4684 71832 4690
rect 71780 4626 71832 4632
rect 71228 4072 71280 4078
rect 71228 4014 71280 4020
rect 71240 3602 71268 4014
rect 71412 4004 71464 4010
rect 71412 3946 71464 3952
rect 71228 3596 71280 3602
rect 71228 3538 71280 3544
rect 71424 3482 71452 3946
rect 71504 3936 71556 3942
rect 71502 3904 71504 3913
rect 71556 3904 71558 3913
rect 71502 3839 71558 3848
rect 71240 3454 71452 3482
rect 71240 3398 71268 3454
rect 71228 3392 71280 3398
rect 71228 3334 71280 3340
rect 71596 2984 71648 2990
rect 71318 2952 71374 2961
rect 71318 2887 71320 2896
rect 71372 2887 71374 2896
rect 71516 2944 71596 2972
rect 71320 2858 71372 2864
rect 71136 2644 71188 2650
rect 71136 2586 71188 2592
rect 71320 2644 71372 2650
rect 71320 2586 71372 2592
rect 71332 800 71360 2586
rect 71412 2372 71464 2378
rect 71412 2314 71464 2320
rect 71424 1562 71452 2314
rect 71412 1556 71464 1562
rect 71412 1498 71464 1504
rect 71516 1290 71544 2944
rect 71596 2926 71648 2932
rect 71596 2848 71648 2854
rect 71596 2790 71648 2796
rect 71608 1902 71636 2790
rect 71792 2774 71820 4626
rect 71872 3188 71924 3194
rect 71872 3130 71924 3136
rect 71700 2746 71820 2774
rect 71596 1896 71648 1902
rect 71596 1838 71648 1844
rect 71504 1284 71556 1290
rect 71504 1226 71556 1232
rect 71700 800 71728 2746
rect 71884 2310 71912 3130
rect 71976 3097 72004 5034
rect 72056 4072 72108 4078
rect 72056 4014 72108 4020
rect 71962 3088 72018 3097
rect 71962 3023 72018 3032
rect 71872 2304 71924 2310
rect 71872 2246 71924 2252
rect 71964 2304 72016 2310
rect 71964 2246 72016 2252
rect 71976 2038 72004 2246
rect 71964 2032 72016 2038
rect 71964 1974 72016 1980
rect 72068 800 72096 4014
rect 72424 3664 72476 3670
rect 72146 3632 72202 3641
rect 72424 3606 72476 3612
rect 72146 3567 72202 3576
rect 72160 2990 72188 3567
rect 72332 3392 72384 3398
rect 72332 3334 72384 3340
rect 72344 3194 72372 3334
rect 72332 3188 72384 3194
rect 72332 3130 72384 3136
rect 72436 3074 72464 3606
rect 72528 3194 72556 9590
rect 72608 7948 72660 7954
rect 72608 7890 72660 7896
rect 72620 5778 72648 7890
rect 73250 6216 73306 6225
rect 73250 6151 73306 6160
rect 73264 5778 73292 6151
rect 73620 6112 73672 6118
rect 73620 6054 73672 6060
rect 72608 5772 72660 5778
rect 72608 5714 72660 5720
rect 73252 5772 73304 5778
rect 73252 5714 73304 5720
rect 72792 4684 72844 4690
rect 72792 4626 72844 4632
rect 72700 3732 72752 3738
rect 72700 3674 72752 3680
rect 72712 3466 72740 3674
rect 72700 3460 72752 3466
rect 72700 3402 72752 3408
rect 72516 3188 72568 3194
rect 72516 3130 72568 3136
rect 72608 3188 72660 3194
rect 72608 3130 72660 3136
rect 72620 3074 72648 3130
rect 72436 3046 72648 3074
rect 72148 2984 72200 2990
rect 72148 2926 72200 2932
rect 72424 2304 72476 2310
rect 72424 2246 72476 2252
rect 72436 800 72464 2246
rect 72804 800 72832 4626
rect 73436 4140 73488 4146
rect 73436 4082 73488 4088
rect 73160 4072 73212 4078
rect 73160 4014 73212 4020
rect 73250 4040 73306 4049
rect 72976 3392 73028 3398
rect 72976 3334 73028 3340
rect 72988 2106 73016 3334
rect 72976 2100 73028 2106
rect 72976 2042 73028 2048
rect 73172 800 73200 4014
rect 73250 3975 73306 3984
rect 73264 3738 73292 3975
rect 73252 3732 73304 3738
rect 73252 3674 73304 3680
rect 73448 3602 73476 4082
rect 73436 3596 73488 3602
rect 73436 3538 73488 3544
rect 73434 3088 73490 3097
rect 73434 3023 73490 3032
rect 73448 2854 73476 3023
rect 73632 2990 73660 6054
rect 73712 5908 73764 5914
rect 73712 5850 73764 5856
rect 73620 2984 73672 2990
rect 73620 2926 73672 2932
rect 73436 2848 73488 2854
rect 73436 2790 73488 2796
rect 73528 2848 73580 2854
rect 73528 2790 73580 2796
rect 73436 2576 73488 2582
rect 73436 2518 73488 2524
rect 73448 1630 73476 2518
rect 73436 1624 73488 1630
rect 73436 1566 73488 1572
rect 73540 800 73568 2790
rect 73724 2582 73752 5850
rect 73804 5568 73856 5574
rect 73804 5510 73856 5516
rect 73816 2582 73844 5510
rect 73908 4826 73936 13262
rect 96380 13084 96676 13104
rect 96436 13082 96460 13084
rect 96516 13082 96540 13084
rect 96596 13082 96620 13084
rect 96458 13030 96460 13082
rect 96522 13030 96534 13082
rect 96596 13030 96598 13082
rect 96436 13028 96460 13030
rect 96516 13028 96540 13030
rect 96596 13028 96620 13030
rect 96380 13008 96676 13028
rect 81020 12540 81316 12560
rect 81076 12538 81100 12540
rect 81156 12538 81180 12540
rect 81236 12538 81260 12540
rect 81098 12486 81100 12538
rect 81162 12486 81174 12538
rect 81236 12486 81238 12538
rect 81076 12484 81100 12486
rect 81156 12484 81180 12486
rect 81236 12484 81260 12486
rect 81020 12464 81316 12484
rect 93952 12300 94004 12306
rect 93952 12242 94004 12248
rect 81020 11452 81316 11472
rect 81076 11450 81100 11452
rect 81156 11450 81180 11452
rect 81236 11450 81260 11452
rect 81098 11398 81100 11450
rect 81162 11398 81174 11450
rect 81236 11398 81238 11450
rect 81076 11396 81100 11398
rect 81156 11396 81180 11398
rect 81236 11396 81260 11398
rect 81020 11376 81316 11396
rect 81020 10364 81316 10384
rect 81076 10362 81100 10364
rect 81156 10362 81180 10364
rect 81236 10362 81260 10364
rect 81098 10310 81100 10362
rect 81162 10310 81174 10362
rect 81236 10310 81238 10362
rect 81076 10308 81100 10310
rect 81156 10308 81180 10310
rect 81236 10308 81260 10310
rect 81020 10288 81316 10308
rect 81020 9276 81316 9296
rect 81076 9274 81100 9276
rect 81156 9274 81180 9276
rect 81236 9274 81260 9276
rect 81098 9222 81100 9274
rect 81162 9222 81174 9274
rect 81236 9222 81238 9274
rect 81076 9220 81100 9222
rect 81156 9220 81180 9222
rect 81236 9220 81260 9222
rect 81020 9200 81316 9220
rect 81020 8188 81316 8208
rect 81076 8186 81100 8188
rect 81156 8186 81180 8188
rect 81236 8186 81260 8188
rect 81098 8134 81100 8186
rect 81162 8134 81174 8186
rect 81236 8134 81238 8186
rect 81076 8132 81100 8134
rect 81156 8132 81180 8134
rect 81236 8132 81260 8134
rect 81020 8112 81316 8132
rect 86592 7336 86644 7342
rect 86592 7278 86644 7284
rect 81020 7100 81316 7120
rect 81076 7098 81100 7100
rect 81156 7098 81180 7100
rect 81236 7098 81260 7100
rect 81098 7046 81100 7098
rect 81162 7046 81174 7098
rect 81236 7046 81238 7098
rect 81076 7044 81100 7046
rect 81156 7044 81180 7046
rect 81236 7044 81260 7046
rect 81020 7024 81316 7044
rect 84844 6996 84896 7002
rect 84844 6938 84896 6944
rect 74080 6928 74132 6934
rect 74080 6870 74132 6876
rect 74092 5778 74120 6870
rect 80520 6860 80572 6866
rect 80520 6802 80572 6808
rect 82912 6860 82964 6866
rect 82912 6802 82964 6808
rect 80244 6656 80296 6662
rect 80244 6598 80296 6604
rect 80336 6656 80388 6662
rect 80336 6598 80388 6604
rect 75552 6452 75604 6458
rect 75552 6394 75604 6400
rect 75092 6384 75144 6390
rect 75092 6326 75144 6332
rect 75104 5914 75132 6326
rect 75092 5908 75144 5914
rect 75092 5850 75144 5856
rect 74080 5772 74132 5778
rect 74080 5714 74132 5720
rect 74632 5772 74684 5778
rect 74632 5714 74684 5720
rect 73896 4820 73948 4826
rect 73896 4762 73948 4768
rect 73896 4072 73948 4078
rect 73896 4014 73948 4020
rect 74264 4072 74316 4078
rect 74264 4014 74316 4020
rect 73712 2576 73764 2582
rect 73712 2518 73764 2524
rect 73804 2576 73856 2582
rect 73804 2518 73856 2524
rect 73908 800 73936 4014
rect 74276 800 74304 4014
rect 74540 3188 74592 3194
rect 74540 3130 74592 3136
rect 74552 2038 74580 3130
rect 74644 2961 74672 5714
rect 75184 5568 75236 5574
rect 75184 5510 75236 5516
rect 75000 4684 75052 4690
rect 75000 4626 75052 4632
rect 74724 4480 74776 4486
rect 74724 4422 74776 4428
rect 74736 3466 74764 4422
rect 74724 3460 74776 3466
rect 74724 3402 74776 3408
rect 74908 3052 74960 3058
rect 74908 2994 74960 3000
rect 74630 2952 74686 2961
rect 74630 2887 74686 2896
rect 74920 2417 74948 2994
rect 74906 2408 74962 2417
rect 74906 2343 74962 2352
rect 74540 2032 74592 2038
rect 74540 1974 74592 1980
rect 74632 1420 74684 1426
rect 74632 1362 74684 1368
rect 74644 800 74672 1362
rect 75012 800 75040 4626
rect 75092 3936 75144 3942
rect 75092 3878 75144 3884
rect 75104 3505 75132 3878
rect 75090 3496 75146 3505
rect 75090 3431 75146 3440
rect 75092 3392 75144 3398
rect 75092 3334 75144 3340
rect 75104 3194 75132 3334
rect 75092 3188 75144 3194
rect 75092 3130 75144 3136
rect 75196 2582 75224 5510
rect 75368 4684 75420 4690
rect 75368 4626 75420 4632
rect 75274 4584 75330 4593
rect 75274 4519 75330 4528
rect 75288 3738 75316 4519
rect 75276 3732 75328 3738
rect 75276 3674 75328 3680
rect 75276 3392 75328 3398
rect 75276 3334 75328 3340
rect 75184 2576 75236 2582
rect 75184 2518 75236 2524
rect 75288 1018 75316 3334
rect 75276 1012 75328 1018
rect 75276 954 75328 960
rect 75380 800 75408 4626
rect 75460 4548 75512 4554
rect 75460 4490 75512 4496
rect 75472 2922 75500 4490
rect 75564 3097 75592 6394
rect 79140 6316 79192 6322
rect 79140 6258 79192 6264
rect 77208 6248 77260 6254
rect 77208 6190 77260 6196
rect 78312 6248 78364 6254
rect 78312 6190 78364 6196
rect 76564 5364 76616 5370
rect 76564 5306 76616 5312
rect 76104 5160 76156 5166
rect 76104 5102 76156 5108
rect 76472 5160 76524 5166
rect 76472 5102 76524 5108
rect 75920 5024 75972 5030
rect 75920 4966 75972 4972
rect 75932 4690 75960 4966
rect 75920 4684 75972 4690
rect 75920 4626 75972 4632
rect 75644 4480 75696 4486
rect 75644 4422 75696 4428
rect 75550 3088 75606 3097
rect 75550 3023 75606 3032
rect 75460 2916 75512 2922
rect 75460 2858 75512 2864
rect 75552 2848 75604 2854
rect 75656 2825 75684 4422
rect 75828 3732 75880 3738
rect 75828 3674 75880 3680
rect 75840 3641 75868 3674
rect 75826 3632 75882 3641
rect 75736 3596 75788 3602
rect 75826 3567 75882 3576
rect 76012 3596 76064 3602
rect 75736 3538 75788 3544
rect 76012 3538 76064 3544
rect 75552 2790 75604 2796
rect 75642 2816 75698 2825
rect 75564 1086 75592 2790
rect 75642 2751 75698 2760
rect 75748 2774 75776 3538
rect 75828 3528 75880 3534
rect 75826 3496 75828 3505
rect 75880 3496 75882 3505
rect 76024 3482 76052 3538
rect 75826 3431 75882 3440
rect 75932 3454 76052 3482
rect 75932 3126 75960 3454
rect 75920 3120 75972 3126
rect 75920 3062 75972 3068
rect 75748 2746 75868 2774
rect 75840 2514 75868 2746
rect 75828 2508 75880 2514
rect 75828 2450 75880 2456
rect 75736 1488 75788 1494
rect 75736 1430 75788 1436
rect 75552 1080 75604 1086
rect 75552 1022 75604 1028
rect 75748 800 75776 1430
rect 76116 800 76144 5102
rect 76380 5024 76432 5030
rect 76380 4966 76432 4972
rect 76288 3664 76340 3670
rect 76286 3632 76288 3641
rect 76340 3632 76342 3641
rect 76286 3567 76342 3576
rect 76288 3392 76340 3398
rect 76288 3334 76340 3340
rect 76300 3194 76328 3334
rect 76288 3188 76340 3194
rect 76288 3130 76340 3136
rect 76300 2378 76328 3130
rect 76288 2372 76340 2378
rect 76288 2314 76340 2320
rect 76392 1902 76420 4966
rect 76380 1896 76432 1902
rect 76380 1838 76432 1844
rect 76484 800 76512 5102
rect 76576 3194 76604 5306
rect 76656 4684 76708 4690
rect 76656 4626 76708 4632
rect 76668 3398 76696 4626
rect 76748 4480 76800 4486
rect 76748 4422 76800 4428
rect 76760 4078 76788 4422
rect 76748 4072 76800 4078
rect 76748 4014 76800 4020
rect 76840 3936 76892 3942
rect 76840 3878 76892 3884
rect 76748 3664 76800 3670
rect 76748 3606 76800 3612
rect 76656 3392 76708 3398
rect 76656 3334 76708 3340
rect 76564 3188 76616 3194
rect 76564 3130 76616 3136
rect 76760 3126 76788 3606
rect 76748 3120 76800 3126
rect 76654 3088 76710 3097
rect 76748 3062 76800 3068
rect 76654 3023 76710 3032
rect 76668 2922 76696 3023
rect 76656 2916 76708 2922
rect 76656 2858 76708 2864
rect 76852 800 76880 3878
rect 77116 2576 77168 2582
rect 77116 2518 77168 2524
rect 77024 2372 77076 2378
rect 77024 2314 77076 2320
rect 76932 2304 76984 2310
rect 76932 2246 76984 2252
rect 76944 1426 76972 2246
rect 77036 1494 77064 2314
rect 77128 2106 77156 2518
rect 77116 2100 77168 2106
rect 77116 2042 77168 2048
rect 77024 1488 77076 1494
rect 77024 1430 77076 1436
rect 76932 1420 76984 1426
rect 76932 1362 76984 1368
rect 77220 800 77248 6190
rect 77392 6112 77444 6118
rect 77392 6054 77444 6060
rect 77404 3369 77432 6054
rect 77760 5908 77812 5914
rect 77588 5868 77760 5896
rect 77588 5778 77616 5868
rect 77760 5850 77812 5856
rect 77576 5772 77628 5778
rect 77576 5714 77628 5720
rect 77668 5772 77720 5778
rect 77668 5714 77720 5720
rect 77576 5160 77628 5166
rect 77576 5102 77628 5108
rect 77588 4758 77616 5102
rect 77576 4752 77628 4758
rect 77576 4694 77628 4700
rect 77576 4140 77628 4146
rect 77576 4082 77628 4088
rect 77588 3942 77616 4082
rect 77576 3936 77628 3942
rect 77576 3878 77628 3884
rect 77390 3360 77446 3369
rect 77390 3295 77446 3304
rect 77576 2984 77628 2990
rect 77576 2926 77628 2932
rect 77588 2582 77616 2926
rect 77576 2576 77628 2582
rect 77576 2518 77628 2524
rect 77680 1306 77708 5714
rect 78220 5228 78272 5234
rect 78220 5170 78272 5176
rect 78128 5160 78180 5166
rect 78128 5102 78180 5108
rect 77944 4480 77996 4486
rect 77944 4422 77996 4428
rect 77850 3904 77906 3913
rect 77850 3839 77906 3848
rect 77864 3398 77892 3839
rect 77852 3392 77904 3398
rect 77758 3360 77814 3369
rect 77852 3334 77904 3340
rect 77758 3295 77814 3304
rect 77772 2650 77800 3295
rect 77864 3194 77892 3334
rect 77852 3188 77904 3194
rect 77852 3130 77904 3136
rect 77760 2644 77812 2650
rect 77760 2586 77812 2592
rect 77588 1278 77708 1306
rect 77588 800 77616 1278
rect 77956 800 77984 4422
rect 78036 4276 78088 4282
rect 78036 4218 78088 4224
rect 78048 3176 78076 4218
rect 78140 4078 78168 5102
rect 78128 4072 78180 4078
rect 78128 4014 78180 4020
rect 78232 4010 78260 5170
rect 78220 4004 78272 4010
rect 78220 3946 78272 3952
rect 78232 3602 78260 3946
rect 78220 3596 78272 3602
rect 78220 3538 78272 3544
rect 78128 3188 78180 3194
rect 78048 3148 78128 3176
rect 78128 3130 78180 3136
rect 78324 800 78352 6190
rect 78588 6112 78640 6118
rect 78588 6054 78640 6060
rect 78402 4448 78458 4457
rect 78402 4383 78458 4392
rect 78416 4282 78444 4383
rect 78404 4276 78456 4282
rect 78404 4218 78456 4224
rect 78496 4276 78548 4282
rect 78496 4218 78548 4224
rect 78508 4146 78536 4218
rect 78496 4140 78548 4146
rect 78496 4082 78548 4088
rect 78600 3233 78628 6054
rect 78680 5772 78732 5778
rect 78680 5714 78732 5720
rect 78586 3224 78642 3233
rect 78586 3159 78642 3168
rect 78600 2106 78628 3159
rect 78588 2100 78640 2106
rect 78588 2042 78640 2048
rect 78692 800 78720 5714
rect 79152 5710 79180 6258
rect 80060 6248 80112 6254
rect 80060 6190 80112 6196
rect 79876 5840 79928 5846
rect 79428 5778 79640 5794
rect 79876 5782 79928 5788
rect 79416 5772 79652 5778
rect 79468 5766 79600 5772
rect 79416 5714 79468 5720
rect 79600 5714 79652 5720
rect 79784 5772 79836 5778
rect 79784 5714 79836 5720
rect 79140 5704 79192 5710
rect 79046 5672 79102 5681
rect 79140 5646 79192 5652
rect 79428 5642 79640 5658
rect 79046 5607 79102 5616
rect 79416 5636 79652 5642
rect 78862 5400 78918 5409
rect 78772 5364 78824 5370
rect 78862 5335 78918 5344
rect 78772 5306 78824 5312
rect 78784 5234 78812 5306
rect 78772 5228 78824 5234
rect 78772 5170 78824 5176
rect 78876 3466 78904 5335
rect 79060 3738 79088 5607
rect 79468 5630 79600 5636
rect 79416 5578 79468 5584
rect 79600 5578 79652 5584
rect 79324 5024 79376 5030
rect 79324 4966 79376 4972
rect 79232 4752 79284 4758
rect 79232 4694 79284 4700
rect 79140 4004 79192 4010
rect 79140 3946 79192 3952
rect 79048 3732 79100 3738
rect 79048 3674 79100 3680
rect 78864 3460 78916 3466
rect 78864 3402 78916 3408
rect 79048 3460 79100 3466
rect 79048 3402 79100 3408
rect 79060 3369 79088 3402
rect 79046 3360 79102 3369
rect 79046 3295 79102 3304
rect 78770 3224 78826 3233
rect 78770 3159 78826 3168
rect 78784 2922 78812 3159
rect 78864 3052 78916 3058
rect 78864 2994 78916 3000
rect 78772 2916 78824 2922
rect 78772 2858 78824 2864
rect 78876 2689 78904 2994
rect 78956 2984 79008 2990
rect 78956 2926 79008 2932
rect 79046 2952 79102 2961
rect 78862 2680 78918 2689
rect 78862 2615 78918 2624
rect 78968 2281 78996 2926
rect 79046 2887 79048 2896
rect 79100 2887 79102 2896
rect 79048 2858 79100 2864
rect 79152 2774 79180 3946
rect 79244 3466 79272 4694
rect 79336 3482 79364 4966
rect 79690 4312 79746 4321
rect 79690 4247 79746 4256
rect 79414 4176 79470 4185
rect 79414 4111 79470 4120
rect 79428 3738 79456 4111
rect 79600 3936 79652 3942
rect 79600 3878 79652 3884
rect 79416 3732 79468 3738
rect 79416 3674 79468 3680
rect 79232 3460 79284 3466
rect 79336 3454 79456 3482
rect 79232 3402 79284 3408
rect 79324 3392 79376 3398
rect 79324 3334 79376 3340
rect 79336 3194 79364 3334
rect 79324 3188 79376 3194
rect 79324 3130 79376 3136
rect 79428 2972 79456 3454
rect 79336 2944 79456 2972
rect 79336 2854 79364 2944
rect 79324 2848 79376 2854
rect 79324 2790 79376 2796
rect 79612 2774 79640 3878
rect 79704 3777 79732 4247
rect 79690 3768 79746 3777
rect 79690 3703 79746 3712
rect 79692 2848 79744 2854
rect 79060 2746 79180 2774
rect 79428 2746 79640 2774
rect 79690 2816 79692 2825
rect 79744 2816 79746 2825
rect 79690 2751 79746 2760
rect 78954 2272 79010 2281
rect 78954 2207 79010 2216
rect 79060 800 79088 2746
rect 79428 800 79456 2746
rect 79796 800 79824 5714
rect 79888 3505 79916 5782
rect 79968 5568 80020 5574
rect 79968 5510 80020 5516
rect 79980 4078 80008 5510
rect 79968 4072 80020 4078
rect 79968 4014 80020 4020
rect 80072 3942 80100 6190
rect 80256 5642 80284 6598
rect 80244 5636 80296 5642
rect 80244 5578 80296 5584
rect 80244 5160 80296 5166
rect 80348 5137 80376 6598
rect 80428 6112 80480 6118
rect 80428 6054 80480 6060
rect 80244 5102 80296 5108
rect 80334 5128 80390 5137
rect 80256 4758 80284 5102
rect 80334 5063 80390 5072
rect 80336 5024 80388 5030
rect 80336 4966 80388 4972
rect 80244 4752 80296 4758
rect 80244 4694 80296 4700
rect 80152 4480 80204 4486
rect 80152 4422 80204 4428
rect 80060 3936 80112 3942
rect 80060 3878 80112 3884
rect 80060 3732 80112 3738
rect 80060 3674 80112 3680
rect 80072 3602 80100 3674
rect 80060 3596 80112 3602
rect 80060 3538 80112 3544
rect 79874 3496 79930 3505
rect 79874 3431 79930 3440
rect 80060 2984 80112 2990
rect 80060 2926 80112 2932
rect 80072 1766 80100 2926
rect 80060 1760 80112 1766
rect 80060 1702 80112 1708
rect 80164 800 80192 4422
rect 80244 4140 80296 4146
rect 80244 4082 80296 4088
rect 80256 2514 80284 4082
rect 80348 4060 80376 4966
rect 80440 4321 80468 6054
rect 80426 4312 80482 4321
rect 80426 4247 80482 4256
rect 80440 4214 80468 4247
rect 80428 4208 80480 4214
rect 80428 4150 80480 4156
rect 80428 4072 80480 4078
rect 80348 4032 80428 4060
rect 80428 4014 80480 4020
rect 80336 3936 80388 3942
rect 80336 3878 80388 3884
rect 80348 2990 80376 3878
rect 80428 3664 80480 3670
rect 80428 3606 80480 3612
rect 80336 2984 80388 2990
rect 80336 2926 80388 2932
rect 80348 2666 80376 2926
rect 80440 2854 80468 3606
rect 80428 2848 80480 2854
rect 80428 2790 80480 2796
rect 80348 2638 80468 2666
rect 80244 2508 80296 2514
rect 80244 2450 80296 2456
rect 80244 2304 80296 2310
rect 80244 2246 80296 2252
rect 80336 2304 80388 2310
rect 80336 2246 80388 2252
rect 80256 1834 80284 2246
rect 80348 2038 80376 2246
rect 80440 2145 80468 2638
rect 80426 2136 80482 2145
rect 80426 2071 80482 2080
rect 80336 2032 80388 2038
rect 80336 1974 80388 1980
rect 80244 1828 80296 1834
rect 80244 1770 80296 1776
rect 80532 800 80560 6802
rect 80612 6384 80664 6390
rect 80612 6326 80664 6332
rect 80624 3738 80652 6326
rect 80796 6248 80848 6254
rect 80796 6190 80848 6196
rect 81624 6248 81676 6254
rect 81624 6190 81676 6196
rect 81992 6248 82044 6254
rect 81992 6190 82044 6196
rect 80704 5228 80756 5234
rect 80704 5170 80756 5176
rect 80716 4554 80744 5170
rect 80704 4548 80756 4554
rect 80704 4490 80756 4496
rect 80704 4072 80756 4078
rect 80704 4014 80756 4020
rect 80612 3732 80664 3738
rect 80612 3674 80664 3680
rect 80610 3496 80666 3505
rect 80610 3431 80612 3440
rect 80664 3431 80666 3440
rect 80612 3402 80664 3408
rect 80716 3126 80744 4014
rect 80704 3120 80756 3126
rect 80704 3062 80756 3068
rect 80716 2990 80744 3062
rect 80704 2984 80756 2990
rect 80704 2926 80756 2932
rect 80612 2576 80664 2582
rect 80612 2518 80664 2524
rect 80624 1766 80652 2518
rect 80612 1760 80664 1766
rect 80612 1702 80664 1708
rect 80808 1442 80836 6190
rect 81020 6012 81316 6032
rect 81076 6010 81100 6012
rect 81156 6010 81180 6012
rect 81236 6010 81260 6012
rect 81098 5958 81100 6010
rect 81162 5958 81174 6010
rect 81236 5958 81238 6010
rect 81076 5956 81100 5958
rect 81156 5956 81180 5958
rect 81236 5956 81260 5958
rect 81020 5936 81316 5956
rect 80888 5568 80940 5574
rect 80888 5510 80940 5516
rect 80900 4758 80928 5510
rect 81532 5024 81584 5030
rect 81532 4966 81584 4972
rect 81020 4924 81316 4944
rect 81076 4922 81100 4924
rect 81156 4922 81180 4924
rect 81236 4922 81260 4924
rect 81098 4870 81100 4922
rect 81162 4870 81174 4922
rect 81236 4870 81238 4922
rect 81076 4868 81100 4870
rect 81156 4868 81180 4870
rect 81236 4868 81260 4870
rect 81020 4848 81316 4868
rect 81440 4820 81492 4826
rect 81440 4762 81492 4768
rect 80888 4752 80940 4758
rect 80888 4694 80940 4700
rect 81348 4548 81400 4554
rect 81348 4490 81400 4496
rect 80888 4480 80940 4486
rect 80888 4422 80940 4428
rect 80900 4282 80928 4422
rect 80888 4276 80940 4282
rect 80888 4218 80940 4224
rect 80888 4004 80940 4010
rect 80888 3946 80940 3952
rect 80900 3720 80928 3946
rect 81020 3836 81316 3856
rect 81076 3834 81100 3836
rect 81156 3834 81180 3836
rect 81236 3834 81260 3836
rect 81098 3782 81100 3834
rect 81162 3782 81174 3834
rect 81236 3782 81238 3834
rect 81076 3780 81100 3782
rect 81156 3780 81180 3782
rect 81236 3780 81260 3782
rect 81020 3760 81316 3780
rect 80900 3692 81020 3720
rect 80992 3602 81020 3692
rect 80980 3596 81032 3602
rect 80980 3538 81032 3544
rect 80888 3528 80940 3534
rect 80888 3470 80940 3476
rect 81070 3496 81126 3505
rect 80900 3126 80928 3470
rect 81070 3431 81126 3440
rect 81084 3398 81112 3431
rect 81072 3392 81124 3398
rect 81072 3334 81124 3340
rect 81164 3392 81216 3398
rect 81164 3334 81216 3340
rect 81176 3194 81204 3334
rect 81164 3188 81216 3194
rect 81164 3130 81216 3136
rect 80888 3120 80940 3126
rect 80888 3062 80940 3068
rect 80888 2984 80940 2990
rect 80888 2926 80940 2932
rect 80900 2825 80928 2926
rect 80886 2816 80942 2825
rect 80886 2751 80942 2760
rect 81020 2748 81316 2768
rect 81076 2746 81100 2748
rect 81156 2746 81180 2748
rect 81236 2746 81260 2748
rect 81098 2694 81100 2746
rect 81162 2694 81174 2746
rect 81236 2694 81238 2746
rect 81076 2692 81100 2694
rect 81156 2692 81180 2694
rect 81236 2692 81260 2694
rect 81020 2672 81316 2692
rect 81360 2258 81388 4490
rect 81452 3738 81480 4762
rect 81440 3732 81492 3738
rect 81440 3674 81492 3680
rect 81544 3602 81572 4966
rect 81532 3596 81584 3602
rect 81532 3538 81584 3544
rect 81544 3466 81572 3538
rect 81440 3460 81492 3466
rect 81440 3402 81492 3408
rect 81532 3460 81584 3466
rect 81532 3402 81584 3408
rect 81268 2230 81388 2258
rect 80808 1414 80928 1442
rect 80900 800 80928 1414
rect 81268 800 81296 2230
rect 81452 1562 81480 3402
rect 81532 3120 81584 3126
rect 81532 3062 81584 3068
rect 81544 2990 81572 3062
rect 81532 2984 81584 2990
rect 81532 2926 81584 2932
rect 81440 1556 81492 1562
rect 81440 1498 81492 1504
rect 81636 800 81664 6190
rect 81716 5772 81768 5778
rect 81716 5714 81768 5720
rect 81728 4865 81756 5714
rect 81808 5364 81860 5370
rect 81808 5306 81860 5312
rect 81820 5273 81848 5306
rect 81806 5264 81862 5273
rect 81806 5199 81862 5208
rect 81714 4856 81770 4865
rect 81714 4791 81770 4800
rect 81728 4486 81756 4791
rect 81716 4480 81768 4486
rect 81716 4422 81768 4428
rect 81900 4140 81952 4146
rect 81900 4082 81952 4088
rect 81808 4004 81860 4010
rect 81808 3946 81860 3952
rect 81716 3936 81768 3942
rect 81716 3878 81768 3884
rect 81728 2689 81756 3878
rect 81820 3738 81848 3946
rect 81912 3942 81940 4082
rect 81900 3936 81952 3942
rect 81900 3878 81952 3884
rect 81808 3732 81860 3738
rect 81808 3674 81860 3680
rect 81808 3596 81860 3602
rect 81808 3538 81860 3544
rect 81820 3194 81848 3538
rect 81900 3528 81952 3534
rect 81900 3470 81952 3476
rect 81808 3188 81860 3194
rect 81808 3130 81860 3136
rect 81714 2680 81770 2689
rect 81912 2650 81940 3470
rect 81714 2615 81770 2624
rect 81900 2644 81952 2650
rect 81900 2586 81952 2592
rect 81808 2576 81860 2582
rect 81808 2518 81860 2524
rect 81820 2446 81848 2518
rect 81808 2440 81860 2446
rect 81808 2382 81860 2388
rect 82004 800 82032 6190
rect 82084 6112 82136 6118
rect 82084 6054 82136 6060
rect 82820 6112 82872 6118
rect 82820 6054 82872 6060
rect 82096 3058 82124 6054
rect 82832 5914 82860 6054
rect 82820 5908 82872 5914
rect 82820 5850 82872 5856
rect 82542 5808 82598 5817
rect 82542 5743 82598 5752
rect 82820 5772 82872 5778
rect 82176 5636 82228 5642
rect 82176 5578 82228 5584
rect 82188 3670 82216 5578
rect 82452 5568 82504 5574
rect 82452 5510 82504 5516
rect 82464 5370 82492 5510
rect 82452 5364 82504 5370
rect 82452 5306 82504 5312
rect 82266 5128 82322 5137
rect 82266 5063 82268 5072
rect 82320 5063 82322 5072
rect 82268 5034 82320 5040
rect 82268 4480 82320 4486
rect 82268 4422 82320 4428
rect 82176 3664 82228 3670
rect 82176 3606 82228 3612
rect 82084 3052 82136 3058
rect 82084 2994 82136 3000
rect 82280 2990 82308 4422
rect 82464 4282 82492 5306
rect 82556 4622 82584 5743
rect 82820 5714 82872 5720
rect 82636 5228 82688 5234
rect 82636 5170 82688 5176
rect 82544 4616 82596 4622
rect 82544 4558 82596 4564
rect 82452 4276 82504 4282
rect 82452 4218 82504 4224
rect 82360 4208 82412 4214
rect 82360 4150 82412 4156
rect 82372 3670 82400 4150
rect 82360 3664 82412 3670
rect 82360 3606 82412 3612
rect 82360 3052 82412 3058
rect 82360 2994 82412 3000
rect 82176 2984 82228 2990
rect 82176 2926 82228 2932
rect 82268 2984 82320 2990
rect 82268 2926 82320 2932
rect 82188 2854 82216 2926
rect 82084 2848 82136 2854
rect 82084 2790 82136 2796
rect 82176 2848 82228 2854
rect 82176 2790 82228 2796
rect 82096 1562 82124 2790
rect 82176 2508 82228 2514
rect 82176 2450 82228 2456
rect 82268 2508 82320 2514
rect 82268 2450 82320 2456
rect 82188 1834 82216 2450
rect 82280 2106 82308 2450
rect 82268 2100 82320 2106
rect 82268 2042 82320 2048
rect 82176 1828 82228 1834
rect 82176 1770 82228 1776
rect 82084 1556 82136 1562
rect 82084 1498 82136 1504
rect 82372 800 82400 2994
rect 82464 2310 82492 4218
rect 82544 3460 82596 3466
rect 82544 3402 82596 3408
rect 82556 2990 82584 3402
rect 82544 2984 82596 2990
rect 82544 2926 82596 2932
rect 82556 2514 82584 2926
rect 82648 2854 82676 5170
rect 82832 5166 82860 5714
rect 82820 5160 82872 5166
rect 82820 5102 82872 5108
rect 82820 4684 82872 4690
rect 82820 4626 82872 4632
rect 82832 4010 82860 4626
rect 82820 4004 82872 4010
rect 82820 3946 82872 3952
rect 82818 3904 82874 3913
rect 82818 3839 82874 3848
rect 82728 3120 82780 3126
rect 82728 3062 82780 3068
rect 82740 2922 82768 3062
rect 82832 2990 82860 3839
rect 82820 2984 82872 2990
rect 82820 2926 82872 2932
rect 82728 2916 82780 2922
rect 82728 2858 82780 2864
rect 82636 2848 82688 2854
rect 82636 2790 82688 2796
rect 82924 2774 82952 6802
rect 83188 6656 83240 6662
rect 83188 6598 83240 6604
rect 83096 6248 83148 6254
rect 83096 6190 83148 6196
rect 83004 4616 83056 4622
rect 83004 4558 83056 4564
rect 83016 4457 83044 4558
rect 83002 4448 83058 4457
rect 83002 4383 83058 4392
rect 83004 4140 83056 4146
rect 83004 4082 83056 4088
rect 83016 2922 83044 4082
rect 83004 2916 83056 2922
rect 83004 2858 83056 2864
rect 82740 2746 82952 2774
rect 82544 2508 82596 2514
rect 82544 2450 82596 2456
rect 82636 2440 82688 2446
rect 82636 2382 82688 2388
rect 82648 2310 82676 2382
rect 82452 2304 82504 2310
rect 82452 2246 82504 2252
rect 82636 2304 82688 2310
rect 82636 2246 82688 2252
rect 82740 800 82768 2746
rect 82820 2508 82872 2514
rect 82820 2450 82872 2456
rect 82832 2106 82860 2450
rect 83016 2378 83044 2858
rect 83004 2372 83056 2378
rect 83004 2314 83056 2320
rect 82820 2100 82872 2106
rect 82820 2042 82872 2048
rect 83108 800 83136 6190
rect 83200 2417 83228 6598
rect 84856 6254 84884 6938
rect 85304 6316 85356 6322
rect 85304 6258 85356 6264
rect 83832 6248 83884 6254
rect 83832 6190 83884 6196
rect 84844 6248 84896 6254
rect 84844 6190 84896 6196
rect 83556 5568 83608 5574
rect 83370 5536 83426 5545
rect 83556 5510 83608 5516
rect 83370 5471 83426 5480
rect 83384 5166 83412 5471
rect 83372 5160 83424 5166
rect 83372 5102 83424 5108
rect 83464 5160 83516 5166
rect 83464 5102 83516 5108
rect 83280 5024 83332 5030
rect 83280 4966 83332 4972
rect 83372 5024 83424 5030
rect 83372 4966 83424 4972
rect 83292 3194 83320 4966
rect 83280 3188 83332 3194
rect 83280 3130 83332 3136
rect 83384 2650 83412 4966
rect 83476 3738 83504 5102
rect 83464 3732 83516 3738
rect 83464 3674 83516 3680
rect 83568 3534 83596 5510
rect 83738 5400 83794 5409
rect 83738 5335 83794 5344
rect 83648 5024 83700 5030
rect 83648 4966 83700 4972
rect 83660 4758 83688 4966
rect 83648 4752 83700 4758
rect 83648 4694 83700 4700
rect 83648 4616 83700 4622
rect 83648 4558 83700 4564
rect 83556 3528 83608 3534
rect 83556 3470 83608 3476
rect 83372 2644 83424 2650
rect 83372 2586 83424 2592
rect 83660 2582 83688 4558
rect 83752 4078 83780 5335
rect 83740 4072 83792 4078
rect 83740 4014 83792 4020
rect 83740 3392 83792 3398
rect 83740 3334 83792 3340
rect 83752 3126 83780 3334
rect 83740 3120 83792 3126
rect 83740 3062 83792 3068
rect 83740 2984 83792 2990
rect 83740 2926 83792 2932
rect 83752 2825 83780 2926
rect 83738 2816 83794 2825
rect 83738 2751 83794 2760
rect 83648 2576 83700 2582
rect 83648 2518 83700 2524
rect 83186 2408 83242 2417
rect 83186 2343 83242 2352
rect 83200 1834 83228 2343
rect 83188 1828 83240 1834
rect 83188 1770 83240 1776
rect 83464 1284 83516 1290
rect 83464 1226 83516 1232
rect 83476 800 83504 1226
rect 83844 800 83872 6190
rect 84016 6112 84068 6118
rect 84016 6054 84068 6060
rect 84028 5681 84056 6054
rect 84566 5808 84622 5817
rect 84476 5772 84528 5778
rect 84566 5743 84622 5752
rect 84936 5772 84988 5778
rect 84476 5714 84528 5720
rect 84014 5672 84070 5681
rect 84014 5607 84070 5616
rect 84028 4690 84056 5607
rect 84292 5024 84344 5030
rect 84292 4966 84344 4972
rect 84108 4820 84160 4826
rect 84108 4762 84160 4768
rect 83924 4684 83976 4690
rect 83924 4626 83976 4632
rect 84016 4684 84068 4690
rect 84016 4626 84068 4632
rect 83936 4570 83964 4626
rect 83936 4542 84056 4570
rect 83922 4448 83978 4457
rect 83922 4383 83978 4392
rect 83936 4282 83964 4383
rect 84028 4282 84056 4542
rect 83924 4276 83976 4282
rect 83924 4218 83976 4224
rect 84016 4276 84068 4282
rect 84016 4218 84068 4224
rect 83924 4004 83976 4010
rect 83924 3946 83976 3952
rect 83936 3194 83964 3946
rect 83924 3188 83976 3194
rect 83924 3130 83976 3136
rect 84028 3074 84056 4218
rect 84120 4214 84148 4762
rect 84198 4312 84254 4321
rect 84198 4247 84254 4256
rect 84108 4208 84160 4214
rect 84108 4150 84160 4156
rect 84212 4078 84240 4247
rect 84200 4072 84252 4078
rect 84200 4014 84252 4020
rect 84106 3768 84162 3777
rect 84106 3703 84162 3712
rect 84120 3602 84148 3703
rect 84108 3596 84160 3602
rect 84108 3538 84160 3544
rect 84304 3466 84332 4966
rect 84384 3596 84436 3602
rect 84384 3538 84436 3544
rect 84292 3460 84344 3466
rect 84292 3402 84344 3408
rect 84028 3046 84148 3074
rect 84016 2984 84068 2990
rect 84016 2926 84068 2932
rect 84028 1902 84056 2926
rect 84120 2650 84148 3046
rect 84304 2990 84332 3402
rect 84292 2984 84344 2990
rect 84292 2926 84344 2932
rect 84292 2848 84344 2854
rect 84198 2816 84254 2825
rect 84292 2790 84344 2796
rect 84198 2751 84254 2760
rect 84108 2644 84160 2650
rect 84108 2586 84160 2592
rect 84212 2038 84240 2751
rect 84304 2650 84332 2790
rect 84396 2650 84424 3538
rect 84292 2644 84344 2650
rect 84292 2586 84344 2592
rect 84384 2644 84436 2650
rect 84384 2586 84436 2592
rect 84200 2032 84252 2038
rect 84200 1974 84252 1980
rect 84016 1896 84068 1902
rect 84016 1838 84068 1844
rect 84488 1442 84516 5714
rect 84580 4214 84608 5743
rect 84936 5714 84988 5720
rect 84750 5400 84806 5409
rect 84660 5364 84712 5370
rect 84750 5335 84752 5344
rect 84660 5306 84712 5312
rect 84804 5335 84806 5344
rect 84752 5306 84804 5312
rect 84672 4486 84700 5306
rect 84842 4992 84898 5001
rect 84842 4927 84898 4936
rect 84856 4570 84884 4927
rect 84764 4542 84884 4570
rect 84660 4480 84712 4486
rect 84660 4422 84712 4428
rect 84568 4208 84620 4214
rect 84568 4150 84620 4156
rect 84568 4004 84620 4010
rect 84568 3946 84620 3952
rect 84580 3398 84608 3946
rect 84660 3528 84712 3534
rect 84660 3470 84712 3476
rect 84568 3392 84620 3398
rect 84568 3334 84620 3340
rect 84672 2990 84700 3470
rect 84660 2984 84712 2990
rect 84660 2926 84712 2932
rect 84764 2774 84792 4542
rect 84842 4312 84898 4321
rect 84842 4247 84898 4256
rect 84856 3126 84884 4247
rect 84844 3120 84896 3126
rect 84844 3062 84896 3068
rect 84764 2746 84884 2774
rect 84856 2514 84884 2746
rect 84568 2508 84620 2514
rect 84568 2450 84620 2456
rect 84844 2508 84896 2514
rect 84844 2450 84896 2456
rect 84580 2417 84608 2450
rect 84566 2408 84622 2417
rect 84566 2343 84622 2352
rect 84580 2310 84608 2343
rect 84568 2304 84620 2310
rect 84568 2246 84620 2252
rect 84212 1414 84516 1442
rect 84568 1420 84620 1426
rect 84212 800 84240 1414
rect 84568 1362 84620 1368
rect 84580 800 84608 1362
rect 84948 800 84976 5714
rect 85120 5568 85172 5574
rect 85120 5510 85172 5516
rect 85026 5264 85082 5273
rect 85026 5199 85082 5208
rect 85040 4214 85068 5199
rect 85028 4208 85080 4214
rect 85028 4150 85080 4156
rect 85028 3936 85080 3942
rect 85028 3878 85080 3884
rect 85040 3738 85068 3878
rect 85028 3732 85080 3738
rect 85028 3674 85080 3680
rect 85132 1630 85160 5510
rect 85212 4276 85264 4282
rect 85212 4218 85264 4224
rect 85224 3670 85252 4218
rect 85212 3664 85264 3670
rect 85212 3606 85264 3612
rect 85316 2922 85344 6258
rect 86040 5772 86092 5778
rect 86040 5714 86092 5720
rect 85762 5536 85818 5545
rect 85762 5471 85818 5480
rect 85580 5160 85632 5166
rect 85580 5102 85632 5108
rect 85488 4548 85540 4554
rect 85488 4490 85540 4496
rect 85396 4004 85448 4010
rect 85396 3946 85448 3952
rect 85408 3913 85436 3946
rect 85394 3904 85450 3913
rect 85394 3839 85450 3848
rect 85500 3777 85528 4490
rect 85486 3768 85542 3777
rect 85486 3703 85542 3712
rect 85488 3596 85540 3602
rect 85488 3538 85540 3544
rect 85396 3528 85448 3534
rect 85396 3470 85448 3476
rect 85304 2916 85356 2922
rect 85304 2858 85356 2864
rect 85210 2136 85266 2145
rect 85210 2071 85266 2080
rect 85224 1630 85252 2071
rect 85408 1902 85436 3470
rect 85500 2854 85528 3538
rect 85488 2848 85540 2854
rect 85488 2790 85540 2796
rect 85488 2644 85540 2650
rect 85488 2586 85540 2592
rect 85500 2514 85528 2586
rect 85488 2508 85540 2514
rect 85488 2450 85540 2456
rect 85396 1896 85448 1902
rect 85396 1838 85448 1844
rect 85592 1748 85620 5102
rect 85672 3936 85724 3942
rect 85672 3878 85724 3884
rect 85684 3602 85712 3878
rect 85776 3738 85804 5471
rect 85854 4448 85910 4457
rect 85854 4383 85910 4392
rect 85764 3732 85816 3738
rect 85764 3674 85816 3680
rect 85672 3596 85724 3602
rect 85672 3538 85724 3544
rect 85684 3505 85712 3538
rect 85670 3496 85726 3505
rect 85670 3431 85726 3440
rect 85764 3188 85816 3194
rect 85764 3130 85816 3136
rect 85776 3097 85804 3130
rect 85762 3088 85818 3097
rect 85762 3023 85818 3032
rect 85868 2990 85896 4383
rect 85856 2984 85908 2990
rect 85856 2926 85908 2932
rect 85856 2508 85908 2514
rect 85856 2450 85908 2456
rect 85868 1834 85896 2450
rect 85856 1828 85908 1834
rect 85856 1770 85908 1776
rect 85316 1720 85620 1748
rect 85120 1624 85172 1630
rect 85120 1566 85172 1572
rect 85212 1624 85264 1630
rect 85212 1566 85264 1572
rect 85316 800 85344 1720
rect 85672 1352 85724 1358
rect 85672 1294 85724 1300
rect 85684 800 85712 1294
rect 86052 800 86080 5714
rect 86224 5228 86276 5234
rect 86276 5188 86356 5216
rect 86224 5170 86276 5176
rect 86224 5024 86276 5030
rect 86224 4966 86276 4972
rect 86132 4480 86184 4486
rect 86132 4422 86184 4428
rect 86144 2650 86172 4422
rect 86236 4049 86264 4966
rect 86222 4040 86278 4049
rect 86222 3975 86278 3984
rect 86224 3936 86276 3942
rect 86222 3904 86224 3913
rect 86276 3904 86278 3913
rect 86222 3839 86278 3848
rect 86328 3040 86356 5188
rect 86500 5024 86552 5030
rect 86500 4966 86552 4972
rect 86512 4729 86540 4966
rect 86498 4720 86554 4729
rect 86498 4655 86554 4664
rect 86500 4616 86552 4622
rect 86500 4558 86552 4564
rect 86512 3602 86540 4558
rect 86604 3942 86632 7278
rect 87328 6792 87380 6798
rect 87328 6734 87380 6740
rect 86776 5160 86828 5166
rect 86776 5102 86828 5108
rect 87144 5160 87196 5166
rect 87144 5102 87196 5108
rect 86684 5092 86736 5098
rect 86684 5034 86736 5040
rect 86696 4078 86724 5034
rect 86788 4321 86816 5102
rect 86960 4480 87012 4486
rect 86960 4422 87012 4428
rect 86774 4312 86830 4321
rect 86774 4247 86830 4256
rect 86868 4276 86920 4282
rect 86868 4218 86920 4224
rect 86684 4072 86736 4078
rect 86684 4014 86736 4020
rect 86774 4040 86830 4049
rect 86774 3975 86830 3984
rect 86788 3942 86816 3975
rect 86592 3936 86644 3942
rect 86592 3878 86644 3884
rect 86776 3936 86828 3942
rect 86776 3878 86828 3884
rect 86880 3670 86908 4218
rect 86972 4078 87000 4422
rect 87052 4208 87104 4214
rect 87052 4150 87104 4156
rect 86960 4072 87012 4078
rect 86960 4014 87012 4020
rect 86868 3664 86920 3670
rect 86868 3606 86920 3612
rect 86500 3596 86552 3602
rect 86500 3538 86552 3544
rect 86512 3097 86540 3538
rect 86776 3460 86828 3466
rect 86776 3402 86828 3408
rect 86592 3392 86644 3398
rect 86592 3334 86644 3340
rect 86236 3012 86356 3040
rect 86498 3088 86554 3097
rect 86498 3023 86554 3032
rect 86132 2644 86184 2650
rect 86132 2586 86184 2592
rect 86236 2446 86264 3012
rect 86604 2990 86632 3334
rect 86788 3176 86816 3402
rect 87064 3398 87092 4150
rect 87052 3392 87104 3398
rect 87052 3334 87104 3340
rect 86788 3148 87000 3176
rect 86972 3097 87000 3148
rect 86958 3088 87014 3097
rect 86958 3023 87014 3032
rect 86592 2984 86644 2990
rect 86592 2926 86644 2932
rect 86776 2984 86828 2990
rect 86776 2926 86828 2932
rect 86500 2916 86552 2922
rect 86500 2858 86552 2864
rect 86406 2816 86462 2825
rect 86406 2751 86462 2760
rect 86224 2440 86276 2446
rect 86224 2382 86276 2388
rect 86420 800 86448 2751
rect 86512 2145 86540 2858
rect 86592 2848 86644 2854
rect 86592 2790 86644 2796
rect 86684 2848 86736 2854
rect 86788 2825 86816 2926
rect 86868 2916 86920 2922
rect 86868 2858 86920 2864
rect 86684 2790 86736 2796
rect 86774 2816 86830 2825
rect 86604 2582 86632 2790
rect 86592 2576 86644 2582
rect 86592 2518 86644 2524
rect 86696 2417 86724 2790
rect 86774 2751 86830 2760
rect 86776 2576 86828 2582
rect 86880 2564 86908 2858
rect 86828 2536 86908 2564
rect 86776 2518 86828 2524
rect 86682 2408 86738 2417
rect 86682 2343 86738 2352
rect 87064 2310 87092 3334
rect 86960 2304 87012 2310
rect 86960 2246 87012 2252
rect 87052 2304 87104 2310
rect 87052 2246 87104 2252
rect 86498 2136 86554 2145
rect 86498 2071 86554 2080
rect 86774 2000 86830 2009
rect 86774 1935 86830 1944
rect 86788 800 86816 1935
rect 86972 1698 87000 2246
rect 86960 1692 87012 1698
rect 86960 1634 87012 1640
rect 87156 800 87184 5102
rect 87340 3738 87368 6734
rect 88892 6724 88944 6730
rect 88892 6666 88944 6672
rect 88708 6180 88760 6186
rect 88708 6122 88760 6128
rect 87878 4856 87934 4865
rect 87878 4791 87934 4800
rect 88522 4856 88578 4865
rect 88522 4791 88578 4800
rect 87512 4684 87564 4690
rect 87512 4626 87564 4632
rect 87328 3732 87380 3738
rect 87328 3674 87380 3680
rect 87328 3596 87380 3602
rect 87328 3538 87380 3544
rect 87236 3120 87288 3126
rect 87234 3088 87236 3097
rect 87288 3088 87290 3097
rect 87234 3023 87290 3032
rect 87340 2825 87368 3538
rect 87326 2816 87382 2825
rect 87326 2751 87382 2760
rect 87328 2576 87380 2582
rect 87328 2518 87380 2524
rect 87236 2508 87288 2514
rect 87236 2450 87288 2456
rect 87248 1630 87276 2450
rect 87340 1834 87368 2518
rect 87420 2508 87472 2514
rect 87420 2450 87472 2456
rect 87432 2310 87460 2450
rect 87420 2304 87472 2310
rect 87420 2246 87472 2252
rect 87328 1828 87380 1834
rect 87328 1770 87380 1776
rect 87236 1624 87288 1630
rect 87236 1566 87288 1572
rect 87524 800 87552 4626
rect 87602 4448 87658 4457
rect 87602 4383 87658 4392
rect 87616 4146 87644 4383
rect 87604 4140 87656 4146
rect 87604 4082 87656 4088
rect 87788 4072 87840 4078
rect 87788 4014 87840 4020
rect 87696 3188 87748 3194
rect 87696 3130 87748 3136
rect 87708 2990 87736 3130
rect 87696 2984 87748 2990
rect 87696 2926 87748 2932
rect 87708 2854 87736 2926
rect 87696 2848 87748 2854
rect 87696 2790 87748 2796
rect 87696 2440 87748 2446
rect 87696 2382 87748 2388
rect 87708 2281 87736 2382
rect 87694 2272 87750 2281
rect 87694 2207 87750 2216
rect 87708 2038 87736 2207
rect 87696 2032 87748 2038
rect 87696 1974 87748 1980
rect 87800 1630 87828 4014
rect 87892 2530 87920 4791
rect 88340 4684 88392 4690
rect 88340 4626 88392 4632
rect 88156 4548 88208 4554
rect 88156 4490 88208 4496
rect 87970 4312 88026 4321
rect 87970 4247 88026 4256
rect 87984 3369 88012 4247
rect 88064 3460 88116 3466
rect 88064 3402 88116 3408
rect 87970 3360 88026 3369
rect 87970 3295 88026 3304
rect 87984 2990 88012 3295
rect 88076 3097 88104 3402
rect 88062 3088 88118 3097
rect 88062 3023 88118 3032
rect 87972 2984 88024 2990
rect 87972 2926 88024 2932
rect 87892 2502 88012 2530
rect 88076 2514 88104 3023
rect 88168 2990 88196 4490
rect 88352 3754 88380 4626
rect 88430 4584 88486 4593
rect 88430 4519 88432 4528
rect 88484 4519 88486 4528
rect 88432 4490 88484 4496
rect 88536 4282 88564 4791
rect 88720 4282 88748 6122
rect 88524 4276 88576 4282
rect 88524 4218 88576 4224
rect 88708 4276 88760 4282
rect 88708 4218 88760 4224
rect 88904 4060 88932 6666
rect 89812 6248 89864 6254
rect 89812 6190 89864 6196
rect 89076 5908 89128 5914
rect 89076 5850 89128 5856
rect 88984 5364 89036 5370
rect 88984 5306 89036 5312
rect 88996 4554 89024 5306
rect 88984 4548 89036 4554
rect 88984 4490 89036 4496
rect 88614 4040 88670 4049
rect 88904 4032 89024 4060
rect 88614 3975 88616 3984
rect 88668 3975 88670 3984
rect 88616 3946 88668 3952
rect 88260 3726 88380 3754
rect 88628 3862 88932 3890
rect 88156 2984 88208 2990
rect 88156 2926 88208 2932
rect 88156 2576 88208 2582
rect 88156 2518 88208 2524
rect 87880 2440 87932 2446
rect 87880 2382 87932 2388
rect 87984 2394 88012 2502
rect 88064 2508 88116 2514
rect 88064 2450 88116 2456
rect 87788 1624 87840 1630
rect 87788 1566 87840 1572
rect 87892 800 87920 2382
rect 87984 2366 88104 2394
rect 88076 2310 88104 2366
rect 87972 2304 88024 2310
rect 87972 2246 88024 2252
rect 88064 2304 88116 2310
rect 88064 2246 88116 2252
rect 87984 1970 88012 2246
rect 88168 1970 88196 2518
rect 87972 1964 88024 1970
rect 87972 1906 88024 1912
rect 88156 1964 88208 1970
rect 88156 1906 88208 1912
rect 88260 800 88288 3726
rect 88628 3641 88656 3862
rect 88706 3768 88762 3777
rect 88904 3738 88932 3862
rect 88706 3703 88708 3712
rect 88760 3703 88762 3712
rect 88892 3732 88944 3738
rect 88708 3674 88760 3680
rect 88892 3674 88944 3680
rect 88614 3632 88670 3641
rect 88614 3567 88670 3576
rect 88430 3496 88486 3505
rect 88430 3431 88486 3440
rect 88340 2984 88392 2990
rect 88340 2926 88392 2932
rect 88352 2038 88380 2926
rect 88444 2854 88472 3431
rect 88524 3392 88576 3398
rect 88524 3334 88576 3340
rect 88536 3194 88564 3334
rect 88524 3188 88576 3194
rect 88524 3130 88576 3136
rect 88432 2848 88484 2854
rect 88432 2790 88484 2796
rect 88892 2848 88944 2854
rect 88996 2836 89024 4032
rect 89088 3398 89116 5850
rect 89626 4856 89682 4865
rect 89626 4791 89682 4800
rect 89352 4684 89404 4690
rect 89352 4626 89404 4632
rect 89168 4480 89220 4486
rect 89168 4422 89220 4428
rect 89180 3602 89208 4422
rect 89168 3596 89220 3602
rect 89168 3538 89220 3544
rect 89076 3392 89128 3398
rect 89076 3334 89128 3340
rect 89168 3392 89220 3398
rect 89168 3334 89220 3340
rect 89180 2961 89208 3334
rect 89166 2952 89222 2961
rect 89166 2887 89222 2896
rect 88944 2808 89024 2836
rect 89168 2848 89220 2854
rect 88892 2790 88944 2796
rect 89168 2790 89220 2796
rect 88524 2508 88576 2514
rect 88524 2450 88576 2456
rect 88340 2032 88392 2038
rect 88340 1974 88392 1980
rect 88536 1902 88564 2450
rect 88524 1896 88576 1902
rect 88524 1838 88576 1844
rect 89180 1442 89208 2790
rect 88996 1414 89208 1442
rect 88616 1012 88668 1018
rect 88616 954 88668 960
rect 88628 800 88656 954
rect 88996 800 89024 1414
rect 89364 800 89392 4626
rect 89444 4276 89496 4282
rect 89444 4218 89496 4224
rect 89536 4276 89588 4282
rect 89536 4218 89588 4224
rect 89456 2990 89484 4218
rect 89548 3670 89576 4218
rect 89536 3664 89588 3670
rect 89536 3606 89588 3612
rect 89640 3398 89668 4791
rect 89718 4448 89774 4457
rect 89718 4383 89774 4392
rect 89732 4146 89760 4383
rect 89720 4140 89772 4146
rect 89720 4082 89772 4088
rect 89720 3664 89772 3670
rect 89720 3606 89772 3612
rect 89628 3392 89680 3398
rect 89628 3334 89680 3340
rect 89444 2984 89496 2990
rect 89444 2926 89496 2932
rect 89626 2816 89682 2825
rect 89626 2751 89682 2760
rect 89640 2038 89668 2751
rect 89628 2032 89680 2038
rect 89628 1974 89680 1980
rect 89732 800 89760 3606
rect 89824 3398 89852 6190
rect 89996 5704 90048 5710
rect 89996 5646 90048 5652
rect 89812 3392 89864 3398
rect 89812 3334 89864 3340
rect 89812 2644 89864 2650
rect 89812 2586 89864 2592
rect 89824 1290 89852 2586
rect 90008 2514 90036 5646
rect 92202 5128 92258 5137
rect 92202 5063 92258 5072
rect 90836 4270 91140 4298
rect 90836 4214 90864 4270
rect 91112 4214 91140 4270
rect 90824 4208 90876 4214
rect 91100 4208 91152 4214
rect 90824 4150 90876 4156
rect 91006 4176 91062 4185
rect 91100 4150 91152 4156
rect 91006 4111 91008 4120
rect 91060 4111 91062 4120
rect 91008 4082 91060 4088
rect 90456 4072 90508 4078
rect 90456 4014 90508 4020
rect 91560 4072 91612 4078
rect 91560 4014 91612 4020
rect 91652 4072 91704 4078
rect 91652 4014 91704 4020
rect 90180 3596 90232 3602
rect 90180 3538 90232 3544
rect 90088 2848 90140 2854
rect 90088 2790 90140 2796
rect 89996 2508 90048 2514
rect 89996 2450 90048 2456
rect 89812 1284 89864 1290
rect 89812 1226 89864 1232
rect 90100 800 90128 2790
rect 90192 1018 90220 3538
rect 90272 2508 90324 2514
rect 90272 2450 90324 2456
rect 90284 2310 90312 2450
rect 90364 2372 90416 2378
rect 90364 2314 90416 2320
rect 90272 2304 90324 2310
rect 90272 2246 90324 2252
rect 90376 2106 90404 2314
rect 90364 2100 90416 2106
rect 90364 2042 90416 2048
rect 90180 1012 90232 1018
rect 90180 954 90232 960
rect 90468 800 90496 4014
rect 90916 3596 90968 3602
rect 90916 3538 90968 3544
rect 90824 3460 90876 3466
rect 90824 3402 90876 3408
rect 90836 3233 90864 3402
rect 90822 3224 90878 3233
rect 90822 3159 90878 3168
rect 90928 2774 90956 3538
rect 90836 2746 90956 2774
rect 90640 2372 90692 2378
rect 90640 2314 90692 2320
rect 90652 1426 90680 2314
rect 90640 1420 90692 1426
rect 90640 1362 90692 1368
rect 90836 800 90864 2746
rect 91376 2372 91428 2378
rect 91376 2314 91428 2320
rect 91284 2304 91336 2310
rect 91284 2246 91336 2252
rect 91296 1358 91324 2246
rect 91284 1352 91336 1358
rect 91284 1294 91336 1300
rect 91388 1170 91416 2314
rect 91204 1142 91416 1170
rect 91204 800 91232 1142
rect 91572 800 91600 4014
rect 91664 3942 91692 4014
rect 91652 3936 91704 3942
rect 91652 3878 91704 3884
rect 91836 3936 91888 3942
rect 91836 3878 91888 3884
rect 91652 3732 91704 3738
rect 91652 3674 91704 3680
rect 91664 1494 91692 3674
rect 91848 2145 91876 3878
rect 91928 3596 91980 3602
rect 91928 3538 91980 3544
rect 91834 2136 91890 2145
rect 91834 2071 91890 2080
rect 91652 1488 91704 1494
rect 91652 1430 91704 1436
rect 91940 800 91968 3538
rect 92216 2922 92244 5063
rect 93768 4684 93820 4690
rect 93768 4626 93820 4632
rect 92388 4208 92440 4214
rect 92388 4150 92440 4156
rect 92204 2916 92256 2922
rect 92204 2858 92256 2864
rect 92400 2582 92428 4150
rect 92664 4072 92716 4078
rect 92664 4014 92716 4020
rect 93032 4072 93084 4078
rect 93032 4014 93084 4020
rect 92572 2848 92624 2854
rect 92572 2790 92624 2796
rect 92388 2576 92440 2582
rect 92388 2518 92440 2524
rect 92296 2508 92348 2514
rect 92296 2450 92348 2456
rect 92308 800 92336 2450
rect 92584 2310 92612 2790
rect 92572 2304 92624 2310
rect 92572 2246 92624 2252
rect 92676 800 92704 4014
rect 92756 2916 92808 2922
rect 92756 2858 92808 2864
rect 92768 1902 92796 2858
rect 92756 1896 92808 1902
rect 92756 1838 92808 1844
rect 93044 800 93072 4014
rect 93216 3936 93268 3942
rect 93216 3878 93268 3884
rect 93228 3369 93256 3878
rect 93308 3528 93360 3534
rect 93308 3470 93360 3476
rect 93214 3360 93270 3369
rect 93214 3295 93270 3304
rect 93320 3126 93348 3470
rect 93492 3392 93544 3398
rect 93492 3334 93544 3340
rect 93124 3120 93176 3126
rect 93124 3062 93176 3068
rect 93308 3120 93360 3126
rect 93308 3062 93360 3068
rect 93136 2582 93164 3062
rect 93216 3052 93268 3058
rect 93216 2994 93268 3000
rect 93228 2582 93256 2994
rect 93308 2984 93360 2990
rect 93308 2926 93360 2932
rect 93124 2576 93176 2582
rect 93124 2518 93176 2524
rect 93216 2576 93268 2582
rect 93216 2518 93268 2524
rect 93320 2514 93348 2926
rect 93400 2644 93452 2650
rect 93400 2586 93452 2592
rect 93308 2508 93360 2514
rect 93308 2450 93360 2456
rect 93412 800 93440 2586
rect 93504 1698 93532 3334
rect 93584 3052 93636 3058
rect 93584 2994 93636 3000
rect 93596 2281 93624 2994
rect 93582 2272 93638 2281
rect 93582 2207 93638 2216
rect 93492 1692 93544 1698
rect 93492 1634 93544 1640
rect 93780 800 93808 4626
rect 93964 3670 93992 12242
rect 96380 11996 96676 12016
rect 96436 11994 96460 11996
rect 96516 11994 96540 11996
rect 96596 11994 96620 11996
rect 96458 11942 96460 11994
rect 96522 11942 96534 11994
rect 96596 11942 96598 11994
rect 96436 11940 96460 11942
rect 96516 11940 96540 11942
rect 96596 11940 96620 11942
rect 96380 11920 96676 11940
rect 96380 10908 96676 10928
rect 96436 10906 96460 10908
rect 96516 10906 96540 10908
rect 96596 10906 96620 10908
rect 96458 10854 96460 10906
rect 96522 10854 96534 10906
rect 96596 10854 96598 10906
rect 96436 10852 96460 10854
rect 96516 10852 96540 10854
rect 96596 10852 96620 10854
rect 96380 10832 96676 10852
rect 96380 9820 96676 9840
rect 96436 9818 96460 9820
rect 96516 9818 96540 9820
rect 96596 9818 96620 9820
rect 96458 9766 96460 9818
rect 96522 9766 96534 9818
rect 96596 9766 96598 9818
rect 96436 9764 96460 9766
rect 96516 9764 96540 9766
rect 96596 9764 96620 9766
rect 96380 9744 96676 9764
rect 96380 8732 96676 8752
rect 96436 8730 96460 8732
rect 96516 8730 96540 8732
rect 96596 8730 96620 8732
rect 96458 8678 96460 8730
rect 96522 8678 96534 8730
rect 96596 8678 96598 8730
rect 96436 8676 96460 8678
rect 96516 8676 96540 8678
rect 96596 8676 96620 8678
rect 96380 8656 96676 8676
rect 96380 7644 96676 7664
rect 96436 7642 96460 7644
rect 96516 7642 96540 7644
rect 96596 7642 96620 7644
rect 96458 7590 96460 7642
rect 96522 7590 96534 7642
rect 96596 7590 96598 7642
rect 96436 7588 96460 7590
rect 96516 7588 96540 7590
rect 96596 7588 96620 7590
rect 96380 7568 96676 7588
rect 96380 6556 96676 6576
rect 96436 6554 96460 6556
rect 96516 6554 96540 6556
rect 96596 6554 96620 6556
rect 96458 6502 96460 6554
rect 96522 6502 96534 6554
rect 96596 6502 96598 6554
rect 96436 6500 96460 6502
rect 96516 6500 96540 6502
rect 96596 6500 96620 6502
rect 96380 6480 96676 6500
rect 96380 5468 96676 5488
rect 96436 5466 96460 5468
rect 96516 5466 96540 5468
rect 96596 5466 96620 5468
rect 96458 5414 96460 5466
rect 96522 5414 96534 5466
rect 96596 5414 96598 5466
rect 96436 5412 96460 5414
rect 96516 5412 96540 5414
rect 96596 5412 96620 5414
rect 96380 5392 96676 5412
rect 94412 5364 94464 5370
rect 94412 5306 94464 5312
rect 94424 4146 94452 5306
rect 98092 4752 98144 4758
rect 98092 4694 98144 4700
rect 94504 4480 94556 4486
rect 94504 4422 94556 4428
rect 94516 4214 94544 4422
rect 96380 4380 96676 4400
rect 96436 4378 96460 4380
rect 96516 4378 96540 4380
rect 96596 4378 96620 4380
rect 96458 4326 96460 4378
rect 96522 4326 96534 4378
rect 96596 4326 96598 4378
rect 96436 4324 96460 4326
rect 96516 4324 96540 4326
rect 96596 4324 96620 4326
rect 95054 4312 95110 4321
rect 96380 4304 96676 4324
rect 95054 4247 95110 4256
rect 94504 4208 94556 4214
rect 94504 4150 94556 4156
rect 94412 4140 94464 4146
rect 94412 4082 94464 4088
rect 94136 4072 94188 4078
rect 94136 4014 94188 4020
rect 94872 4072 94924 4078
rect 94872 4014 94924 4020
rect 93952 3664 94004 3670
rect 93952 3606 94004 3612
rect 94148 800 94176 4014
rect 94688 3596 94740 3602
rect 94688 3538 94740 3544
rect 94412 2984 94464 2990
rect 94412 2926 94464 2932
rect 94424 2582 94452 2926
rect 94412 2576 94464 2582
rect 94700 2553 94728 3538
rect 94412 2518 94464 2524
rect 94686 2544 94742 2553
rect 94686 2479 94742 2488
rect 94504 2372 94556 2378
rect 94504 2314 94556 2320
rect 94516 800 94544 2314
rect 94884 800 94912 4014
rect 95068 3942 95096 4247
rect 98000 4140 98052 4146
rect 98000 4082 98052 4088
rect 95976 4072 96028 4078
rect 95976 4014 96028 4020
rect 97080 4072 97132 4078
rect 97080 4014 97132 4020
rect 95056 3936 95108 3942
rect 95056 3878 95108 3884
rect 95608 3664 95660 3670
rect 95606 3632 95608 3641
rect 95660 3632 95662 3641
rect 95516 3596 95568 3602
rect 95606 3567 95662 3576
rect 95516 3538 95568 3544
rect 95148 3460 95200 3466
rect 95148 3402 95200 3408
rect 95160 2689 95188 3402
rect 95528 2774 95556 3538
rect 95252 2746 95556 2774
rect 95146 2680 95202 2689
rect 95146 2615 95202 2624
rect 95148 2508 95200 2514
rect 95148 2450 95200 2456
rect 95160 2106 95188 2450
rect 95148 2100 95200 2106
rect 95148 2042 95200 2048
rect 95252 800 95280 2746
rect 95608 2440 95660 2446
rect 95608 2382 95660 2388
rect 95620 800 95648 2382
rect 95988 800 96016 4014
rect 96252 3596 96304 3602
rect 96252 3538 96304 3544
rect 96068 2984 96120 2990
rect 96068 2926 96120 2932
rect 96080 2582 96108 2926
rect 96068 2576 96120 2582
rect 96068 2518 96120 2524
rect 96264 1170 96292 3538
rect 96380 3292 96676 3312
rect 96436 3290 96460 3292
rect 96516 3290 96540 3292
rect 96596 3290 96620 3292
rect 96458 3238 96460 3290
rect 96522 3238 96534 3290
rect 96596 3238 96598 3290
rect 96436 3236 96460 3238
rect 96516 3236 96540 3238
rect 96596 3236 96620 3238
rect 96380 3216 96676 3236
rect 96620 2984 96672 2990
rect 96620 2926 96672 2932
rect 96632 2582 96660 2926
rect 96620 2576 96672 2582
rect 96620 2518 96672 2524
rect 96712 2372 96764 2378
rect 96712 2314 96764 2320
rect 96380 2204 96676 2224
rect 96436 2202 96460 2204
rect 96516 2202 96540 2204
rect 96596 2202 96620 2204
rect 96458 2150 96460 2202
rect 96522 2150 96534 2202
rect 96596 2150 96598 2202
rect 96436 2148 96460 2150
rect 96516 2148 96540 2150
rect 96596 2148 96620 2150
rect 96380 2128 96676 2148
rect 96264 1142 96384 1170
rect 96356 800 96384 1142
rect 96724 800 96752 2314
rect 97092 800 97120 4014
rect 97264 3936 97316 3942
rect 98012 3913 98040 4082
rect 97264 3878 97316 3884
rect 97998 3904 98054 3913
rect 97276 2922 97304 3878
rect 97998 3839 98054 3848
rect 97448 3596 97500 3602
rect 97448 3538 97500 3544
rect 97264 2916 97316 2922
rect 97264 2858 97316 2864
rect 97460 800 97488 3538
rect 98104 3466 98132 4694
rect 98184 4072 98236 4078
rect 98184 4014 98236 4020
rect 99288 4072 99340 4078
rect 99288 4014 99340 4020
rect 100392 4072 100444 4078
rect 100392 4014 100444 4020
rect 98092 3460 98144 3466
rect 98092 3402 98144 3408
rect 97632 3392 97684 3398
rect 97632 3334 97684 3340
rect 97644 1562 97672 3334
rect 98000 2440 98052 2446
rect 98000 2382 98052 2388
rect 97632 1556 97684 1562
rect 97632 1498 97684 1504
rect 98012 1442 98040 2382
rect 97828 1414 98040 1442
rect 97828 800 97856 1414
rect 98196 800 98224 4014
rect 98368 3936 98420 3942
rect 98368 3878 98420 3884
rect 98380 1766 98408 3878
rect 98552 3596 98604 3602
rect 98552 3538 98604 3544
rect 98460 3052 98512 3058
rect 98460 2994 98512 3000
rect 98472 2582 98500 2994
rect 98460 2576 98512 2582
rect 98460 2518 98512 2524
rect 98368 1760 98420 1766
rect 98368 1702 98420 1708
rect 98564 800 98592 3538
rect 98828 3392 98880 3398
rect 98828 3334 98880 3340
rect 98920 3392 98972 3398
rect 98920 3334 98972 3340
rect 98736 2984 98788 2990
rect 98736 2926 98788 2932
rect 98748 2582 98776 2926
rect 98840 2854 98868 3334
rect 98932 3194 98960 3334
rect 98920 3188 98972 3194
rect 98920 3130 98972 3136
rect 98828 2848 98880 2854
rect 98828 2790 98880 2796
rect 98736 2576 98788 2582
rect 98736 2518 98788 2524
rect 98920 2372 98972 2378
rect 98920 2314 98972 2320
rect 98932 800 98960 2314
rect 99300 800 99328 4014
rect 99656 3596 99708 3602
rect 99656 3538 99708 3544
rect 99668 800 99696 3538
rect 99932 2984 99984 2990
rect 99932 2926 99984 2932
rect 99944 2582 99972 2926
rect 99932 2576 99984 2582
rect 99932 2518 99984 2524
rect 100024 2440 100076 2446
rect 100024 2382 100076 2388
rect 100036 800 100064 2382
rect 100404 800 100432 4014
rect 101036 4004 101088 4010
rect 101036 3946 101088 3952
rect 100760 3596 100812 3602
rect 100760 3538 100812 3544
rect 100484 3392 100536 3398
rect 100484 3334 100536 3340
rect 100496 3194 100524 3334
rect 100484 3188 100536 3194
rect 100484 3130 100536 3136
rect 100772 800 100800 3538
rect 101048 2825 101076 3946
rect 101324 3058 101352 14282
rect 127100 14172 127396 14192
rect 127156 14170 127180 14172
rect 127236 14170 127260 14172
rect 127316 14170 127340 14172
rect 127178 14118 127180 14170
rect 127242 14118 127254 14170
rect 127316 14118 127318 14170
rect 127156 14116 127180 14118
rect 127236 14116 127260 14118
rect 127316 14116 127340 14118
rect 127100 14096 127396 14116
rect 157820 14172 158116 14192
rect 157876 14170 157900 14172
rect 157956 14170 157980 14172
rect 158036 14170 158060 14172
rect 157898 14118 157900 14170
rect 157962 14118 157974 14170
rect 158036 14118 158038 14170
rect 157876 14116 157900 14118
rect 157956 14116 157980 14118
rect 158036 14116 158060 14118
rect 157820 14096 158116 14116
rect 111740 13628 112036 13648
rect 111796 13626 111820 13628
rect 111876 13626 111900 13628
rect 111956 13626 111980 13628
rect 111818 13574 111820 13626
rect 111882 13574 111894 13626
rect 111956 13574 111958 13626
rect 111796 13572 111820 13574
rect 111876 13572 111900 13574
rect 111956 13572 111980 13574
rect 111740 13552 112036 13572
rect 142460 13628 142756 13648
rect 142516 13626 142540 13628
rect 142596 13626 142620 13628
rect 142676 13626 142700 13628
rect 142538 13574 142540 13626
rect 142602 13574 142614 13626
rect 142676 13574 142678 13626
rect 142516 13572 142540 13574
rect 142596 13572 142620 13574
rect 142676 13572 142700 13574
rect 142460 13552 142756 13572
rect 173180 13628 173476 13648
rect 173236 13626 173260 13628
rect 173316 13626 173340 13628
rect 173396 13626 173420 13628
rect 173258 13574 173260 13626
rect 173322 13574 173334 13626
rect 173396 13574 173398 13626
rect 173236 13572 173260 13574
rect 173316 13572 173340 13574
rect 173396 13572 173420 13574
rect 173180 13552 173476 13572
rect 127100 13084 127396 13104
rect 127156 13082 127180 13084
rect 127236 13082 127260 13084
rect 127316 13082 127340 13084
rect 127178 13030 127180 13082
rect 127242 13030 127254 13082
rect 127316 13030 127318 13082
rect 127156 13028 127180 13030
rect 127236 13028 127260 13030
rect 127316 13028 127340 13030
rect 127100 13008 127396 13028
rect 157820 13084 158116 13104
rect 157876 13082 157900 13084
rect 157956 13082 157980 13084
rect 158036 13082 158060 13084
rect 157898 13030 157900 13082
rect 157962 13030 157974 13082
rect 158036 13030 158038 13082
rect 157876 13028 157900 13030
rect 157956 13028 157980 13030
rect 158036 13028 158060 13030
rect 157820 13008 158116 13028
rect 111740 12540 112036 12560
rect 111796 12538 111820 12540
rect 111876 12538 111900 12540
rect 111956 12538 111980 12540
rect 111818 12486 111820 12538
rect 111882 12486 111894 12538
rect 111956 12486 111958 12538
rect 111796 12484 111820 12486
rect 111876 12484 111900 12486
rect 111956 12484 111980 12486
rect 111740 12464 112036 12484
rect 142460 12540 142756 12560
rect 142516 12538 142540 12540
rect 142596 12538 142620 12540
rect 142676 12538 142700 12540
rect 142538 12486 142540 12538
rect 142602 12486 142614 12538
rect 142676 12486 142678 12538
rect 142516 12484 142540 12486
rect 142596 12484 142620 12486
rect 142676 12484 142700 12486
rect 142460 12464 142756 12484
rect 173180 12540 173476 12560
rect 173236 12538 173260 12540
rect 173316 12538 173340 12540
rect 173396 12538 173420 12540
rect 173258 12486 173260 12538
rect 173322 12486 173334 12538
rect 173396 12486 173398 12538
rect 173236 12484 173260 12486
rect 173316 12484 173340 12486
rect 173396 12484 173420 12486
rect 173180 12464 173476 12484
rect 127100 11996 127396 12016
rect 127156 11994 127180 11996
rect 127236 11994 127260 11996
rect 127316 11994 127340 11996
rect 127178 11942 127180 11994
rect 127242 11942 127254 11994
rect 127316 11942 127318 11994
rect 127156 11940 127180 11942
rect 127236 11940 127260 11942
rect 127316 11940 127340 11942
rect 127100 11920 127396 11940
rect 157820 11996 158116 12016
rect 157876 11994 157900 11996
rect 157956 11994 157980 11996
rect 158036 11994 158060 11996
rect 157898 11942 157900 11994
rect 157962 11942 157974 11994
rect 158036 11942 158038 11994
rect 157876 11940 157900 11942
rect 157956 11940 157980 11942
rect 158036 11940 158060 11942
rect 157820 11920 158116 11940
rect 111740 11452 112036 11472
rect 111796 11450 111820 11452
rect 111876 11450 111900 11452
rect 111956 11450 111980 11452
rect 111818 11398 111820 11450
rect 111882 11398 111894 11450
rect 111956 11398 111958 11450
rect 111796 11396 111820 11398
rect 111876 11396 111900 11398
rect 111956 11396 111980 11398
rect 111740 11376 112036 11396
rect 142460 11452 142756 11472
rect 142516 11450 142540 11452
rect 142596 11450 142620 11452
rect 142676 11450 142700 11452
rect 142538 11398 142540 11450
rect 142602 11398 142614 11450
rect 142676 11398 142678 11450
rect 142516 11396 142540 11398
rect 142596 11396 142620 11398
rect 142676 11396 142700 11398
rect 142460 11376 142756 11396
rect 173180 11452 173476 11472
rect 173236 11450 173260 11452
rect 173316 11450 173340 11452
rect 173396 11450 173420 11452
rect 173258 11398 173260 11450
rect 173322 11398 173334 11450
rect 173396 11398 173398 11450
rect 173236 11396 173260 11398
rect 173316 11396 173340 11398
rect 173396 11396 173420 11398
rect 173180 11376 173476 11396
rect 127100 10908 127396 10928
rect 127156 10906 127180 10908
rect 127236 10906 127260 10908
rect 127316 10906 127340 10908
rect 127178 10854 127180 10906
rect 127242 10854 127254 10906
rect 127316 10854 127318 10906
rect 127156 10852 127180 10854
rect 127236 10852 127260 10854
rect 127316 10852 127340 10854
rect 127100 10832 127396 10852
rect 157820 10908 158116 10928
rect 157876 10906 157900 10908
rect 157956 10906 157980 10908
rect 158036 10906 158060 10908
rect 157898 10854 157900 10906
rect 157962 10854 157974 10906
rect 158036 10854 158038 10906
rect 157876 10852 157900 10854
rect 157956 10852 157980 10854
rect 158036 10852 158060 10854
rect 157820 10832 158116 10852
rect 111740 10364 112036 10384
rect 111796 10362 111820 10364
rect 111876 10362 111900 10364
rect 111956 10362 111980 10364
rect 111818 10310 111820 10362
rect 111882 10310 111894 10362
rect 111956 10310 111958 10362
rect 111796 10308 111820 10310
rect 111876 10308 111900 10310
rect 111956 10308 111980 10310
rect 111740 10288 112036 10308
rect 142460 10364 142756 10384
rect 142516 10362 142540 10364
rect 142596 10362 142620 10364
rect 142676 10362 142700 10364
rect 142538 10310 142540 10362
rect 142602 10310 142614 10362
rect 142676 10310 142678 10362
rect 142516 10308 142540 10310
rect 142596 10308 142620 10310
rect 142676 10308 142700 10310
rect 142460 10288 142756 10308
rect 173180 10364 173476 10384
rect 173236 10362 173260 10364
rect 173316 10362 173340 10364
rect 173396 10362 173420 10364
rect 173258 10310 173260 10362
rect 173322 10310 173334 10362
rect 173396 10310 173398 10362
rect 173236 10308 173260 10310
rect 173316 10308 173340 10310
rect 173396 10308 173420 10310
rect 173180 10288 173476 10308
rect 127100 9820 127396 9840
rect 127156 9818 127180 9820
rect 127236 9818 127260 9820
rect 127316 9818 127340 9820
rect 127178 9766 127180 9818
rect 127242 9766 127254 9818
rect 127316 9766 127318 9818
rect 127156 9764 127180 9766
rect 127236 9764 127260 9766
rect 127316 9764 127340 9766
rect 127100 9744 127396 9764
rect 157820 9820 158116 9840
rect 157876 9818 157900 9820
rect 157956 9818 157980 9820
rect 158036 9818 158060 9820
rect 157898 9766 157900 9818
rect 157962 9766 157974 9818
rect 158036 9766 158038 9818
rect 157876 9764 157900 9766
rect 157956 9764 157980 9766
rect 158036 9764 158060 9766
rect 157820 9744 158116 9764
rect 111740 9276 112036 9296
rect 111796 9274 111820 9276
rect 111876 9274 111900 9276
rect 111956 9274 111980 9276
rect 111818 9222 111820 9274
rect 111882 9222 111894 9274
rect 111956 9222 111958 9274
rect 111796 9220 111820 9222
rect 111876 9220 111900 9222
rect 111956 9220 111980 9222
rect 111740 9200 112036 9220
rect 142460 9276 142756 9296
rect 142516 9274 142540 9276
rect 142596 9274 142620 9276
rect 142676 9274 142700 9276
rect 142538 9222 142540 9274
rect 142602 9222 142614 9274
rect 142676 9222 142678 9274
rect 142516 9220 142540 9222
rect 142596 9220 142620 9222
rect 142676 9220 142700 9222
rect 142460 9200 142756 9220
rect 173180 9276 173476 9296
rect 173236 9274 173260 9276
rect 173316 9274 173340 9276
rect 173396 9274 173420 9276
rect 173258 9222 173260 9274
rect 173322 9222 173334 9274
rect 173396 9222 173398 9274
rect 173236 9220 173260 9222
rect 173316 9220 173340 9222
rect 173396 9220 173420 9222
rect 173180 9200 173476 9220
rect 127100 8732 127396 8752
rect 127156 8730 127180 8732
rect 127236 8730 127260 8732
rect 127316 8730 127340 8732
rect 127178 8678 127180 8730
rect 127242 8678 127254 8730
rect 127316 8678 127318 8730
rect 127156 8676 127180 8678
rect 127236 8676 127260 8678
rect 127316 8676 127340 8678
rect 127100 8656 127396 8676
rect 157820 8732 158116 8752
rect 157876 8730 157900 8732
rect 157956 8730 157980 8732
rect 158036 8730 158060 8732
rect 157898 8678 157900 8730
rect 157962 8678 157974 8730
rect 158036 8678 158038 8730
rect 157876 8676 157900 8678
rect 157956 8676 157980 8678
rect 158036 8676 158060 8678
rect 157820 8656 158116 8676
rect 111740 8188 112036 8208
rect 111796 8186 111820 8188
rect 111876 8186 111900 8188
rect 111956 8186 111980 8188
rect 111818 8134 111820 8186
rect 111882 8134 111894 8186
rect 111956 8134 111958 8186
rect 111796 8132 111820 8134
rect 111876 8132 111900 8134
rect 111956 8132 111980 8134
rect 111740 8112 112036 8132
rect 142460 8188 142756 8208
rect 142516 8186 142540 8188
rect 142596 8186 142620 8188
rect 142676 8186 142700 8188
rect 142538 8134 142540 8186
rect 142602 8134 142614 8186
rect 142676 8134 142678 8186
rect 142516 8132 142540 8134
rect 142596 8132 142620 8134
rect 142676 8132 142700 8134
rect 142460 8112 142756 8132
rect 173180 8188 173476 8208
rect 173236 8186 173260 8188
rect 173316 8186 173340 8188
rect 173396 8186 173420 8188
rect 173258 8134 173260 8186
rect 173322 8134 173334 8186
rect 173396 8134 173398 8186
rect 173236 8132 173260 8134
rect 173316 8132 173340 8134
rect 173396 8132 173420 8134
rect 173180 8112 173476 8132
rect 127100 7644 127396 7664
rect 127156 7642 127180 7644
rect 127236 7642 127260 7644
rect 127316 7642 127340 7644
rect 127178 7590 127180 7642
rect 127242 7590 127254 7642
rect 127316 7590 127318 7642
rect 127156 7588 127180 7590
rect 127236 7588 127260 7590
rect 127316 7588 127340 7590
rect 127100 7568 127396 7588
rect 157820 7644 158116 7664
rect 157876 7642 157900 7644
rect 157956 7642 157980 7644
rect 158036 7642 158060 7644
rect 157898 7590 157900 7642
rect 157962 7590 157974 7642
rect 158036 7590 158038 7642
rect 157876 7588 157900 7590
rect 157956 7588 157980 7590
rect 158036 7588 158060 7590
rect 157820 7568 158116 7588
rect 111740 7100 112036 7120
rect 111796 7098 111820 7100
rect 111876 7098 111900 7100
rect 111956 7098 111980 7100
rect 111818 7046 111820 7098
rect 111882 7046 111894 7098
rect 111956 7046 111958 7098
rect 111796 7044 111820 7046
rect 111876 7044 111900 7046
rect 111956 7044 111980 7046
rect 111740 7024 112036 7044
rect 142460 7100 142756 7120
rect 142516 7098 142540 7100
rect 142596 7098 142620 7100
rect 142676 7098 142700 7100
rect 142538 7046 142540 7098
rect 142602 7046 142614 7098
rect 142676 7046 142678 7098
rect 142516 7044 142540 7046
rect 142596 7044 142620 7046
rect 142676 7044 142700 7046
rect 142460 7024 142756 7044
rect 173180 7100 173476 7120
rect 173236 7098 173260 7100
rect 173316 7098 173340 7100
rect 173396 7098 173420 7100
rect 173258 7046 173260 7098
rect 173322 7046 173334 7098
rect 173396 7046 173398 7098
rect 173236 7044 173260 7046
rect 173316 7044 173340 7046
rect 173396 7044 173420 7046
rect 173180 7024 173476 7044
rect 127100 6556 127396 6576
rect 127156 6554 127180 6556
rect 127236 6554 127260 6556
rect 127316 6554 127340 6556
rect 127178 6502 127180 6554
rect 127242 6502 127254 6554
rect 127316 6502 127318 6554
rect 127156 6500 127180 6502
rect 127236 6500 127260 6502
rect 127316 6500 127340 6502
rect 127100 6480 127396 6500
rect 157820 6556 158116 6576
rect 157876 6554 157900 6556
rect 157956 6554 157980 6556
rect 158036 6554 158060 6556
rect 157898 6502 157900 6554
rect 157962 6502 157974 6554
rect 158036 6502 158038 6554
rect 157876 6500 157900 6502
rect 157956 6500 157980 6502
rect 158036 6500 158060 6502
rect 157820 6480 158116 6500
rect 111740 6012 112036 6032
rect 111796 6010 111820 6012
rect 111876 6010 111900 6012
rect 111956 6010 111980 6012
rect 111818 5958 111820 6010
rect 111882 5958 111894 6010
rect 111956 5958 111958 6010
rect 111796 5956 111820 5958
rect 111876 5956 111900 5958
rect 111956 5956 111980 5958
rect 111740 5936 112036 5956
rect 142460 6012 142756 6032
rect 142516 6010 142540 6012
rect 142596 6010 142620 6012
rect 142676 6010 142700 6012
rect 142538 5958 142540 6010
rect 142602 5958 142614 6010
rect 142676 5958 142678 6010
rect 142516 5956 142540 5958
rect 142596 5956 142620 5958
rect 142676 5956 142700 5958
rect 142460 5936 142756 5956
rect 173180 6012 173476 6032
rect 173236 6010 173260 6012
rect 173316 6010 173340 6012
rect 173396 6010 173420 6012
rect 173258 5958 173260 6010
rect 173322 5958 173334 6010
rect 173396 5958 173398 6010
rect 173236 5956 173260 5958
rect 173316 5956 173340 5958
rect 173396 5956 173420 5958
rect 173180 5936 173476 5956
rect 178684 5772 178736 5778
rect 178684 5714 178736 5720
rect 127100 5468 127396 5488
rect 127156 5466 127180 5468
rect 127236 5466 127260 5468
rect 127316 5466 127340 5468
rect 127178 5414 127180 5466
rect 127242 5414 127254 5466
rect 127316 5414 127318 5466
rect 127156 5412 127180 5414
rect 127236 5412 127260 5414
rect 127316 5412 127340 5414
rect 127100 5392 127396 5412
rect 157820 5468 158116 5488
rect 157876 5466 157900 5468
rect 157956 5466 157980 5468
rect 158036 5466 158060 5468
rect 157898 5414 157900 5466
rect 157962 5414 157974 5466
rect 158036 5414 158038 5466
rect 157876 5412 157900 5414
rect 157956 5412 157980 5414
rect 158036 5412 158060 5414
rect 157820 5392 158116 5412
rect 177580 5160 177632 5166
rect 177580 5102 177632 5108
rect 102784 5024 102836 5030
rect 102784 4966 102836 4972
rect 102796 4826 102824 4966
rect 111740 4924 112036 4944
rect 111796 4922 111820 4924
rect 111876 4922 111900 4924
rect 111956 4922 111980 4924
rect 111818 4870 111820 4922
rect 111882 4870 111894 4922
rect 111956 4870 111958 4922
rect 111796 4868 111820 4870
rect 111876 4868 111900 4870
rect 111956 4868 111980 4870
rect 111740 4848 112036 4868
rect 142460 4924 142756 4944
rect 142516 4922 142540 4924
rect 142596 4922 142620 4924
rect 142676 4922 142700 4924
rect 142538 4870 142540 4922
rect 142602 4870 142614 4922
rect 142676 4870 142678 4922
rect 142516 4868 142540 4870
rect 142596 4868 142620 4870
rect 142676 4868 142700 4870
rect 142460 4848 142756 4868
rect 173180 4924 173476 4944
rect 173236 4922 173260 4924
rect 173316 4922 173340 4924
rect 173396 4922 173420 4924
rect 173258 4870 173260 4922
rect 173322 4870 173334 4922
rect 173396 4870 173398 4922
rect 173236 4868 173260 4870
rect 173316 4868 173340 4870
rect 173396 4868 173420 4870
rect 173180 4848 173476 4868
rect 102784 4820 102836 4826
rect 102784 4762 102836 4768
rect 102600 4684 102652 4690
rect 102600 4626 102652 4632
rect 175372 4684 175424 4690
rect 175372 4626 175424 4632
rect 176660 4684 176712 4690
rect 176660 4626 176712 4632
rect 101496 4072 101548 4078
rect 101496 4014 101548 4020
rect 101586 4040 101642 4049
rect 101404 3936 101456 3942
rect 101404 3878 101456 3884
rect 101416 3670 101444 3878
rect 101404 3664 101456 3670
rect 101404 3606 101456 3612
rect 101404 3528 101456 3534
rect 101404 3470 101456 3476
rect 101312 3052 101364 3058
rect 101312 2994 101364 3000
rect 101128 2984 101180 2990
rect 101416 2961 101444 3470
rect 101128 2926 101180 2932
rect 101402 2952 101458 2961
rect 101034 2816 101090 2825
rect 101034 2751 101090 2760
rect 101140 2582 101168 2926
rect 101402 2887 101458 2896
rect 101128 2576 101180 2582
rect 101128 2518 101180 2524
rect 101128 2372 101180 2378
rect 101128 2314 101180 2320
rect 101140 800 101168 2314
rect 101508 800 101536 4014
rect 101586 3975 101642 3984
rect 101600 3534 101628 3975
rect 102048 3936 102100 3942
rect 102048 3878 102100 3884
rect 101862 3768 101918 3777
rect 101680 3732 101732 3738
rect 101680 3674 101732 3680
rect 101772 3732 101824 3738
rect 101862 3703 101918 3712
rect 101772 3674 101824 3680
rect 101588 3528 101640 3534
rect 101588 3470 101640 3476
rect 101692 3194 101720 3674
rect 101784 3641 101812 3674
rect 101876 3670 101904 3703
rect 101864 3664 101916 3670
rect 101770 3632 101826 3641
rect 101864 3606 101916 3612
rect 101770 3567 101826 3576
rect 101956 3596 102008 3602
rect 101956 3538 102008 3544
rect 101864 3392 101916 3398
rect 101864 3334 101916 3340
rect 101680 3188 101732 3194
rect 101680 3130 101732 3136
rect 101876 2582 101904 3334
rect 101864 2576 101916 2582
rect 101864 2518 101916 2524
rect 101968 1816 101996 3538
rect 102060 3466 102088 3878
rect 102048 3460 102100 3466
rect 102048 3402 102100 3408
rect 102324 3460 102376 3466
rect 102324 3402 102376 3408
rect 102232 3392 102284 3398
rect 102232 3334 102284 3340
rect 102138 3088 102194 3097
rect 102138 3023 102140 3032
rect 102192 3023 102194 3032
rect 102140 2994 102192 3000
rect 102244 2582 102272 3334
rect 102336 2854 102364 3402
rect 102324 2848 102376 2854
rect 102324 2790 102376 2796
rect 102508 2848 102560 2854
rect 102508 2790 102560 2796
rect 102232 2576 102284 2582
rect 102232 2518 102284 2524
rect 102520 2514 102548 2790
rect 102508 2508 102560 2514
rect 102508 2450 102560 2456
rect 102232 2304 102284 2310
rect 102232 2246 102284 2252
rect 101876 1788 101996 1816
rect 101876 800 101904 1788
rect 102244 800 102272 2246
rect 102612 800 102640 4626
rect 127100 4380 127396 4400
rect 127156 4378 127180 4380
rect 127236 4378 127260 4380
rect 127316 4378 127340 4380
rect 127178 4326 127180 4378
rect 127242 4326 127254 4378
rect 127316 4326 127318 4378
rect 127156 4324 127180 4326
rect 127236 4324 127260 4326
rect 127316 4324 127340 4326
rect 127100 4304 127396 4324
rect 157820 4380 158116 4400
rect 157876 4378 157900 4380
rect 157956 4378 157980 4380
rect 158036 4378 158060 4380
rect 157898 4326 157900 4378
rect 157962 4326 157974 4378
rect 158036 4326 158038 4378
rect 157876 4324 157900 4326
rect 157956 4324 157980 4326
rect 158036 4324 158060 4326
rect 157820 4304 158116 4324
rect 109316 4276 109368 4282
rect 109316 4218 109368 4224
rect 102876 4140 102928 4146
rect 102876 4082 102928 4088
rect 102888 3398 102916 4082
rect 102968 4072 103020 4078
rect 102968 4014 103020 4020
rect 103796 4072 103848 4078
rect 103796 4014 103848 4020
rect 104808 4072 104860 4078
rect 104808 4014 104860 4020
rect 105912 4072 105964 4078
rect 105912 4014 105964 4020
rect 107016 4072 107068 4078
rect 107016 4014 107068 4020
rect 102876 3392 102928 3398
rect 102876 3334 102928 3340
rect 102874 2952 102930 2961
rect 102874 2887 102876 2896
rect 102928 2887 102930 2896
rect 102876 2858 102928 2864
rect 102980 800 103008 4014
rect 103520 4004 103572 4010
rect 103520 3946 103572 3952
rect 103060 3936 103112 3942
rect 103060 3878 103112 3884
rect 103072 1834 103100 3878
rect 103532 3233 103560 3946
rect 103518 3224 103574 3233
rect 103518 3159 103574 3168
rect 103704 2984 103756 2990
rect 103704 2926 103756 2932
rect 103716 2582 103744 2926
rect 103152 2576 103204 2582
rect 103152 2518 103204 2524
rect 103704 2576 103756 2582
rect 103704 2518 103756 2524
rect 103164 1970 103192 2518
rect 103336 2304 103388 2310
rect 103336 2246 103388 2252
rect 103152 1964 103204 1970
rect 103152 1906 103204 1912
rect 103060 1828 103112 1834
rect 103060 1770 103112 1776
rect 103348 800 103376 2246
rect 103808 2122 103836 4014
rect 103888 3936 103940 3942
rect 103888 3878 103940 3884
rect 103900 3126 103928 3878
rect 104072 3596 104124 3602
rect 104072 3538 104124 3544
rect 103888 3120 103940 3126
rect 103888 3062 103940 3068
rect 103716 2094 103836 2122
rect 103716 800 103744 2094
rect 104084 800 104112 3538
rect 104440 2984 104492 2990
rect 104440 2926 104492 2932
rect 104452 2582 104480 2926
rect 104440 2576 104492 2582
rect 104440 2518 104492 2524
rect 104440 2304 104492 2310
rect 104440 2246 104492 2252
rect 104452 800 104480 2246
rect 104820 800 104848 4014
rect 105176 3596 105228 3602
rect 105176 3538 105228 3544
rect 105188 800 105216 3538
rect 105544 2984 105596 2990
rect 105544 2926 105596 2932
rect 105556 2582 105584 2926
rect 105544 2576 105596 2582
rect 105544 2518 105596 2524
rect 105544 2304 105596 2310
rect 105544 2246 105596 2252
rect 105556 800 105584 2246
rect 105924 800 105952 4014
rect 106280 3596 106332 3602
rect 106280 3538 106332 3544
rect 106292 800 106320 3538
rect 106464 3392 106516 3398
rect 106464 3334 106516 3340
rect 106476 2650 106504 3334
rect 106648 2984 106700 2990
rect 106648 2926 106700 2932
rect 106464 2644 106516 2650
rect 106464 2586 106516 2592
rect 106660 2582 106688 2926
rect 106648 2576 106700 2582
rect 106648 2518 106700 2524
rect 106648 2304 106700 2310
rect 106648 2246 106700 2252
rect 106924 2304 106976 2310
rect 106924 2246 106976 2252
rect 106660 800 106688 2246
rect 106936 1698 106964 2246
rect 106924 1692 106976 1698
rect 106924 1634 106976 1640
rect 107028 800 107056 4014
rect 107292 3936 107344 3942
rect 107292 3878 107344 3884
rect 107476 3936 107528 3942
rect 107476 3878 107528 3884
rect 107200 2916 107252 2922
rect 107200 2858 107252 2864
rect 107212 2650 107240 2858
rect 107304 2854 107332 3878
rect 107384 3596 107436 3602
rect 107384 3538 107436 3544
rect 107292 2848 107344 2854
rect 107292 2790 107344 2796
rect 107200 2644 107252 2650
rect 107200 2586 107252 2592
rect 107396 800 107424 3538
rect 107488 3058 107516 3878
rect 109328 3738 109356 4218
rect 109960 4208 110012 4214
rect 109960 4150 110012 4156
rect 109972 3738 110000 4150
rect 111432 4072 111484 4078
rect 111432 4014 111484 4020
rect 112536 4072 112588 4078
rect 112536 4014 112588 4020
rect 113640 4072 113692 4078
rect 113640 4014 113692 4020
rect 114744 4072 114796 4078
rect 114744 4014 114796 4020
rect 115848 4072 115900 4078
rect 115848 4014 115900 4020
rect 116952 4072 117004 4078
rect 116952 4014 117004 4020
rect 118056 4072 118108 4078
rect 118056 4014 118108 4020
rect 119160 4072 119212 4078
rect 119160 4014 119212 4020
rect 120172 4072 120224 4078
rect 120172 4014 120224 4020
rect 121276 4072 121328 4078
rect 121276 4014 121328 4020
rect 122288 4072 122340 4078
rect 122288 4014 122340 4020
rect 123484 4072 123536 4078
rect 123484 4014 123536 4020
rect 124588 4072 124640 4078
rect 124588 4014 124640 4020
rect 125692 4072 125744 4078
rect 125692 4014 125744 4020
rect 126796 4072 126848 4078
rect 126796 4014 126848 4020
rect 127900 4072 127952 4078
rect 127900 4014 127952 4020
rect 131212 4072 131264 4078
rect 131212 4014 131264 4020
rect 133420 4072 133472 4078
rect 133420 4014 133472 4020
rect 134524 4072 134576 4078
rect 134524 4014 134576 4020
rect 136732 4072 136784 4078
rect 136732 4014 136784 4020
rect 137836 4072 137888 4078
rect 137836 4014 137888 4020
rect 138940 4072 138992 4078
rect 138940 4014 138992 4020
rect 140044 4072 140096 4078
rect 140044 4014 140096 4020
rect 141148 4072 141200 4078
rect 141148 4014 141200 4020
rect 142252 4072 142304 4078
rect 142252 4014 142304 4020
rect 143448 4072 143500 4078
rect 143448 4014 143500 4020
rect 144460 4072 144512 4078
rect 144460 4014 144512 4020
rect 145564 4072 145616 4078
rect 145564 4014 145616 4020
rect 146668 4072 146720 4078
rect 146668 4014 146720 4020
rect 147772 4072 147824 4078
rect 147772 4014 147824 4020
rect 148876 4072 148928 4078
rect 148876 4014 148928 4020
rect 152188 4072 152240 4078
rect 152188 4014 152240 4020
rect 153292 4072 153344 4078
rect 153292 4014 153344 4020
rect 154396 4072 154448 4078
rect 154396 4014 154448 4020
rect 155500 4072 155552 4078
rect 155500 4014 155552 4020
rect 157708 4072 157760 4078
rect 157708 4014 157760 4020
rect 158812 4072 158864 4078
rect 158812 4014 158864 4020
rect 159916 4072 159968 4078
rect 159916 4014 159968 4020
rect 161020 4072 161072 4078
rect 161020 4014 161072 4020
rect 162124 4072 162176 4078
rect 162124 4014 162176 4020
rect 165436 4072 165488 4078
rect 165436 4014 165488 4020
rect 166540 4072 166592 4078
rect 166540 4014 166592 4020
rect 167644 4072 167696 4078
rect 167644 4014 167696 4020
rect 168748 4072 168800 4078
rect 168748 4014 168800 4020
rect 169852 4072 169904 4078
rect 169852 4014 169904 4020
rect 173072 4072 173124 4078
rect 173072 4014 173124 4020
rect 174268 4072 174320 4078
rect 174268 4014 174320 4020
rect 109316 3732 109368 3738
rect 109316 3674 109368 3680
rect 109960 3732 110012 3738
rect 109960 3674 110012 3680
rect 108488 3596 108540 3602
rect 108488 3538 108540 3544
rect 109224 3596 109276 3602
rect 109224 3538 109276 3544
rect 110696 3596 110748 3602
rect 110696 3538 110748 3544
rect 107476 3052 107528 3058
rect 107476 2994 107528 3000
rect 108120 2508 108172 2514
rect 108120 2450 108172 2456
rect 107752 2440 107804 2446
rect 107752 2382 107804 2388
rect 107764 800 107792 2382
rect 108132 800 108160 2450
rect 108500 800 108528 3538
rect 109132 3052 109184 3058
rect 109132 2994 109184 3000
rect 109144 2582 109172 2994
rect 109132 2576 109184 2582
rect 109132 2518 109184 2524
rect 108856 2372 108908 2378
rect 108856 2314 108908 2320
rect 108868 800 108896 2314
rect 109236 800 109264 3538
rect 109868 2984 109920 2990
rect 109868 2926 109920 2932
rect 109592 2916 109644 2922
rect 109592 2858 109644 2864
rect 109604 800 109632 2858
rect 109880 2582 109908 2926
rect 109868 2576 109920 2582
rect 109868 2518 109920 2524
rect 110328 2508 110380 2514
rect 110328 2450 110380 2456
rect 109960 2440 110012 2446
rect 109960 2382 110012 2388
rect 109972 800 110000 2382
rect 110340 800 110368 2450
rect 110708 800 110736 3538
rect 111064 2372 111116 2378
rect 111064 2314 111116 2320
rect 111076 800 111104 2314
rect 111444 800 111472 4014
rect 111740 3836 112036 3856
rect 111796 3834 111820 3836
rect 111876 3834 111900 3836
rect 111956 3834 111980 3836
rect 111818 3782 111820 3834
rect 111882 3782 111894 3834
rect 111956 3782 111958 3834
rect 111796 3780 111820 3782
rect 111876 3780 111900 3782
rect 111956 3780 111980 3782
rect 111740 3760 112036 3780
rect 112076 3596 112128 3602
rect 112076 3538 112128 3544
rect 111616 3052 111668 3058
rect 111616 2994 111668 3000
rect 111628 2582 111656 2994
rect 111740 2748 112036 2768
rect 111796 2746 111820 2748
rect 111876 2746 111900 2748
rect 111956 2746 111980 2748
rect 111818 2694 111820 2746
rect 111882 2694 111894 2746
rect 111956 2694 111958 2746
rect 111796 2692 111820 2694
rect 111876 2692 111900 2694
rect 111956 2692 111980 2694
rect 111740 2672 112036 2692
rect 111616 2576 111668 2582
rect 111616 2518 111668 2524
rect 112088 1850 112116 3538
rect 112444 2984 112496 2990
rect 112444 2926 112496 2932
rect 112456 2582 112484 2926
rect 112444 2576 112496 2582
rect 112444 2518 112496 2524
rect 112168 2372 112220 2378
rect 112168 2314 112220 2320
rect 111812 1822 112116 1850
rect 111812 800 111840 1822
rect 112180 800 112208 2314
rect 112548 800 112576 4014
rect 112904 3596 112956 3602
rect 112904 3538 112956 3544
rect 112916 800 112944 3538
rect 113180 2984 113232 2990
rect 113180 2926 113232 2932
rect 113192 2582 113220 2926
rect 113180 2576 113232 2582
rect 113180 2518 113232 2524
rect 113272 2304 113324 2310
rect 113272 2246 113324 2252
rect 113284 800 113312 2246
rect 113652 800 113680 4014
rect 114008 3596 114060 3602
rect 114008 3538 114060 3544
rect 114020 800 114048 3538
rect 114284 2984 114336 2990
rect 114284 2926 114336 2932
rect 114296 2582 114324 2926
rect 114284 2576 114336 2582
rect 114284 2518 114336 2524
rect 114376 2372 114428 2378
rect 114376 2314 114428 2320
rect 114388 800 114416 2314
rect 114756 800 114784 4014
rect 115112 3596 115164 3602
rect 115112 3538 115164 3544
rect 115124 800 115152 3538
rect 115204 2984 115256 2990
rect 115204 2926 115256 2932
rect 115216 2582 115244 2926
rect 115204 2576 115256 2582
rect 115204 2518 115256 2524
rect 115480 2304 115532 2310
rect 115480 2246 115532 2252
rect 115492 800 115520 2246
rect 115860 800 115888 4014
rect 116216 3596 116268 3602
rect 116216 3538 116268 3544
rect 116228 800 116256 3538
rect 116400 2984 116452 2990
rect 116400 2926 116452 2932
rect 116412 2582 116440 2926
rect 116400 2576 116452 2582
rect 116400 2518 116452 2524
rect 116584 2372 116636 2378
rect 116584 2314 116636 2320
rect 116596 800 116624 2314
rect 116964 800 116992 4014
rect 117320 3596 117372 3602
rect 117320 3538 117372 3544
rect 117136 2984 117188 2990
rect 117136 2926 117188 2932
rect 117148 2582 117176 2926
rect 117136 2576 117188 2582
rect 117136 2518 117188 2524
rect 117332 800 117360 3538
rect 117780 2984 117832 2990
rect 117780 2926 117832 2932
rect 117792 2582 117820 2926
rect 117780 2576 117832 2582
rect 117780 2518 117832 2524
rect 117688 2304 117740 2310
rect 117688 2246 117740 2252
rect 117700 800 117728 2246
rect 118068 800 118096 4014
rect 118424 3596 118476 3602
rect 118424 3538 118476 3544
rect 118436 800 118464 3538
rect 118792 2984 118844 2990
rect 118792 2926 118844 2932
rect 118804 2582 118832 2926
rect 118792 2576 118844 2582
rect 118792 2518 118844 2524
rect 118792 2304 118844 2310
rect 118792 2246 118844 2252
rect 118804 800 118832 2246
rect 119172 800 119200 4014
rect 119528 3596 119580 3602
rect 119528 3538 119580 3544
rect 119540 800 119568 3538
rect 119896 2984 119948 2990
rect 119896 2926 119948 2932
rect 119908 2582 119936 2926
rect 119896 2576 119948 2582
rect 119896 2518 119948 2524
rect 119896 2304 119948 2310
rect 119896 2246 119948 2252
rect 119908 800 119936 2246
rect 120184 800 120212 4014
rect 120540 3596 120592 3602
rect 120540 3538 120592 3544
rect 120552 800 120580 3538
rect 120908 2304 120960 2310
rect 120908 2246 120960 2252
rect 120920 800 120948 2246
rect 121288 800 121316 4014
rect 121644 3596 121696 3602
rect 121644 3538 121696 3544
rect 121656 800 121684 3538
rect 121736 2984 121788 2990
rect 121736 2926 121788 2932
rect 121748 2582 121776 2926
rect 121736 2576 121788 2582
rect 121736 2518 121788 2524
rect 122012 2304 122064 2310
rect 122012 2246 122064 2252
rect 122024 800 122052 2246
rect 122300 1442 122328 4014
rect 122748 3596 122800 3602
rect 122748 3538 122800 3544
rect 122380 2984 122432 2990
rect 122380 2926 122432 2932
rect 122392 2582 122420 2926
rect 122380 2576 122432 2582
rect 122380 2518 122432 2524
rect 122300 1414 122420 1442
rect 122392 800 122420 1414
rect 122760 800 122788 3538
rect 123116 2984 123168 2990
rect 123116 2926 123168 2932
rect 123128 2582 123156 2926
rect 123116 2576 123168 2582
rect 123116 2518 123168 2524
rect 123116 2304 123168 2310
rect 123116 2246 123168 2252
rect 123128 800 123156 2246
rect 123496 800 123524 4014
rect 123852 3596 123904 3602
rect 123852 3538 123904 3544
rect 123864 800 123892 3538
rect 124220 2984 124272 2990
rect 124220 2926 124272 2932
rect 124232 2582 124260 2926
rect 124220 2576 124272 2582
rect 124220 2518 124272 2524
rect 124220 2304 124272 2310
rect 124220 2246 124272 2252
rect 124232 800 124260 2246
rect 124600 800 124628 4014
rect 124956 3596 125008 3602
rect 124956 3538 125008 3544
rect 124968 800 124996 3538
rect 125324 2984 125376 2990
rect 125324 2926 125376 2932
rect 125336 2582 125364 2926
rect 125324 2576 125376 2582
rect 125324 2518 125376 2524
rect 125324 2372 125376 2378
rect 125324 2314 125376 2320
rect 125336 800 125364 2314
rect 125704 800 125732 4014
rect 126060 3596 126112 3602
rect 126060 3538 126112 3544
rect 126072 800 126100 3538
rect 126428 2304 126480 2310
rect 126428 2246 126480 2252
rect 126440 800 126468 2246
rect 126808 800 126836 4014
rect 126980 3596 127032 3602
rect 126980 3538 127032 3544
rect 126992 1850 127020 3538
rect 127100 3292 127396 3312
rect 127156 3290 127180 3292
rect 127236 3290 127260 3292
rect 127316 3290 127340 3292
rect 127178 3238 127180 3290
rect 127242 3238 127254 3290
rect 127316 3238 127318 3290
rect 127156 3236 127180 3238
rect 127236 3236 127260 3238
rect 127316 3236 127340 3238
rect 127100 3216 127396 3236
rect 127072 2984 127124 2990
rect 127072 2926 127124 2932
rect 127624 2984 127676 2990
rect 127624 2926 127676 2932
rect 127084 2582 127112 2926
rect 127636 2582 127664 2926
rect 127072 2576 127124 2582
rect 127072 2518 127124 2524
rect 127624 2576 127676 2582
rect 127624 2518 127676 2524
rect 127532 2304 127584 2310
rect 127532 2246 127584 2252
rect 127100 2204 127396 2224
rect 127156 2202 127180 2204
rect 127236 2202 127260 2204
rect 127316 2202 127340 2204
rect 127178 2150 127180 2202
rect 127242 2150 127254 2202
rect 127316 2150 127318 2202
rect 127156 2148 127180 2150
rect 127236 2148 127260 2150
rect 127316 2148 127340 2150
rect 127100 2128 127396 2148
rect 126992 1822 127204 1850
rect 127176 800 127204 1822
rect 127544 800 127572 2246
rect 127912 800 127940 4014
rect 128268 3596 128320 3602
rect 128268 3538 128320 3544
rect 129004 3596 129056 3602
rect 129004 3538 129056 3544
rect 129372 3596 129424 3602
rect 130200 3596 130252 3602
rect 129372 3538 129424 3544
rect 130120 3556 130200 3584
rect 128280 800 128308 3538
rect 128636 2984 128688 2990
rect 128636 2926 128688 2932
rect 128648 2582 128676 2926
rect 128636 2576 128688 2582
rect 128636 2518 128688 2524
rect 128636 2304 128688 2310
rect 128636 2246 128688 2252
rect 128648 800 128676 2246
rect 129016 800 129044 3538
rect 129384 800 129412 3538
rect 129740 2984 129792 2990
rect 129740 2926 129792 2932
rect 129752 2582 129780 2926
rect 129740 2576 129792 2582
rect 129740 2518 129792 2524
rect 129740 2304 129792 2310
rect 129740 2246 129792 2252
rect 129752 800 129780 2246
rect 130120 800 130148 3556
rect 130200 3538 130252 3544
rect 130844 2984 130896 2990
rect 130844 2926 130896 2932
rect 130476 2916 130528 2922
rect 130476 2858 130528 2864
rect 130488 800 130516 2858
rect 130856 2582 130884 2926
rect 130844 2576 130896 2582
rect 130844 2518 130896 2524
rect 130844 2372 130896 2378
rect 130844 2314 130896 2320
rect 130856 800 130884 2314
rect 131224 800 131252 4014
rect 131580 3596 131632 3602
rect 131580 3538 131632 3544
rect 131592 800 131620 3538
rect 132316 3528 132368 3534
rect 132316 3470 132368 3476
rect 131948 3392 132000 3398
rect 131948 3334 132000 3340
rect 131960 2582 131988 3334
rect 131948 2576 132000 2582
rect 131948 2518 132000 2524
rect 131948 2304 132000 2310
rect 131948 2246 132000 2252
rect 131960 800 131988 2246
rect 132328 800 132356 3470
rect 133052 2984 133104 2990
rect 133052 2926 133104 2932
rect 133064 2582 133092 2926
rect 133052 2576 133104 2582
rect 133052 2518 133104 2524
rect 132684 2508 132736 2514
rect 132684 2450 132736 2456
rect 132696 800 132724 2450
rect 133052 2304 133104 2310
rect 133052 2246 133104 2252
rect 133064 800 133092 2246
rect 133432 800 133460 4014
rect 133788 3596 133840 3602
rect 133788 3538 133840 3544
rect 133800 800 133828 3538
rect 134156 2984 134208 2990
rect 134156 2926 134208 2932
rect 134168 2582 134196 2926
rect 134156 2576 134208 2582
rect 134156 2518 134208 2524
rect 134156 2304 134208 2310
rect 134156 2246 134208 2252
rect 134168 800 134196 2246
rect 134536 800 134564 4014
rect 134892 3596 134944 3602
rect 134892 3538 134944 3544
rect 135628 3596 135680 3602
rect 135628 3538 135680 3544
rect 134904 800 134932 3538
rect 135260 2984 135312 2990
rect 135260 2926 135312 2932
rect 135272 2582 135300 2926
rect 135260 2576 135312 2582
rect 135260 2518 135312 2524
rect 135260 2304 135312 2310
rect 135260 2246 135312 2252
rect 135272 800 135300 2246
rect 135640 800 135668 3538
rect 136364 2984 136416 2990
rect 136364 2926 136416 2932
rect 135996 2916 136048 2922
rect 135996 2858 136048 2864
rect 136008 800 136036 2858
rect 136376 2582 136404 2926
rect 136364 2576 136416 2582
rect 136364 2518 136416 2524
rect 136364 2304 136416 2310
rect 136364 2246 136416 2252
rect 136376 800 136404 2246
rect 136744 800 136772 4014
rect 137100 3596 137152 3602
rect 137100 3538 137152 3544
rect 137112 800 137140 3538
rect 137468 2304 137520 2310
rect 137468 2246 137520 2252
rect 137480 800 137508 2246
rect 137848 800 137876 4014
rect 138204 3596 138256 3602
rect 138204 3538 138256 3544
rect 138112 2984 138164 2990
rect 138112 2926 138164 2932
rect 138124 2582 138152 2926
rect 138112 2576 138164 2582
rect 138112 2518 138164 2524
rect 138216 800 138244 3538
rect 138756 2984 138808 2990
rect 138756 2926 138808 2932
rect 138768 2582 138796 2926
rect 138756 2576 138808 2582
rect 138756 2518 138808 2524
rect 138572 2304 138624 2310
rect 138572 2246 138624 2252
rect 138584 800 138612 2246
rect 138952 800 138980 4014
rect 139308 3596 139360 3602
rect 139308 3538 139360 3544
rect 139320 800 139348 3538
rect 139676 2984 139728 2990
rect 139676 2926 139728 2932
rect 139688 2582 139716 2926
rect 139676 2576 139728 2582
rect 139676 2518 139728 2524
rect 139676 2304 139728 2310
rect 139676 2246 139728 2252
rect 139688 800 139716 2246
rect 140056 800 140084 4014
rect 140412 3596 140464 3602
rect 140412 3538 140464 3544
rect 140424 800 140452 3538
rect 140780 2984 140832 2990
rect 140780 2926 140832 2932
rect 140792 2582 140820 2926
rect 140780 2576 140832 2582
rect 140780 2518 140832 2524
rect 140780 2304 140832 2310
rect 140780 2246 140832 2252
rect 140792 800 140820 2246
rect 141160 800 141188 4014
rect 141516 3596 141568 3602
rect 141516 3538 141568 3544
rect 141528 800 141556 3538
rect 141884 2984 141936 2990
rect 141884 2926 141936 2932
rect 141896 2582 141924 2926
rect 141884 2576 141936 2582
rect 141884 2518 141936 2524
rect 141884 2304 141936 2310
rect 141884 2246 141936 2252
rect 141896 800 141924 2246
rect 142264 800 142292 4014
rect 142460 3836 142756 3856
rect 142516 3834 142540 3836
rect 142596 3834 142620 3836
rect 142676 3834 142700 3836
rect 142538 3782 142540 3834
rect 142602 3782 142614 3834
rect 142676 3782 142678 3834
rect 142516 3780 142540 3782
rect 142596 3780 142620 3782
rect 142676 3780 142700 3782
rect 142460 3760 142756 3780
rect 142804 3596 142856 3602
rect 142804 3538 142856 3544
rect 142460 2748 142756 2768
rect 142516 2746 142540 2748
rect 142596 2746 142620 2748
rect 142676 2746 142700 2748
rect 142538 2694 142540 2746
rect 142602 2694 142614 2746
rect 142676 2694 142678 2746
rect 142516 2692 142540 2694
rect 142596 2692 142620 2694
rect 142676 2692 142700 2694
rect 142460 2672 142756 2692
rect 142816 1850 142844 3538
rect 143356 2984 143408 2990
rect 143356 2926 143408 2932
rect 143368 2582 143396 2926
rect 143356 2576 143408 2582
rect 143356 2518 143408 2524
rect 142988 2304 143040 2310
rect 142988 2246 143040 2252
rect 142632 1822 142844 1850
rect 142632 800 142660 1822
rect 143000 800 143028 2246
rect 143460 2122 143488 4014
rect 143724 3596 143776 3602
rect 143724 3538 143776 3544
rect 143368 2094 143488 2122
rect 143368 800 143396 2094
rect 143736 800 143764 3538
rect 144092 2984 144144 2990
rect 144092 2926 144144 2932
rect 144104 2582 144132 2926
rect 144092 2576 144144 2582
rect 144092 2518 144144 2524
rect 144092 2304 144144 2310
rect 144092 2246 144144 2252
rect 144104 800 144132 2246
rect 144472 800 144500 4014
rect 144828 3596 144880 3602
rect 144828 3538 144880 3544
rect 144840 800 144868 3538
rect 145196 2984 145248 2990
rect 145196 2926 145248 2932
rect 145208 2582 145236 2926
rect 145196 2576 145248 2582
rect 145196 2518 145248 2524
rect 145196 2304 145248 2310
rect 145196 2246 145248 2252
rect 145208 800 145236 2246
rect 145576 800 145604 4014
rect 145932 3596 145984 3602
rect 145932 3538 145984 3544
rect 145944 800 145972 3538
rect 146300 2984 146352 2990
rect 146300 2926 146352 2932
rect 146312 2582 146340 2926
rect 146300 2576 146352 2582
rect 146300 2518 146352 2524
rect 146300 2304 146352 2310
rect 146300 2246 146352 2252
rect 146312 800 146340 2246
rect 146680 800 146708 4014
rect 147036 3596 147088 3602
rect 147036 3538 147088 3544
rect 147048 800 147076 3538
rect 147404 2984 147456 2990
rect 147404 2926 147456 2932
rect 147416 2582 147444 2926
rect 147404 2576 147456 2582
rect 147404 2518 147456 2524
rect 147404 2372 147456 2378
rect 147404 2314 147456 2320
rect 147416 800 147444 2314
rect 147784 800 147812 4014
rect 148140 3596 148192 3602
rect 148140 3538 148192 3544
rect 148152 800 148180 3538
rect 148600 2984 148652 2990
rect 148600 2926 148652 2932
rect 148612 2582 148640 2926
rect 148600 2576 148652 2582
rect 148600 2518 148652 2524
rect 148508 2304 148560 2310
rect 148508 2246 148560 2252
rect 148520 800 148548 2246
rect 148888 800 148916 4014
rect 149244 3596 149296 3602
rect 149244 3538 149296 3544
rect 149980 3596 150032 3602
rect 149980 3538 150032 3544
rect 150348 3596 150400 3602
rect 150348 3538 150400 3544
rect 151176 3596 151228 3602
rect 151176 3538 151228 3544
rect 149256 800 149284 3538
rect 149612 2984 149664 2990
rect 149612 2926 149664 2932
rect 149624 2582 149652 2926
rect 149612 2576 149664 2582
rect 149612 2518 149664 2524
rect 149612 2304 149664 2310
rect 149612 2246 149664 2252
rect 149624 800 149652 2246
rect 149992 800 150020 3538
rect 150360 800 150388 3538
rect 150716 2984 150768 2990
rect 150716 2926 150768 2932
rect 150728 2582 150756 2926
rect 150716 2576 150768 2582
rect 150716 2518 150768 2524
rect 150716 2304 150768 2310
rect 150716 2246 150768 2252
rect 150728 800 150756 2246
rect 151188 1850 151216 3538
rect 151820 2984 151872 2990
rect 151820 2926 151872 2932
rect 151832 2582 151860 2926
rect 151820 2576 151872 2582
rect 151820 2518 151872 2524
rect 151452 2508 151504 2514
rect 151452 2450 151504 2456
rect 151096 1822 151216 1850
rect 151096 800 151124 1822
rect 151464 800 151492 2450
rect 151820 2304 151872 2310
rect 151820 2246 151872 2252
rect 151832 800 151860 2246
rect 152200 800 152228 4014
rect 152556 2984 152608 2990
rect 152556 2926 152608 2932
rect 152568 800 152596 2926
rect 152924 2304 152976 2310
rect 152924 2246 152976 2252
rect 152936 800 152964 2246
rect 153304 800 153332 4014
rect 153660 3596 153712 3602
rect 153660 3538 153712 3544
rect 153672 800 153700 3538
rect 153752 3392 153804 3398
rect 153752 3334 153804 3340
rect 153764 2582 153792 3334
rect 154028 2984 154080 2990
rect 154028 2926 154080 2932
rect 154040 2582 154068 2926
rect 153752 2576 153804 2582
rect 153752 2518 153804 2524
rect 154028 2576 154080 2582
rect 154028 2518 154080 2524
rect 154028 2304 154080 2310
rect 154028 2246 154080 2252
rect 154040 800 154068 2246
rect 154408 800 154436 4014
rect 154764 3596 154816 3602
rect 154764 3538 154816 3544
rect 154776 800 154804 3538
rect 155132 2984 155184 2990
rect 155132 2926 155184 2932
rect 155144 2582 155172 2926
rect 155132 2576 155184 2582
rect 155132 2518 155184 2524
rect 155132 2304 155184 2310
rect 155132 2246 155184 2252
rect 155144 800 155172 2246
rect 155512 800 155540 4014
rect 155868 3596 155920 3602
rect 155868 3538 155920 3544
rect 156604 3596 156656 3602
rect 156604 3538 156656 3544
rect 155880 800 155908 3538
rect 156236 2984 156288 2990
rect 156236 2926 156288 2932
rect 156248 2582 156276 2926
rect 156236 2576 156288 2582
rect 156236 2518 156288 2524
rect 156236 2304 156288 2310
rect 156236 2246 156288 2252
rect 156248 800 156276 2246
rect 156616 800 156644 3538
rect 157340 2984 157392 2990
rect 157340 2926 157392 2932
rect 156972 2916 157024 2922
rect 156972 2858 157024 2864
rect 156984 800 157012 2858
rect 157352 2582 157380 2926
rect 157340 2576 157392 2582
rect 157340 2518 157392 2524
rect 157340 2304 157392 2310
rect 157340 2246 157392 2252
rect 157352 800 157380 2246
rect 157720 800 157748 4014
rect 158168 3596 158220 3602
rect 158168 3538 158220 3544
rect 157820 3292 158116 3312
rect 157876 3290 157900 3292
rect 157956 3290 157980 3292
rect 158036 3290 158060 3292
rect 157898 3238 157900 3290
rect 157962 3238 157974 3290
rect 158036 3238 158038 3290
rect 157876 3236 157900 3238
rect 157956 3236 157980 3238
rect 158036 3236 158060 3238
rect 157820 3216 158116 3236
rect 157820 2204 158116 2224
rect 157876 2202 157900 2204
rect 157956 2202 157980 2204
rect 158036 2202 158060 2204
rect 157898 2150 157900 2202
rect 157962 2150 157974 2202
rect 158036 2150 158038 2202
rect 157876 2148 157900 2150
rect 157956 2148 157980 2150
rect 158036 2148 158060 2150
rect 157820 2128 158116 2148
rect 158180 1850 158208 3538
rect 158444 2304 158496 2310
rect 158444 2246 158496 2252
rect 158088 1822 158208 1850
rect 158088 800 158116 1822
rect 158456 800 158484 2246
rect 158824 800 158852 4014
rect 159180 3596 159232 3602
rect 159180 3538 159232 3544
rect 159088 2984 159140 2990
rect 159088 2926 159140 2932
rect 159100 2582 159128 2926
rect 159088 2576 159140 2582
rect 159088 2518 159140 2524
rect 159192 800 159220 3538
rect 159732 2984 159784 2990
rect 159732 2926 159784 2932
rect 159744 2582 159772 2926
rect 159732 2576 159784 2582
rect 159732 2518 159784 2524
rect 159548 2304 159600 2310
rect 159548 2246 159600 2252
rect 159560 800 159588 2246
rect 159928 800 159956 4014
rect 160284 3596 160336 3602
rect 160284 3538 160336 3544
rect 160296 800 160324 3538
rect 160652 2984 160704 2990
rect 160652 2926 160704 2932
rect 160664 2582 160692 2926
rect 160652 2576 160704 2582
rect 160652 2518 160704 2524
rect 160652 2304 160704 2310
rect 160652 2246 160704 2252
rect 160664 800 160692 2246
rect 161032 800 161060 4014
rect 161388 3596 161440 3602
rect 161388 3538 161440 3544
rect 161400 800 161428 3538
rect 161756 2984 161808 2990
rect 161756 2926 161808 2932
rect 161768 2582 161796 2926
rect 161756 2576 161808 2582
rect 161756 2518 161808 2524
rect 161756 2304 161808 2310
rect 161756 2246 161808 2252
rect 161768 800 161796 2246
rect 162136 800 162164 4014
rect 162492 3596 162544 3602
rect 162492 3538 162544 3544
rect 163596 3596 163648 3602
rect 163596 3538 163648 3544
rect 164424 3596 164476 3602
rect 164424 3538 164476 3544
rect 162504 800 162532 3538
rect 163228 3528 163280 3534
rect 163228 3470 163280 3476
rect 162860 2984 162912 2990
rect 162860 2926 162912 2932
rect 162872 2582 162900 2926
rect 162860 2576 162912 2582
rect 162860 2518 162912 2524
rect 162860 2304 162912 2310
rect 162860 2246 162912 2252
rect 162872 800 162900 2246
rect 163240 800 163268 3470
rect 163608 800 163636 3538
rect 164332 2984 164384 2990
rect 164332 2926 164384 2932
rect 164344 2582 164372 2926
rect 164332 2576 164384 2582
rect 164332 2518 164384 2524
rect 163964 2304 164016 2310
rect 163964 2246 164016 2252
rect 163976 800 164004 2246
rect 164436 1850 164464 3538
rect 165068 2984 165120 2990
rect 165068 2926 165120 2932
rect 165080 2582 165108 2926
rect 165068 2576 165120 2582
rect 165068 2518 165120 2524
rect 164700 2508 164752 2514
rect 164700 2450 164752 2456
rect 164344 1822 164464 1850
rect 164344 800 164372 1822
rect 164712 800 164740 2450
rect 165068 2304 165120 2310
rect 165068 2246 165120 2252
rect 165080 800 165108 2246
rect 165448 800 165476 4014
rect 165804 3596 165856 3602
rect 165804 3538 165856 3544
rect 165816 800 165844 3538
rect 166172 2304 166224 2310
rect 166172 2246 166224 2252
rect 166184 800 166212 2246
rect 166552 800 166580 4014
rect 166908 3596 166960 3602
rect 166908 3538 166960 3544
rect 166920 800 166948 3538
rect 167092 2984 167144 2990
rect 167092 2926 167144 2932
rect 167276 2984 167328 2990
rect 167276 2926 167328 2932
rect 167104 2582 167132 2926
rect 167288 2582 167316 2926
rect 167092 2576 167144 2582
rect 167092 2518 167144 2524
rect 167276 2576 167328 2582
rect 167276 2518 167328 2524
rect 167276 2304 167328 2310
rect 167276 2246 167328 2252
rect 167288 800 167316 2246
rect 167656 800 167684 4014
rect 168012 3596 168064 3602
rect 168012 3538 168064 3544
rect 168024 800 168052 3538
rect 168380 2984 168432 2990
rect 168380 2926 168432 2932
rect 168392 2582 168420 2926
rect 168380 2576 168432 2582
rect 168380 2518 168432 2524
rect 168380 2304 168432 2310
rect 168380 2246 168432 2252
rect 168392 800 168420 2246
rect 168760 800 168788 4014
rect 169116 3596 169168 3602
rect 169116 3538 169168 3544
rect 169128 800 169156 3538
rect 169760 2984 169812 2990
rect 169760 2926 169812 2932
rect 169772 2582 169800 2926
rect 169760 2576 169812 2582
rect 169760 2518 169812 2524
rect 169484 2304 169536 2310
rect 169484 2246 169536 2252
rect 169496 800 169524 2246
rect 169864 800 169892 4014
rect 170220 3596 170272 3602
rect 170220 3538 170272 3544
rect 170956 3596 171008 3602
rect 170956 3538 171008 3544
rect 171324 3596 171376 3602
rect 172152 3596 172204 3602
rect 171324 3538 171376 3544
rect 172072 3556 172152 3584
rect 170232 800 170260 3538
rect 170588 2984 170640 2990
rect 170588 2926 170640 2932
rect 170600 2582 170628 2926
rect 170588 2576 170640 2582
rect 170588 2518 170640 2524
rect 170588 2304 170640 2310
rect 170588 2246 170640 2252
rect 170600 800 170628 2246
rect 170968 800 170996 3538
rect 171336 800 171364 3538
rect 171692 2984 171744 2990
rect 171692 2926 171744 2932
rect 171704 2582 171732 2926
rect 171692 2576 171744 2582
rect 171692 2518 171744 2524
rect 171692 2304 171744 2310
rect 171692 2246 171744 2252
rect 171704 800 171732 2246
rect 172072 800 172100 3556
rect 172152 3538 172204 3544
rect 172796 2984 172848 2990
rect 172796 2926 172848 2932
rect 172428 2916 172480 2922
rect 172428 2858 172480 2864
rect 172440 800 172468 2858
rect 172808 2582 172836 2926
rect 172796 2576 172848 2582
rect 172796 2518 172848 2524
rect 172796 2304 172848 2310
rect 172796 2246 172848 2252
rect 172808 800 172836 2246
rect 173084 1578 173112 4014
rect 173180 3836 173476 3856
rect 173236 3834 173260 3836
rect 173316 3834 173340 3836
rect 173396 3834 173420 3836
rect 173258 3782 173260 3834
rect 173322 3782 173334 3834
rect 173396 3782 173398 3834
rect 173236 3780 173260 3782
rect 173316 3780 173340 3782
rect 173396 3780 173420 3782
rect 173180 3760 173476 3780
rect 173532 3596 173584 3602
rect 173532 3538 173584 3544
rect 173180 2748 173476 2768
rect 173236 2746 173260 2748
rect 173316 2746 173340 2748
rect 173396 2746 173420 2748
rect 173258 2694 173260 2746
rect 173322 2694 173334 2746
rect 173396 2694 173398 2746
rect 173236 2692 173260 2694
rect 173316 2692 173340 2694
rect 173396 2692 173420 2694
rect 173180 2672 173476 2692
rect 173084 1550 173204 1578
rect 173176 800 173204 1550
rect 173544 800 173572 3538
rect 173900 3392 173952 3398
rect 173900 3334 173952 3340
rect 173912 2582 173940 3334
rect 173900 2576 173952 2582
rect 173900 2518 173952 2524
rect 173900 2304 173952 2310
rect 173900 2246 173952 2252
rect 173912 800 173940 2246
rect 174280 800 174308 4014
rect 174636 3596 174688 3602
rect 174636 3538 174688 3544
rect 174648 800 174676 3538
rect 175004 2984 175056 2990
rect 175004 2926 175056 2932
rect 175016 2582 175044 2926
rect 175004 2576 175056 2582
rect 175004 2518 175056 2524
rect 175004 2372 175056 2378
rect 175004 2314 175056 2320
rect 175016 800 175044 2314
rect 175384 800 175412 4626
rect 175740 4072 175792 4078
rect 175740 4014 175792 4020
rect 175752 800 175780 4014
rect 176108 2984 176160 2990
rect 176108 2926 176160 2932
rect 176120 2582 176148 2926
rect 176672 2802 176700 4626
rect 177304 4072 177356 4078
rect 177304 4014 177356 4020
rect 176844 4004 176896 4010
rect 176844 3946 176896 3952
rect 176488 2774 176700 2802
rect 176108 2576 176160 2582
rect 176108 2518 176160 2524
rect 176108 2304 176160 2310
rect 176108 2246 176160 2252
rect 176120 800 176148 2246
rect 176488 800 176516 2774
rect 176856 800 176884 3946
rect 177316 2990 177344 4014
rect 176936 2984 176988 2990
rect 176936 2926 176988 2932
rect 177304 2984 177356 2990
rect 177304 2926 177356 2932
rect 176948 2582 176976 2926
rect 176936 2576 176988 2582
rect 176936 2518 176988 2524
rect 177212 2304 177264 2310
rect 177212 2246 177264 2252
rect 177224 800 177252 2246
rect 177592 800 177620 5102
rect 177948 4684 178000 4690
rect 177948 4626 178000 4632
rect 177960 800 177988 4626
rect 178316 2916 178368 2922
rect 178316 2858 178368 2864
rect 178328 800 178356 2858
rect 178696 800 178724 5714
rect 179052 5160 179104 5166
rect 179052 5102 179104 5108
rect 179064 800 179092 5102
rect 179788 4616 179840 4622
rect 179788 4558 179840 4564
rect 179420 3460 179472 3466
rect 179420 3402 179472 3408
rect 179432 800 179460 3402
rect 179800 800 179828 4558
rect 68836 604 68888 610
rect 68836 546 68888 552
rect 69110 0 69166 800
rect 69478 0 69534 800
rect 69846 0 69902 800
rect 70214 0 70270 800
rect 70582 0 70638 800
rect 70950 0 71006 800
rect 71318 0 71374 800
rect 71686 0 71742 800
rect 72054 0 72110 800
rect 72422 0 72478 800
rect 72790 0 72846 800
rect 73158 0 73214 800
rect 73526 0 73582 800
rect 73894 0 73950 800
rect 74262 0 74318 800
rect 74630 0 74686 800
rect 74998 0 75054 800
rect 75366 0 75422 800
rect 75734 0 75790 800
rect 76102 0 76158 800
rect 76470 0 76526 800
rect 76838 0 76894 800
rect 77206 0 77262 800
rect 77574 0 77630 800
rect 77942 0 77998 800
rect 78310 0 78366 800
rect 78678 0 78734 800
rect 79046 0 79102 800
rect 79414 0 79470 800
rect 79782 0 79838 800
rect 80150 0 80206 800
rect 80518 0 80574 800
rect 80886 0 80942 800
rect 81254 0 81310 800
rect 81622 0 81678 800
rect 81990 0 82046 800
rect 82358 0 82414 800
rect 82726 0 82782 800
rect 83094 0 83150 800
rect 83462 0 83518 800
rect 83830 0 83886 800
rect 84198 0 84254 800
rect 84566 0 84622 800
rect 84934 0 84990 800
rect 85302 0 85358 800
rect 85670 0 85726 800
rect 86038 0 86094 800
rect 86406 0 86462 800
rect 86774 0 86830 800
rect 87142 0 87198 800
rect 87510 0 87566 800
rect 87878 0 87934 800
rect 88246 0 88302 800
rect 88614 0 88670 800
rect 88982 0 89038 800
rect 89350 0 89406 800
rect 89718 0 89774 800
rect 90086 0 90142 800
rect 90454 0 90510 800
rect 90822 0 90878 800
rect 91190 0 91246 800
rect 91558 0 91614 800
rect 91926 0 91982 800
rect 92294 0 92350 800
rect 92662 0 92718 800
rect 93030 0 93086 800
rect 93398 0 93454 800
rect 93766 0 93822 800
rect 94134 0 94190 800
rect 94502 0 94558 800
rect 94870 0 94926 800
rect 95238 0 95294 800
rect 95606 0 95662 800
rect 95974 0 96030 800
rect 96342 0 96398 800
rect 96710 0 96766 800
rect 97078 0 97134 800
rect 97446 0 97502 800
rect 97814 0 97870 800
rect 98182 0 98238 800
rect 98550 0 98606 800
rect 98918 0 98974 800
rect 99286 0 99342 800
rect 99654 0 99710 800
rect 100022 0 100078 800
rect 100390 0 100446 800
rect 100758 0 100814 800
rect 101126 0 101182 800
rect 101494 0 101550 800
rect 101862 0 101918 800
rect 102230 0 102286 800
rect 102598 0 102654 800
rect 102966 0 103022 800
rect 103334 0 103390 800
rect 103702 0 103758 800
rect 104070 0 104126 800
rect 104438 0 104494 800
rect 104806 0 104862 800
rect 105174 0 105230 800
rect 105542 0 105598 800
rect 105910 0 105966 800
rect 106278 0 106334 800
rect 106646 0 106702 800
rect 107014 0 107070 800
rect 107382 0 107438 800
rect 107750 0 107806 800
rect 108118 0 108174 800
rect 108486 0 108542 800
rect 108854 0 108910 800
rect 109222 0 109278 800
rect 109590 0 109646 800
rect 109958 0 110014 800
rect 110326 0 110382 800
rect 110694 0 110750 800
rect 111062 0 111118 800
rect 111430 0 111486 800
rect 111798 0 111854 800
rect 112166 0 112222 800
rect 112534 0 112590 800
rect 112902 0 112958 800
rect 113270 0 113326 800
rect 113638 0 113694 800
rect 114006 0 114062 800
rect 114374 0 114430 800
rect 114742 0 114798 800
rect 115110 0 115166 800
rect 115478 0 115534 800
rect 115846 0 115902 800
rect 116214 0 116270 800
rect 116582 0 116638 800
rect 116950 0 117006 800
rect 117318 0 117374 800
rect 117686 0 117742 800
rect 118054 0 118110 800
rect 118422 0 118478 800
rect 118790 0 118846 800
rect 119158 0 119214 800
rect 119526 0 119582 800
rect 119894 0 119950 800
rect 120170 0 120226 800
rect 120538 0 120594 800
rect 120906 0 120962 800
rect 121274 0 121330 800
rect 121642 0 121698 800
rect 122010 0 122066 800
rect 122378 0 122434 800
rect 122746 0 122802 800
rect 123114 0 123170 800
rect 123482 0 123538 800
rect 123850 0 123906 800
rect 124218 0 124274 800
rect 124586 0 124642 800
rect 124954 0 125010 800
rect 125322 0 125378 800
rect 125690 0 125746 800
rect 126058 0 126114 800
rect 126426 0 126482 800
rect 126794 0 126850 800
rect 127162 0 127218 800
rect 127530 0 127586 800
rect 127898 0 127954 800
rect 128266 0 128322 800
rect 128634 0 128690 800
rect 129002 0 129058 800
rect 129370 0 129426 800
rect 129738 0 129794 800
rect 130106 0 130162 800
rect 130474 0 130530 800
rect 130842 0 130898 800
rect 131210 0 131266 800
rect 131578 0 131634 800
rect 131946 0 132002 800
rect 132314 0 132370 800
rect 132682 0 132738 800
rect 133050 0 133106 800
rect 133418 0 133474 800
rect 133786 0 133842 800
rect 134154 0 134210 800
rect 134522 0 134578 800
rect 134890 0 134946 800
rect 135258 0 135314 800
rect 135626 0 135682 800
rect 135994 0 136050 800
rect 136362 0 136418 800
rect 136730 0 136786 800
rect 137098 0 137154 800
rect 137466 0 137522 800
rect 137834 0 137890 800
rect 138202 0 138258 800
rect 138570 0 138626 800
rect 138938 0 138994 800
rect 139306 0 139362 800
rect 139674 0 139730 800
rect 140042 0 140098 800
rect 140410 0 140466 800
rect 140778 0 140834 800
rect 141146 0 141202 800
rect 141514 0 141570 800
rect 141882 0 141938 800
rect 142250 0 142306 800
rect 142618 0 142674 800
rect 142986 0 143042 800
rect 143354 0 143410 800
rect 143722 0 143778 800
rect 144090 0 144146 800
rect 144458 0 144514 800
rect 144826 0 144882 800
rect 145194 0 145250 800
rect 145562 0 145618 800
rect 145930 0 145986 800
rect 146298 0 146354 800
rect 146666 0 146722 800
rect 147034 0 147090 800
rect 147402 0 147458 800
rect 147770 0 147826 800
rect 148138 0 148194 800
rect 148506 0 148562 800
rect 148874 0 148930 800
rect 149242 0 149298 800
rect 149610 0 149666 800
rect 149978 0 150034 800
rect 150346 0 150402 800
rect 150714 0 150770 800
rect 151082 0 151138 800
rect 151450 0 151506 800
rect 151818 0 151874 800
rect 152186 0 152242 800
rect 152554 0 152610 800
rect 152922 0 152978 800
rect 153290 0 153346 800
rect 153658 0 153714 800
rect 154026 0 154082 800
rect 154394 0 154450 800
rect 154762 0 154818 800
rect 155130 0 155186 800
rect 155498 0 155554 800
rect 155866 0 155922 800
rect 156234 0 156290 800
rect 156602 0 156658 800
rect 156970 0 157026 800
rect 157338 0 157394 800
rect 157706 0 157762 800
rect 158074 0 158130 800
rect 158442 0 158498 800
rect 158810 0 158866 800
rect 159178 0 159234 800
rect 159546 0 159602 800
rect 159914 0 159970 800
rect 160282 0 160338 800
rect 160650 0 160706 800
rect 161018 0 161074 800
rect 161386 0 161442 800
rect 161754 0 161810 800
rect 162122 0 162178 800
rect 162490 0 162546 800
rect 162858 0 162914 800
rect 163226 0 163282 800
rect 163594 0 163650 800
rect 163962 0 164018 800
rect 164330 0 164386 800
rect 164698 0 164754 800
rect 165066 0 165122 800
rect 165434 0 165490 800
rect 165802 0 165858 800
rect 166170 0 166226 800
rect 166538 0 166594 800
rect 166906 0 166962 800
rect 167274 0 167330 800
rect 167642 0 167698 800
rect 168010 0 168066 800
rect 168378 0 168434 800
rect 168746 0 168802 800
rect 169114 0 169170 800
rect 169482 0 169538 800
rect 169850 0 169906 800
rect 170218 0 170274 800
rect 170586 0 170642 800
rect 170954 0 171010 800
rect 171322 0 171378 800
rect 171690 0 171746 800
rect 172058 0 172114 800
rect 172426 0 172482 800
rect 172794 0 172850 800
rect 173162 0 173218 800
rect 173530 0 173586 800
rect 173898 0 173954 800
rect 174266 0 174322 800
rect 174634 0 174690 800
rect 175002 0 175058 800
rect 175370 0 175426 800
rect 175738 0 175794 800
rect 176106 0 176162 800
rect 176474 0 176530 800
rect 176842 0 176898 800
rect 177210 0 177266 800
rect 177578 0 177634 800
rect 177946 0 178002 800
rect 178314 0 178370 800
rect 178682 0 178738 800
rect 179050 0 179106 800
rect 179418 0 179474 800
rect 179786 0 179842 800
<< via2 >>
rect 4220 117530 4276 117532
rect 4300 117530 4356 117532
rect 4380 117530 4436 117532
rect 4460 117530 4516 117532
rect 4220 117478 4246 117530
rect 4246 117478 4276 117530
rect 4300 117478 4310 117530
rect 4310 117478 4356 117530
rect 4380 117478 4426 117530
rect 4426 117478 4436 117530
rect 4460 117478 4490 117530
rect 4490 117478 4516 117530
rect 4220 117476 4276 117478
rect 4300 117476 4356 117478
rect 4380 117476 4436 117478
rect 4460 117476 4516 117478
rect 34940 117530 34996 117532
rect 35020 117530 35076 117532
rect 35100 117530 35156 117532
rect 35180 117530 35236 117532
rect 34940 117478 34966 117530
rect 34966 117478 34996 117530
rect 35020 117478 35030 117530
rect 35030 117478 35076 117530
rect 35100 117478 35146 117530
rect 35146 117478 35156 117530
rect 35180 117478 35210 117530
rect 35210 117478 35236 117530
rect 34940 117476 34996 117478
rect 35020 117476 35076 117478
rect 35100 117476 35156 117478
rect 35180 117476 35236 117478
rect 65660 117530 65716 117532
rect 65740 117530 65796 117532
rect 65820 117530 65876 117532
rect 65900 117530 65956 117532
rect 65660 117478 65686 117530
rect 65686 117478 65716 117530
rect 65740 117478 65750 117530
rect 65750 117478 65796 117530
rect 65820 117478 65866 117530
rect 65866 117478 65876 117530
rect 65900 117478 65930 117530
rect 65930 117478 65956 117530
rect 65660 117476 65716 117478
rect 65740 117476 65796 117478
rect 65820 117476 65876 117478
rect 65900 117476 65956 117478
rect 96380 117530 96436 117532
rect 96460 117530 96516 117532
rect 96540 117530 96596 117532
rect 96620 117530 96676 117532
rect 96380 117478 96406 117530
rect 96406 117478 96436 117530
rect 96460 117478 96470 117530
rect 96470 117478 96516 117530
rect 96540 117478 96586 117530
rect 96586 117478 96596 117530
rect 96620 117478 96650 117530
rect 96650 117478 96676 117530
rect 96380 117476 96436 117478
rect 96460 117476 96516 117478
rect 96540 117476 96596 117478
rect 96620 117476 96676 117478
rect 127100 117530 127156 117532
rect 127180 117530 127236 117532
rect 127260 117530 127316 117532
rect 127340 117530 127396 117532
rect 127100 117478 127126 117530
rect 127126 117478 127156 117530
rect 127180 117478 127190 117530
rect 127190 117478 127236 117530
rect 127260 117478 127306 117530
rect 127306 117478 127316 117530
rect 127340 117478 127370 117530
rect 127370 117478 127396 117530
rect 127100 117476 127156 117478
rect 127180 117476 127236 117478
rect 127260 117476 127316 117478
rect 127340 117476 127396 117478
rect 157820 117530 157876 117532
rect 157900 117530 157956 117532
rect 157980 117530 158036 117532
rect 158060 117530 158116 117532
rect 157820 117478 157846 117530
rect 157846 117478 157876 117530
rect 157900 117478 157910 117530
rect 157910 117478 157956 117530
rect 157980 117478 158026 117530
rect 158026 117478 158036 117530
rect 158060 117478 158090 117530
rect 158090 117478 158116 117530
rect 157820 117476 157876 117478
rect 157900 117476 157956 117478
rect 157980 117476 158036 117478
rect 158060 117476 158116 117478
rect 4220 116442 4276 116444
rect 4300 116442 4356 116444
rect 4380 116442 4436 116444
rect 4460 116442 4516 116444
rect 4220 116390 4246 116442
rect 4246 116390 4276 116442
rect 4300 116390 4310 116442
rect 4310 116390 4356 116442
rect 4380 116390 4426 116442
rect 4426 116390 4436 116442
rect 4460 116390 4490 116442
rect 4490 116390 4516 116442
rect 4220 116388 4276 116390
rect 4300 116388 4356 116390
rect 4380 116388 4436 116390
rect 4460 116388 4516 116390
rect 19580 116986 19636 116988
rect 19660 116986 19716 116988
rect 19740 116986 19796 116988
rect 19820 116986 19876 116988
rect 19580 116934 19606 116986
rect 19606 116934 19636 116986
rect 19660 116934 19670 116986
rect 19670 116934 19716 116986
rect 19740 116934 19786 116986
rect 19786 116934 19796 116986
rect 19820 116934 19850 116986
rect 19850 116934 19876 116986
rect 19580 116932 19636 116934
rect 19660 116932 19716 116934
rect 19740 116932 19796 116934
rect 19820 116932 19876 116934
rect 19580 115898 19636 115900
rect 19660 115898 19716 115900
rect 19740 115898 19796 115900
rect 19820 115898 19876 115900
rect 19580 115846 19606 115898
rect 19606 115846 19636 115898
rect 19660 115846 19670 115898
rect 19670 115846 19716 115898
rect 19740 115846 19786 115898
rect 19786 115846 19796 115898
rect 19820 115846 19850 115898
rect 19850 115846 19876 115898
rect 19580 115844 19636 115846
rect 19660 115844 19716 115846
rect 19740 115844 19796 115846
rect 19820 115844 19876 115846
rect 4220 115354 4276 115356
rect 4300 115354 4356 115356
rect 4380 115354 4436 115356
rect 4460 115354 4516 115356
rect 4220 115302 4246 115354
rect 4246 115302 4276 115354
rect 4300 115302 4310 115354
rect 4310 115302 4356 115354
rect 4380 115302 4426 115354
rect 4426 115302 4436 115354
rect 4460 115302 4490 115354
rect 4490 115302 4516 115354
rect 4220 115300 4276 115302
rect 4300 115300 4356 115302
rect 4380 115300 4436 115302
rect 4460 115300 4516 115302
rect 19580 114810 19636 114812
rect 19660 114810 19716 114812
rect 19740 114810 19796 114812
rect 19820 114810 19876 114812
rect 19580 114758 19606 114810
rect 19606 114758 19636 114810
rect 19660 114758 19670 114810
rect 19670 114758 19716 114810
rect 19740 114758 19786 114810
rect 19786 114758 19796 114810
rect 19820 114758 19850 114810
rect 19850 114758 19876 114810
rect 19580 114756 19636 114758
rect 19660 114756 19716 114758
rect 19740 114756 19796 114758
rect 19820 114756 19876 114758
rect 4220 114266 4276 114268
rect 4300 114266 4356 114268
rect 4380 114266 4436 114268
rect 4460 114266 4516 114268
rect 4220 114214 4246 114266
rect 4246 114214 4276 114266
rect 4300 114214 4310 114266
rect 4310 114214 4356 114266
rect 4380 114214 4426 114266
rect 4426 114214 4436 114266
rect 4460 114214 4490 114266
rect 4490 114214 4516 114266
rect 4220 114212 4276 114214
rect 4300 114212 4356 114214
rect 4380 114212 4436 114214
rect 4460 114212 4516 114214
rect 19580 113722 19636 113724
rect 19660 113722 19716 113724
rect 19740 113722 19796 113724
rect 19820 113722 19876 113724
rect 19580 113670 19606 113722
rect 19606 113670 19636 113722
rect 19660 113670 19670 113722
rect 19670 113670 19716 113722
rect 19740 113670 19786 113722
rect 19786 113670 19796 113722
rect 19820 113670 19850 113722
rect 19850 113670 19876 113722
rect 19580 113668 19636 113670
rect 19660 113668 19716 113670
rect 19740 113668 19796 113670
rect 19820 113668 19876 113670
rect 4220 113178 4276 113180
rect 4300 113178 4356 113180
rect 4380 113178 4436 113180
rect 4460 113178 4516 113180
rect 4220 113126 4246 113178
rect 4246 113126 4276 113178
rect 4300 113126 4310 113178
rect 4310 113126 4356 113178
rect 4380 113126 4426 113178
rect 4426 113126 4436 113178
rect 4460 113126 4490 113178
rect 4490 113126 4516 113178
rect 4220 113124 4276 113126
rect 4300 113124 4356 113126
rect 4380 113124 4436 113126
rect 4460 113124 4516 113126
rect 19580 112634 19636 112636
rect 19660 112634 19716 112636
rect 19740 112634 19796 112636
rect 19820 112634 19876 112636
rect 19580 112582 19606 112634
rect 19606 112582 19636 112634
rect 19660 112582 19670 112634
rect 19670 112582 19716 112634
rect 19740 112582 19786 112634
rect 19786 112582 19796 112634
rect 19820 112582 19850 112634
rect 19850 112582 19876 112634
rect 19580 112580 19636 112582
rect 19660 112580 19716 112582
rect 19740 112580 19796 112582
rect 19820 112580 19876 112582
rect 4220 112090 4276 112092
rect 4300 112090 4356 112092
rect 4380 112090 4436 112092
rect 4460 112090 4516 112092
rect 4220 112038 4246 112090
rect 4246 112038 4276 112090
rect 4300 112038 4310 112090
rect 4310 112038 4356 112090
rect 4380 112038 4426 112090
rect 4426 112038 4436 112090
rect 4460 112038 4490 112090
rect 4490 112038 4516 112090
rect 4220 112036 4276 112038
rect 4300 112036 4356 112038
rect 4380 112036 4436 112038
rect 4460 112036 4516 112038
rect 19580 111546 19636 111548
rect 19660 111546 19716 111548
rect 19740 111546 19796 111548
rect 19820 111546 19876 111548
rect 19580 111494 19606 111546
rect 19606 111494 19636 111546
rect 19660 111494 19670 111546
rect 19670 111494 19716 111546
rect 19740 111494 19786 111546
rect 19786 111494 19796 111546
rect 19820 111494 19850 111546
rect 19850 111494 19876 111546
rect 19580 111492 19636 111494
rect 19660 111492 19716 111494
rect 19740 111492 19796 111494
rect 19820 111492 19876 111494
rect 4220 111002 4276 111004
rect 4300 111002 4356 111004
rect 4380 111002 4436 111004
rect 4460 111002 4516 111004
rect 4220 110950 4246 111002
rect 4246 110950 4276 111002
rect 4300 110950 4310 111002
rect 4310 110950 4356 111002
rect 4380 110950 4426 111002
rect 4426 110950 4436 111002
rect 4460 110950 4490 111002
rect 4490 110950 4516 111002
rect 4220 110948 4276 110950
rect 4300 110948 4356 110950
rect 4380 110948 4436 110950
rect 4460 110948 4516 110950
rect 19580 110458 19636 110460
rect 19660 110458 19716 110460
rect 19740 110458 19796 110460
rect 19820 110458 19876 110460
rect 19580 110406 19606 110458
rect 19606 110406 19636 110458
rect 19660 110406 19670 110458
rect 19670 110406 19716 110458
rect 19740 110406 19786 110458
rect 19786 110406 19796 110458
rect 19820 110406 19850 110458
rect 19850 110406 19876 110458
rect 19580 110404 19636 110406
rect 19660 110404 19716 110406
rect 19740 110404 19796 110406
rect 19820 110404 19876 110406
rect 4220 109914 4276 109916
rect 4300 109914 4356 109916
rect 4380 109914 4436 109916
rect 4460 109914 4516 109916
rect 4220 109862 4246 109914
rect 4246 109862 4276 109914
rect 4300 109862 4310 109914
rect 4310 109862 4356 109914
rect 4380 109862 4426 109914
rect 4426 109862 4436 109914
rect 4460 109862 4490 109914
rect 4490 109862 4516 109914
rect 4220 109860 4276 109862
rect 4300 109860 4356 109862
rect 4380 109860 4436 109862
rect 4460 109860 4516 109862
rect 19580 109370 19636 109372
rect 19660 109370 19716 109372
rect 19740 109370 19796 109372
rect 19820 109370 19876 109372
rect 19580 109318 19606 109370
rect 19606 109318 19636 109370
rect 19660 109318 19670 109370
rect 19670 109318 19716 109370
rect 19740 109318 19786 109370
rect 19786 109318 19796 109370
rect 19820 109318 19850 109370
rect 19850 109318 19876 109370
rect 19580 109316 19636 109318
rect 19660 109316 19716 109318
rect 19740 109316 19796 109318
rect 19820 109316 19876 109318
rect 4220 108826 4276 108828
rect 4300 108826 4356 108828
rect 4380 108826 4436 108828
rect 4460 108826 4516 108828
rect 4220 108774 4246 108826
rect 4246 108774 4276 108826
rect 4300 108774 4310 108826
rect 4310 108774 4356 108826
rect 4380 108774 4426 108826
rect 4426 108774 4436 108826
rect 4460 108774 4490 108826
rect 4490 108774 4516 108826
rect 4220 108772 4276 108774
rect 4300 108772 4356 108774
rect 4380 108772 4436 108774
rect 4460 108772 4516 108774
rect 19580 108282 19636 108284
rect 19660 108282 19716 108284
rect 19740 108282 19796 108284
rect 19820 108282 19876 108284
rect 19580 108230 19606 108282
rect 19606 108230 19636 108282
rect 19660 108230 19670 108282
rect 19670 108230 19716 108282
rect 19740 108230 19786 108282
rect 19786 108230 19796 108282
rect 19820 108230 19850 108282
rect 19850 108230 19876 108282
rect 19580 108228 19636 108230
rect 19660 108228 19716 108230
rect 19740 108228 19796 108230
rect 19820 108228 19876 108230
rect 4220 107738 4276 107740
rect 4300 107738 4356 107740
rect 4380 107738 4436 107740
rect 4460 107738 4516 107740
rect 4220 107686 4246 107738
rect 4246 107686 4276 107738
rect 4300 107686 4310 107738
rect 4310 107686 4356 107738
rect 4380 107686 4426 107738
rect 4426 107686 4436 107738
rect 4460 107686 4490 107738
rect 4490 107686 4516 107738
rect 4220 107684 4276 107686
rect 4300 107684 4356 107686
rect 4380 107684 4436 107686
rect 4460 107684 4516 107686
rect 19580 107194 19636 107196
rect 19660 107194 19716 107196
rect 19740 107194 19796 107196
rect 19820 107194 19876 107196
rect 19580 107142 19606 107194
rect 19606 107142 19636 107194
rect 19660 107142 19670 107194
rect 19670 107142 19716 107194
rect 19740 107142 19786 107194
rect 19786 107142 19796 107194
rect 19820 107142 19850 107194
rect 19850 107142 19876 107194
rect 19580 107140 19636 107142
rect 19660 107140 19716 107142
rect 19740 107140 19796 107142
rect 19820 107140 19876 107142
rect 4220 106650 4276 106652
rect 4300 106650 4356 106652
rect 4380 106650 4436 106652
rect 4460 106650 4516 106652
rect 4220 106598 4246 106650
rect 4246 106598 4276 106650
rect 4300 106598 4310 106650
rect 4310 106598 4356 106650
rect 4380 106598 4426 106650
rect 4426 106598 4436 106650
rect 4460 106598 4490 106650
rect 4490 106598 4516 106650
rect 4220 106596 4276 106598
rect 4300 106596 4356 106598
rect 4380 106596 4436 106598
rect 4460 106596 4516 106598
rect 19580 106106 19636 106108
rect 19660 106106 19716 106108
rect 19740 106106 19796 106108
rect 19820 106106 19876 106108
rect 19580 106054 19606 106106
rect 19606 106054 19636 106106
rect 19660 106054 19670 106106
rect 19670 106054 19716 106106
rect 19740 106054 19786 106106
rect 19786 106054 19796 106106
rect 19820 106054 19850 106106
rect 19850 106054 19876 106106
rect 19580 106052 19636 106054
rect 19660 106052 19716 106054
rect 19740 106052 19796 106054
rect 19820 106052 19876 106054
rect 4220 105562 4276 105564
rect 4300 105562 4356 105564
rect 4380 105562 4436 105564
rect 4460 105562 4516 105564
rect 4220 105510 4246 105562
rect 4246 105510 4276 105562
rect 4300 105510 4310 105562
rect 4310 105510 4356 105562
rect 4380 105510 4426 105562
rect 4426 105510 4436 105562
rect 4460 105510 4490 105562
rect 4490 105510 4516 105562
rect 4220 105508 4276 105510
rect 4300 105508 4356 105510
rect 4380 105508 4436 105510
rect 4460 105508 4516 105510
rect 19580 105018 19636 105020
rect 19660 105018 19716 105020
rect 19740 105018 19796 105020
rect 19820 105018 19876 105020
rect 19580 104966 19606 105018
rect 19606 104966 19636 105018
rect 19660 104966 19670 105018
rect 19670 104966 19716 105018
rect 19740 104966 19786 105018
rect 19786 104966 19796 105018
rect 19820 104966 19850 105018
rect 19850 104966 19876 105018
rect 19580 104964 19636 104966
rect 19660 104964 19716 104966
rect 19740 104964 19796 104966
rect 19820 104964 19876 104966
rect 4220 104474 4276 104476
rect 4300 104474 4356 104476
rect 4380 104474 4436 104476
rect 4460 104474 4516 104476
rect 4220 104422 4246 104474
rect 4246 104422 4276 104474
rect 4300 104422 4310 104474
rect 4310 104422 4356 104474
rect 4380 104422 4426 104474
rect 4426 104422 4436 104474
rect 4460 104422 4490 104474
rect 4490 104422 4516 104474
rect 4220 104420 4276 104422
rect 4300 104420 4356 104422
rect 4380 104420 4436 104422
rect 4460 104420 4516 104422
rect 19580 103930 19636 103932
rect 19660 103930 19716 103932
rect 19740 103930 19796 103932
rect 19820 103930 19876 103932
rect 19580 103878 19606 103930
rect 19606 103878 19636 103930
rect 19660 103878 19670 103930
rect 19670 103878 19716 103930
rect 19740 103878 19786 103930
rect 19786 103878 19796 103930
rect 19820 103878 19850 103930
rect 19850 103878 19876 103930
rect 19580 103876 19636 103878
rect 19660 103876 19716 103878
rect 19740 103876 19796 103878
rect 19820 103876 19876 103878
rect 4220 103386 4276 103388
rect 4300 103386 4356 103388
rect 4380 103386 4436 103388
rect 4460 103386 4516 103388
rect 4220 103334 4246 103386
rect 4246 103334 4276 103386
rect 4300 103334 4310 103386
rect 4310 103334 4356 103386
rect 4380 103334 4426 103386
rect 4426 103334 4436 103386
rect 4460 103334 4490 103386
rect 4490 103334 4516 103386
rect 4220 103332 4276 103334
rect 4300 103332 4356 103334
rect 4380 103332 4436 103334
rect 4460 103332 4516 103334
rect 19580 102842 19636 102844
rect 19660 102842 19716 102844
rect 19740 102842 19796 102844
rect 19820 102842 19876 102844
rect 19580 102790 19606 102842
rect 19606 102790 19636 102842
rect 19660 102790 19670 102842
rect 19670 102790 19716 102842
rect 19740 102790 19786 102842
rect 19786 102790 19796 102842
rect 19820 102790 19850 102842
rect 19850 102790 19876 102842
rect 19580 102788 19636 102790
rect 19660 102788 19716 102790
rect 19740 102788 19796 102790
rect 19820 102788 19876 102790
rect 4220 102298 4276 102300
rect 4300 102298 4356 102300
rect 4380 102298 4436 102300
rect 4460 102298 4516 102300
rect 4220 102246 4246 102298
rect 4246 102246 4276 102298
rect 4300 102246 4310 102298
rect 4310 102246 4356 102298
rect 4380 102246 4426 102298
rect 4426 102246 4436 102298
rect 4460 102246 4490 102298
rect 4490 102246 4516 102298
rect 4220 102244 4276 102246
rect 4300 102244 4356 102246
rect 4380 102244 4436 102246
rect 4460 102244 4516 102246
rect 19580 101754 19636 101756
rect 19660 101754 19716 101756
rect 19740 101754 19796 101756
rect 19820 101754 19876 101756
rect 19580 101702 19606 101754
rect 19606 101702 19636 101754
rect 19660 101702 19670 101754
rect 19670 101702 19716 101754
rect 19740 101702 19786 101754
rect 19786 101702 19796 101754
rect 19820 101702 19850 101754
rect 19850 101702 19876 101754
rect 19580 101700 19636 101702
rect 19660 101700 19716 101702
rect 19740 101700 19796 101702
rect 19820 101700 19876 101702
rect 4220 101210 4276 101212
rect 4300 101210 4356 101212
rect 4380 101210 4436 101212
rect 4460 101210 4516 101212
rect 4220 101158 4246 101210
rect 4246 101158 4276 101210
rect 4300 101158 4310 101210
rect 4310 101158 4356 101210
rect 4380 101158 4426 101210
rect 4426 101158 4436 101210
rect 4460 101158 4490 101210
rect 4490 101158 4516 101210
rect 4220 101156 4276 101158
rect 4300 101156 4356 101158
rect 4380 101156 4436 101158
rect 4460 101156 4516 101158
rect 19580 100666 19636 100668
rect 19660 100666 19716 100668
rect 19740 100666 19796 100668
rect 19820 100666 19876 100668
rect 19580 100614 19606 100666
rect 19606 100614 19636 100666
rect 19660 100614 19670 100666
rect 19670 100614 19716 100666
rect 19740 100614 19786 100666
rect 19786 100614 19796 100666
rect 19820 100614 19850 100666
rect 19850 100614 19876 100666
rect 19580 100612 19636 100614
rect 19660 100612 19716 100614
rect 19740 100612 19796 100614
rect 19820 100612 19876 100614
rect 4220 100122 4276 100124
rect 4300 100122 4356 100124
rect 4380 100122 4436 100124
rect 4460 100122 4516 100124
rect 4220 100070 4246 100122
rect 4246 100070 4276 100122
rect 4300 100070 4310 100122
rect 4310 100070 4356 100122
rect 4380 100070 4426 100122
rect 4426 100070 4436 100122
rect 4460 100070 4490 100122
rect 4490 100070 4516 100122
rect 4220 100068 4276 100070
rect 4300 100068 4356 100070
rect 4380 100068 4436 100070
rect 4460 100068 4516 100070
rect 19580 99578 19636 99580
rect 19660 99578 19716 99580
rect 19740 99578 19796 99580
rect 19820 99578 19876 99580
rect 19580 99526 19606 99578
rect 19606 99526 19636 99578
rect 19660 99526 19670 99578
rect 19670 99526 19716 99578
rect 19740 99526 19786 99578
rect 19786 99526 19796 99578
rect 19820 99526 19850 99578
rect 19850 99526 19876 99578
rect 19580 99524 19636 99526
rect 19660 99524 19716 99526
rect 19740 99524 19796 99526
rect 19820 99524 19876 99526
rect 4220 99034 4276 99036
rect 4300 99034 4356 99036
rect 4380 99034 4436 99036
rect 4460 99034 4516 99036
rect 4220 98982 4246 99034
rect 4246 98982 4276 99034
rect 4300 98982 4310 99034
rect 4310 98982 4356 99034
rect 4380 98982 4426 99034
rect 4426 98982 4436 99034
rect 4460 98982 4490 99034
rect 4490 98982 4516 99034
rect 4220 98980 4276 98982
rect 4300 98980 4356 98982
rect 4380 98980 4436 98982
rect 4460 98980 4516 98982
rect 19580 98490 19636 98492
rect 19660 98490 19716 98492
rect 19740 98490 19796 98492
rect 19820 98490 19876 98492
rect 19580 98438 19606 98490
rect 19606 98438 19636 98490
rect 19660 98438 19670 98490
rect 19670 98438 19716 98490
rect 19740 98438 19786 98490
rect 19786 98438 19796 98490
rect 19820 98438 19850 98490
rect 19850 98438 19876 98490
rect 19580 98436 19636 98438
rect 19660 98436 19716 98438
rect 19740 98436 19796 98438
rect 19820 98436 19876 98438
rect 4220 97946 4276 97948
rect 4300 97946 4356 97948
rect 4380 97946 4436 97948
rect 4460 97946 4516 97948
rect 4220 97894 4246 97946
rect 4246 97894 4276 97946
rect 4300 97894 4310 97946
rect 4310 97894 4356 97946
rect 4380 97894 4426 97946
rect 4426 97894 4436 97946
rect 4460 97894 4490 97946
rect 4490 97894 4516 97946
rect 4220 97892 4276 97894
rect 4300 97892 4356 97894
rect 4380 97892 4436 97894
rect 4460 97892 4516 97894
rect 19580 97402 19636 97404
rect 19660 97402 19716 97404
rect 19740 97402 19796 97404
rect 19820 97402 19876 97404
rect 19580 97350 19606 97402
rect 19606 97350 19636 97402
rect 19660 97350 19670 97402
rect 19670 97350 19716 97402
rect 19740 97350 19786 97402
rect 19786 97350 19796 97402
rect 19820 97350 19850 97402
rect 19850 97350 19876 97402
rect 19580 97348 19636 97350
rect 19660 97348 19716 97350
rect 19740 97348 19796 97350
rect 19820 97348 19876 97350
rect 4220 96858 4276 96860
rect 4300 96858 4356 96860
rect 4380 96858 4436 96860
rect 4460 96858 4516 96860
rect 4220 96806 4246 96858
rect 4246 96806 4276 96858
rect 4300 96806 4310 96858
rect 4310 96806 4356 96858
rect 4380 96806 4426 96858
rect 4426 96806 4436 96858
rect 4460 96806 4490 96858
rect 4490 96806 4516 96858
rect 4220 96804 4276 96806
rect 4300 96804 4356 96806
rect 4380 96804 4436 96806
rect 4460 96804 4516 96806
rect 19580 96314 19636 96316
rect 19660 96314 19716 96316
rect 19740 96314 19796 96316
rect 19820 96314 19876 96316
rect 19580 96262 19606 96314
rect 19606 96262 19636 96314
rect 19660 96262 19670 96314
rect 19670 96262 19716 96314
rect 19740 96262 19786 96314
rect 19786 96262 19796 96314
rect 19820 96262 19850 96314
rect 19850 96262 19876 96314
rect 19580 96260 19636 96262
rect 19660 96260 19716 96262
rect 19740 96260 19796 96262
rect 19820 96260 19876 96262
rect 4220 95770 4276 95772
rect 4300 95770 4356 95772
rect 4380 95770 4436 95772
rect 4460 95770 4516 95772
rect 4220 95718 4246 95770
rect 4246 95718 4276 95770
rect 4300 95718 4310 95770
rect 4310 95718 4356 95770
rect 4380 95718 4426 95770
rect 4426 95718 4436 95770
rect 4460 95718 4490 95770
rect 4490 95718 4516 95770
rect 4220 95716 4276 95718
rect 4300 95716 4356 95718
rect 4380 95716 4436 95718
rect 4460 95716 4516 95718
rect 19580 95226 19636 95228
rect 19660 95226 19716 95228
rect 19740 95226 19796 95228
rect 19820 95226 19876 95228
rect 19580 95174 19606 95226
rect 19606 95174 19636 95226
rect 19660 95174 19670 95226
rect 19670 95174 19716 95226
rect 19740 95174 19786 95226
rect 19786 95174 19796 95226
rect 19820 95174 19850 95226
rect 19850 95174 19876 95226
rect 19580 95172 19636 95174
rect 19660 95172 19716 95174
rect 19740 95172 19796 95174
rect 19820 95172 19876 95174
rect 4220 94682 4276 94684
rect 4300 94682 4356 94684
rect 4380 94682 4436 94684
rect 4460 94682 4516 94684
rect 4220 94630 4246 94682
rect 4246 94630 4276 94682
rect 4300 94630 4310 94682
rect 4310 94630 4356 94682
rect 4380 94630 4426 94682
rect 4426 94630 4436 94682
rect 4460 94630 4490 94682
rect 4490 94630 4516 94682
rect 4220 94628 4276 94630
rect 4300 94628 4356 94630
rect 4380 94628 4436 94630
rect 4460 94628 4516 94630
rect 19580 94138 19636 94140
rect 19660 94138 19716 94140
rect 19740 94138 19796 94140
rect 19820 94138 19876 94140
rect 19580 94086 19606 94138
rect 19606 94086 19636 94138
rect 19660 94086 19670 94138
rect 19670 94086 19716 94138
rect 19740 94086 19786 94138
rect 19786 94086 19796 94138
rect 19820 94086 19850 94138
rect 19850 94086 19876 94138
rect 19580 94084 19636 94086
rect 19660 94084 19716 94086
rect 19740 94084 19796 94086
rect 19820 94084 19876 94086
rect 4220 93594 4276 93596
rect 4300 93594 4356 93596
rect 4380 93594 4436 93596
rect 4460 93594 4516 93596
rect 4220 93542 4246 93594
rect 4246 93542 4276 93594
rect 4300 93542 4310 93594
rect 4310 93542 4356 93594
rect 4380 93542 4426 93594
rect 4426 93542 4436 93594
rect 4460 93542 4490 93594
rect 4490 93542 4516 93594
rect 4220 93540 4276 93542
rect 4300 93540 4356 93542
rect 4380 93540 4436 93542
rect 4460 93540 4516 93542
rect 19580 93050 19636 93052
rect 19660 93050 19716 93052
rect 19740 93050 19796 93052
rect 19820 93050 19876 93052
rect 19580 92998 19606 93050
rect 19606 92998 19636 93050
rect 19660 92998 19670 93050
rect 19670 92998 19716 93050
rect 19740 92998 19786 93050
rect 19786 92998 19796 93050
rect 19820 92998 19850 93050
rect 19850 92998 19876 93050
rect 19580 92996 19636 92998
rect 19660 92996 19716 92998
rect 19740 92996 19796 92998
rect 19820 92996 19876 92998
rect 4220 92506 4276 92508
rect 4300 92506 4356 92508
rect 4380 92506 4436 92508
rect 4460 92506 4516 92508
rect 4220 92454 4246 92506
rect 4246 92454 4276 92506
rect 4300 92454 4310 92506
rect 4310 92454 4356 92506
rect 4380 92454 4426 92506
rect 4426 92454 4436 92506
rect 4460 92454 4490 92506
rect 4490 92454 4516 92506
rect 4220 92452 4276 92454
rect 4300 92452 4356 92454
rect 4380 92452 4436 92454
rect 4460 92452 4516 92454
rect 19580 91962 19636 91964
rect 19660 91962 19716 91964
rect 19740 91962 19796 91964
rect 19820 91962 19876 91964
rect 19580 91910 19606 91962
rect 19606 91910 19636 91962
rect 19660 91910 19670 91962
rect 19670 91910 19716 91962
rect 19740 91910 19786 91962
rect 19786 91910 19796 91962
rect 19820 91910 19850 91962
rect 19850 91910 19876 91962
rect 19580 91908 19636 91910
rect 19660 91908 19716 91910
rect 19740 91908 19796 91910
rect 19820 91908 19876 91910
rect 4220 91418 4276 91420
rect 4300 91418 4356 91420
rect 4380 91418 4436 91420
rect 4460 91418 4516 91420
rect 4220 91366 4246 91418
rect 4246 91366 4276 91418
rect 4300 91366 4310 91418
rect 4310 91366 4356 91418
rect 4380 91366 4426 91418
rect 4426 91366 4436 91418
rect 4460 91366 4490 91418
rect 4490 91366 4516 91418
rect 4220 91364 4276 91366
rect 4300 91364 4356 91366
rect 4380 91364 4436 91366
rect 4460 91364 4516 91366
rect 19580 90874 19636 90876
rect 19660 90874 19716 90876
rect 19740 90874 19796 90876
rect 19820 90874 19876 90876
rect 19580 90822 19606 90874
rect 19606 90822 19636 90874
rect 19660 90822 19670 90874
rect 19670 90822 19716 90874
rect 19740 90822 19786 90874
rect 19786 90822 19796 90874
rect 19820 90822 19850 90874
rect 19850 90822 19876 90874
rect 19580 90820 19636 90822
rect 19660 90820 19716 90822
rect 19740 90820 19796 90822
rect 19820 90820 19876 90822
rect 4220 90330 4276 90332
rect 4300 90330 4356 90332
rect 4380 90330 4436 90332
rect 4460 90330 4516 90332
rect 4220 90278 4246 90330
rect 4246 90278 4276 90330
rect 4300 90278 4310 90330
rect 4310 90278 4356 90330
rect 4380 90278 4426 90330
rect 4426 90278 4436 90330
rect 4460 90278 4490 90330
rect 4490 90278 4516 90330
rect 4220 90276 4276 90278
rect 4300 90276 4356 90278
rect 4380 90276 4436 90278
rect 4460 90276 4516 90278
rect 19580 89786 19636 89788
rect 19660 89786 19716 89788
rect 19740 89786 19796 89788
rect 19820 89786 19876 89788
rect 19580 89734 19606 89786
rect 19606 89734 19636 89786
rect 19660 89734 19670 89786
rect 19670 89734 19716 89786
rect 19740 89734 19786 89786
rect 19786 89734 19796 89786
rect 19820 89734 19850 89786
rect 19850 89734 19876 89786
rect 19580 89732 19636 89734
rect 19660 89732 19716 89734
rect 19740 89732 19796 89734
rect 19820 89732 19876 89734
rect 4220 89242 4276 89244
rect 4300 89242 4356 89244
rect 4380 89242 4436 89244
rect 4460 89242 4516 89244
rect 4220 89190 4246 89242
rect 4246 89190 4276 89242
rect 4300 89190 4310 89242
rect 4310 89190 4356 89242
rect 4380 89190 4426 89242
rect 4426 89190 4436 89242
rect 4460 89190 4490 89242
rect 4490 89190 4516 89242
rect 4220 89188 4276 89190
rect 4300 89188 4356 89190
rect 4380 89188 4436 89190
rect 4460 89188 4516 89190
rect 19580 88698 19636 88700
rect 19660 88698 19716 88700
rect 19740 88698 19796 88700
rect 19820 88698 19876 88700
rect 19580 88646 19606 88698
rect 19606 88646 19636 88698
rect 19660 88646 19670 88698
rect 19670 88646 19716 88698
rect 19740 88646 19786 88698
rect 19786 88646 19796 88698
rect 19820 88646 19850 88698
rect 19850 88646 19876 88698
rect 19580 88644 19636 88646
rect 19660 88644 19716 88646
rect 19740 88644 19796 88646
rect 19820 88644 19876 88646
rect 4220 88154 4276 88156
rect 4300 88154 4356 88156
rect 4380 88154 4436 88156
rect 4460 88154 4516 88156
rect 4220 88102 4246 88154
rect 4246 88102 4276 88154
rect 4300 88102 4310 88154
rect 4310 88102 4356 88154
rect 4380 88102 4426 88154
rect 4426 88102 4436 88154
rect 4460 88102 4490 88154
rect 4490 88102 4516 88154
rect 4220 88100 4276 88102
rect 4300 88100 4356 88102
rect 4380 88100 4436 88102
rect 4460 88100 4516 88102
rect 19580 87610 19636 87612
rect 19660 87610 19716 87612
rect 19740 87610 19796 87612
rect 19820 87610 19876 87612
rect 19580 87558 19606 87610
rect 19606 87558 19636 87610
rect 19660 87558 19670 87610
rect 19670 87558 19716 87610
rect 19740 87558 19786 87610
rect 19786 87558 19796 87610
rect 19820 87558 19850 87610
rect 19850 87558 19876 87610
rect 19580 87556 19636 87558
rect 19660 87556 19716 87558
rect 19740 87556 19796 87558
rect 19820 87556 19876 87558
rect 4220 87066 4276 87068
rect 4300 87066 4356 87068
rect 4380 87066 4436 87068
rect 4460 87066 4516 87068
rect 4220 87014 4246 87066
rect 4246 87014 4276 87066
rect 4300 87014 4310 87066
rect 4310 87014 4356 87066
rect 4380 87014 4426 87066
rect 4426 87014 4436 87066
rect 4460 87014 4490 87066
rect 4490 87014 4516 87066
rect 4220 87012 4276 87014
rect 4300 87012 4356 87014
rect 4380 87012 4436 87014
rect 4460 87012 4516 87014
rect 19580 86522 19636 86524
rect 19660 86522 19716 86524
rect 19740 86522 19796 86524
rect 19820 86522 19876 86524
rect 19580 86470 19606 86522
rect 19606 86470 19636 86522
rect 19660 86470 19670 86522
rect 19670 86470 19716 86522
rect 19740 86470 19786 86522
rect 19786 86470 19796 86522
rect 19820 86470 19850 86522
rect 19850 86470 19876 86522
rect 19580 86468 19636 86470
rect 19660 86468 19716 86470
rect 19740 86468 19796 86470
rect 19820 86468 19876 86470
rect 4220 85978 4276 85980
rect 4300 85978 4356 85980
rect 4380 85978 4436 85980
rect 4460 85978 4516 85980
rect 4220 85926 4246 85978
rect 4246 85926 4276 85978
rect 4300 85926 4310 85978
rect 4310 85926 4356 85978
rect 4380 85926 4426 85978
rect 4426 85926 4436 85978
rect 4460 85926 4490 85978
rect 4490 85926 4516 85978
rect 4220 85924 4276 85926
rect 4300 85924 4356 85926
rect 4380 85924 4436 85926
rect 4460 85924 4516 85926
rect 19580 85434 19636 85436
rect 19660 85434 19716 85436
rect 19740 85434 19796 85436
rect 19820 85434 19876 85436
rect 19580 85382 19606 85434
rect 19606 85382 19636 85434
rect 19660 85382 19670 85434
rect 19670 85382 19716 85434
rect 19740 85382 19786 85434
rect 19786 85382 19796 85434
rect 19820 85382 19850 85434
rect 19850 85382 19876 85434
rect 19580 85380 19636 85382
rect 19660 85380 19716 85382
rect 19740 85380 19796 85382
rect 19820 85380 19876 85382
rect 4220 84890 4276 84892
rect 4300 84890 4356 84892
rect 4380 84890 4436 84892
rect 4460 84890 4516 84892
rect 4220 84838 4246 84890
rect 4246 84838 4276 84890
rect 4300 84838 4310 84890
rect 4310 84838 4356 84890
rect 4380 84838 4426 84890
rect 4426 84838 4436 84890
rect 4460 84838 4490 84890
rect 4490 84838 4516 84890
rect 4220 84836 4276 84838
rect 4300 84836 4356 84838
rect 4380 84836 4436 84838
rect 4460 84836 4516 84838
rect 19580 84346 19636 84348
rect 19660 84346 19716 84348
rect 19740 84346 19796 84348
rect 19820 84346 19876 84348
rect 19580 84294 19606 84346
rect 19606 84294 19636 84346
rect 19660 84294 19670 84346
rect 19670 84294 19716 84346
rect 19740 84294 19786 84346
rect 19786 84294 19796 84346
rect 19820 84294 19850 84346
rect 19850 84294 19876 84346
rect 19580 84292 19636 84294
rect 19660 84292 19716 84294
rect 19740 84292 19796 84294
rect 19820 84292 19876 84294
rect 4220 83802 4276 83804
rect 4300 83802 4356 83804
rect 4380 83802 4436 83804
rect 4460 83802 4516 83804
rect 4220 83750 4246 83802
rect 4246 83750 4276 83802
rect 4300 83750 4310 83802
rect 4310 83750 4356 83802
rect 4380 83750 4426 83802
rect 4426 83750 4436 83802
rect 4460 83750 4490 83802
rect 4490 83750 4516 83802
rect 4220 83748 4276 83750
rect 4300 83748 4356 83750
rect 4380 83748 4436 83750
rect 4460 83748 4516 83750
rect 19580 83258 19636 83260
rect 19660 83258 19716 83260
rect 19740 83258 19796 83260
rect 19820 83258 19876 83260
rect 19580 83206 19606 83258
rect 19606 83206 19636 83258
rect 19660 83206 19670 83258
rect 19670 83206 19716 83258
rect 19740 83206 19786 83258
rect 19786 83206 19796 83258
rect 19820 83206 19850 83258
rect 19850 83206 19876 83258
rect 19580 83204 19636 83206
rect 19660 83204 19716 83206
rect 19740 83204 19796 83206
rect 19820 83204 19876 83206
rect 4220 82714 4276 82716
rect 4300 82714 4356 82716
rect 4380 82714 4436 82716
rect 4460 82714 4516 82716
rect 4220 82662 4246 82714
rect 4246 82662 4276 82714
rect 4300 82662 4310 82714
rect 4310 82662 4356 82714
rect 4380 82662 4426 82714
rect 4426 82662 4436 82714
rect 4460 82662 4490 82714
rect 4490 82662 4516 82714
rect 4220 82660 4276 82662
rect 4300 82660 4356 82662
rect 4380 82660 4436 82662
rect 4460 82660 4516 82662
rect 19580 82170 19636 82172
rect 19660 82170 19716 82172
rect 19740 82170 19796 82172
rect 19820 82170 19876 82172
rect 19580 82118 19606 82170
rect 19606 82118 19636 82170
rect 19660 82118 19670 82170
rect 19670 82118 19716 82170
rect 19740 82118 19786 82170
rect 19786 82118 19796 82170
rect 19820 82118 19850 82170
rect 19850 82118 19876 82170
rect 19580 82116 19636 82118
rect 19660 82116 19716 82118
rect 19740 82116 19796 82118
rect 19820 82116 19876 82118
rect 4220 81626 4276 81628
rect 4300 81626 4356 81628
rect 4380 81626 4436 81628
rect 4460 81626 4516 81628
rect 4220 81574 4246 81626
rect 4246 81574 4276 81626
rect 4300 81574 4310 81626
rect 4310 81574 4356 81626
rect 4380 81574 4426 81626
rect 4426 81574 4436 81626
rect 4460 81574 4490 81626
rect 4490 81574 4516 81626
rect 4220 81572 4276 81574
rect 4300 81572 4356 81574
rect 4380 81572 4436 81574
rect 4460 81572 4516 81574
rect 19580 81082 19636 81084
rect 19660 81082 19716 81084
rect 19740 81082 19796 81084
rect 19820 81082 19876 81084
rect 19580 81030 19606 81082
rect 19606 81030 19636 81082
rect 19660 81030 19670 81082
rect 19670 81030 19716 81082
rect 19740 81030 19786 81082
rect 19786 81030 19796 81082
rect 19820 81030 19850 81082
rect 19850 81030 19876 81082
rect 19580 81028 19636 81030
rect 19660 81028 19716 81030
rect 19740 81028 19796 81030
rect 19820 81028 19876 81030
rect 4220 80538 4276 80540
rect 4300 80538 4356 80540
rect 4380 80538 4436 80540
rect 4460 80538 4516 80540
rect 4220 80486 4246 80538
rect 4246 80486 4276 80538
rect 4300 80486 4310 80538
rect 4310 80486 4356 80538
rect 4380 80486 4426 80538
rect 4426 80486 4436 80538
rect 4460 80486 4490 80538
rect 4490 80486 4516 80538
rect 4220 80484 4276 80486
rect 4300 80484 4356 80486
rect 4380 80484 4436 80486
rect 4460 80484 4516 80486
rect 19580 79994 19636 79996
rect 19660 79994 19716 79996
rect 19740 79994 19796 79996
rect 19820 79994 19876 79996
rect 19580 79942 19606 79994
rect 19606 79942 19636 79994
rect 19660 79942 19670 79994
rect 19670 79942 19716 79994
rect 19740 79942 19786 79994
rect 19786 79942 19796 79994
rect 19820 79942 19850 79994
rect 19850 79942 19876 79994
rect 19580 79940 19636 79942
rect 19660 79940 19716 79942
rect 19740 79940 19796 79942
rect 19820 79940 19876 79942
rect 4220 79450 4276 79452
rect 4300 79450 4356 79452
rect 4380 79450 4436 79452
rect 4460 79450 4516 79452
rect 4220 79398 4246 79450
rect 4246 79398 4276 79450
rect 4300 79398 4310 79450
rect 4310 79398 4356 79450
rect 4380 79398 4426 79450
rect 4426 79398 4436 79450
rect 4460 79398 4490 79450
rect 4490 79398 4516 79450
rect 4220 79396 4276 79398
rect 4300 79396 4356 79398
rect 4380 79396 4436 79398
rect 4460 79396 4516 79398
rect 19580 78906 19636 78908
rect 19660 78906 19716 78908
rect 19740 78906 19796 78908
rect 19820 78906 19876 78908
rect 19580 78854 19606 78906
rect 19606 78854 19636 78906
rect 19660 78854 19670 78906
rect 19670 78854 19716 78906
rect 19740 78854 19786 78906
rect 19786 78854 19796 78906
rect 19820 78854 19850 78906
rect 19850 78854 19876 78906
rect 19580 78852 19636 78854
rect 19660 78852 19716 78854
rect 19740 78852 19796 78854
rect 19820 78852 19876 78854
rect 4220 78362 4276 78364
rect 4300 78362 4356 78364
rect 4380 78362 4436 78364
rect 4460 78362 4516 78364
rect 4220 78310 4246 78362
rect 4246 78310 4276 78362
rect 4300 78310 4310 78362
rect 4310 78310 4356 78362
rect 4380 78310 4426 78362
rect 4426 78310 4436 78362
rect 4460 78310 4490 78362
rect 4490 78310 4516 78362
rect 4220 78308 4276 78310
rect 4300 78308 4356 78310
rect 4380 78308 4436 78310
rect 4460 78308 4516 78310
rect 19580 77818 19636 77820
rect 19660 77818 19716 77820
rect 19740 77818 19796 77820
rect 19820 77818 19876 77820
rect 19580 77766 19606 77818
rect 19606 77766 19636 77818
rect 19660 77766 19670 77818
rect 19670 77766 19716 77818
rect 19740 77766 19786 77818
rect 19786 77766 19796 77818
rect 19820 77766 19850 77818
rect 19850 77766 19876 77818
rect 19580 77764 19636 77766
rect 19660 77764 19716 77766
rect 19740 77764 19796 77766
rect 19820 77764 19876 77766
rect 4220 77274 4276 77276
rect 4300 77274 4356 77276
rect 4380 77274 4436 77276
rect 4460 77274 4516 77276
rect 4220 77222 4246 77274
rect 4246 77222 4276 77274
rect 4300 77222 4310 77274
rect 4310 77222 4356 77274
rect 4380 77222 4426 77274
rect 4426 77222 4436 77274
rect 4460 77222 4490 77274
rect 4490 77222 4516 77274
rect 4220 77220 4276 77222
rect 4300 77220 4356 77222
rect 4380 77220 4436 77222
rect 4460 77220 4516 77222
rect 19580 76730 19636 76732
rect 19660 76730 19716 76732
rect 19740 76730 19796 76732
rect 19820 76730 19876 76732
rect 19580 76678 19606 76730
rect 19606 76678 19636 76730
rect 19660 76678 19670 76730
rect 19670 76678 19716 76730
rect 19740 76678 19786 76730
rect 19786 76678 19796 76730
rect 19820 76678 19850 76730
rect 19850 76678 19876 76730
rect 19580 76676 19636 76678
rect 19660 76676 19716 76678
rect 19740 76676 19796 76678
rect 19820 76676 19876 76678
rect 4220 76186 4276 76188
rect 4300 76186 4356 76188
rect 4380 76186 4436 76188
rect 4460 76186 4516 76188
rect 4220 76134 4246 76186
rect 4246 76134 4276 76186
rect 4300 76134 4310 76186
rect 4310 76134 4356 76186
rect 4380 76134 4426 76186
rect 4426 76134 4436 76186
rect 4460 76134 4490 76186
rect 4490 76134 4516 76186
rect 4220 76132 4276 76134
rect 4300 76132 4356 76134
rect 4380 76132 4436 76134
rect 4460 76132 4516 76134
rect 19580 75642 19636 75644
rect 19660 75642 19716 75644
rect 19740 75642 19796 75644
rect 19820 75642 19876 75644
rect 19580 75590 19606 75642
rect 19606 75590 19636 75642
rect 19660 75590 19670 75642
rect 19670 75590 19716 75642
rect 19740 75590 19786 75642
rect 19786 75590 19796 75642
rect 19820 75590 19850 75642
rect 19850 75590 19876 75642
rect 19580 75588 19636 75590
rect 19660 75588 19716 75590
rect 19740 75588 19796 75590
rect 19820 75588 19876 75590
rect 4220 75098 4276 75100
rect 4300 75098 4356 75100
rect 4380 75098 4436 75100
rect 4460 75098 4516 75100
rect 4220 75046 4246 75098
rect 4246 75046 4276 75098
rect 4300 75046 4310 75098
rect 4310 75046 4356 75098
rect 4380 75046 4426 75098
rect 4426 75046 4436 75098
rect 4460 75046 4490 75098
rect 4490 75046 4516 75098
rect 4220 75044 4276 75046
rect 4300 75044 4356 75046
rect 4380 75044 4436 75046
rect 4460 75044 4516 75046
rect 19580 74554 19636 74556
rect 19660 74554 19716 74556
rect 19740 74554 19796 74556
rect 19820 74554 19876 74556
rect 19580 74502 19606 74554
rect 19606 74502 19636 74554
rect 19660 74502 19670 74554
rect 19670 74502 19716 74554
rect 19740 74502 19786 74554
rect 19786 74502 19796 74554
rect 19820 74502 19850 74554
rect 19850 74502 19876 74554
rect 19580 74500 19636 74502
rect 19660 74500 19716 74502
rect 19740 74500 19796 74502
rect 19820 74500 19876 74502
rect 4220 74010 4276 74012
rect 4300 74010 4356 74012
rect 4380 74010 4436 74012
rect 4460 74010 4516 74012
rect 4220 73958 4246 74010
rect 4246 73958 4276 74010
rect 4300 73958 4310 74010
rect 4310 73958 4356 74010
rect 4380 73958 4426 74010
rect 4426 73958 4436 74010
rect 4460 73958 4490 74010
rect 4490 73958 4516 74010
rect 4220 73956 4276 73958
rect 4300 73956 4356 73958
rect 4380 73956 4436 73958
rect 4460 73956 4516 73958
rect 19580 73466 19636 73468
rect 19660 73466 19716 73468
rect 19740 73466 19796 73468
rect 19820 73466 19876 73468
rect 19580 73414 19606 73466
rect 19606 73414 19636 73466
rect 19660 73414 19670 73466
rect 19670 73414 19716 73466
rect 19740 73414 19786 73466
rect 19786 73414 19796 73466
rect 19820 73414 19850 73466
rect 19850 73414 19876 73466
rect 19580 73412 19636 73414
rect 19660 73412 19716 73414
rect 19740 73412 19796 73414
rect 19820 73412 19876 73414
rect 4220 72922 4276 72924
rect 4300 72922 4356 72924
rect 4380 72922 4436 72924
rect 4460 72922 4516 72924
rect 4220 72870 4246 72922
rect 4246 72870 4276 72922
rect 4300 72870 4310 72922
rect 4310 72870 4356 72922
rect 4380 72870 4426 72922
rect 4426 72870 4436 72922
rect 4460 72870 4490 72922
rect 4490 72870 4516 72922
rect 4220 72868 4276 72870
rect 4300 72868 4356 72870
rect 4380 72868 4436 72870
rect 4460 72868 4516 72870
rect 19580 72378 19636 72380
rect 19660 72378 19716 72380
rect 19740 72378 19796 72380
rect 19820 72378 19876 72380
rect 19580 72326 19606 72378
rect 19606 72326 19636 72378
rect 19660 72326 19670 72378
rect 19670 72326 19716 72378
rect 19740 72326 19786 72378
rect 19786 72326 19796 72378
rect 19820 72326 19850 72378
rect 19850 72326 19876 72378
rect 19580 72324 19636 72326
rect 19660 72324 19716 72326
rect 19740 72324 19796 72326
rect 19820 72324 19876 72326
rect 4220 71834 4276 71836
rect 4300 71834 4356 71836
rect 4380 71834 4436 71836
rect 4460 71834 4516 71836
rect 4220 71782 4246 71834
rect 4246 71782 4276 71834
rect 4300 71782 4310 71834
rect 4310 71782 4356 71834
rect 4380 71782 4426 71834
rect 4426 71782 4436 71834
rect 4460 71782 4490 71834
rect 4490 71782 4516 71834
rect 4220 71780 4276 71782
rect 4300 71780 4356 71782
rect 4380 71780 4436 71782
rect 4460 71780 4516 71782
rect 19580 71290 19636 71292
rect 19660 71290 19716 71292
rect 19740 71290 19796 71292
rect 19820 71290 19876 71292
rect 19580 71238 19606 71290
rect 19606 71238 19636 71290
rect 19660 71238 19670 71290
rect 19670 71238 19716 71290
rect 19740 71238 19786 71290
rect 19786 71238 19796 71290
rect 19820 71238 19850 71290
rect 19850 71238 19876 71290
rect 19580 71236 19636 71238
rect 19660 71236 19716 71238
rect 19740 71236 19796 71238
rect 19820 71236 19876 71238
rect 4220 70746 4276 70748
rect 4300 70746 4356 70748
rect 4380 70746 4436 70748
rect 4460 70746 4516 70748
rect 4220 70694 4246 70746
rect 4246 70694 4276 70746
rect 4300 70694 4310 70746
rect 4310 70694 4356 70746
rect 4380 70694 4426 70746
rect 4426 70694 4436 70746
rect 4460 70694 4490 70746
rect 4490 70694 4516 70746
rect 4220 70692 4276 70694
rect 4300 70692 4356 70694
rect 4380 70692 4436 70694
rect 4460 70692 4516 70694
rect 19580 70202 19636 70204
rect 19660 70202 19716 70204
rect 19740 70202 19796 70204
rect 19820 70202 19876 70204
rect 19580 70150 19606 70202
rect 19606 70150 19636 70202
rect 19660 70150 19670 70202
rect 19670 70150 19716 70202
rect 19740 70150 19786 70202
rect 19786 70150 19796 70202
rect 19820 70150 19850 70202
rect 19850 70150 19876 70202
rect 19580 70148 19636 70150
rect 19660 70148 19716 70150
rect 19740 70148 19796 70150
rect 19820 70148 19876 70150
rect 4220 69658 4276 69660
rect 4300 69658 4356 69660
rect 4380 69658 4436 69660
rect 4460 69658 4516 69660
rect 4220 69606 4246 69658
rect 4246 69606 4276 69658
rect 4300 69606 4310 69658
rect 4310 69606 4356 69658
rect 4380 69606 4426 69658
rect 4426 69606 4436 69658
rect 4460 69606 4490 69658
rect 4490 69606 4516 69658
rect 4220 69604 4276 69606
rect 4300 69604 4356 69606
rect 4380 69604 4436 69606
rect 4460 69604 4516 69606
rect 19580 69114 19636 69116
rect 19660 69114 19716 69116
rect 19740 69114 19796 69116
rect 19820 69114 19876 69116
rect 19580 69062 19606 69114
rect 19606 69062 19636 69114
rect 19660 69062 19670 69114
rect 19670 69062 19716 69114
rect 19740 69062 19786 69114
rect 19786 69062 19796 69114
rect 19820 69062 19850 69114
rect 19850 69062 19876 69114
rect 19580 69060 19636 69062
rect 19660 69060 19716 69062
rect 19740 69060 19796 69062
rect 19820 69060 19876 69062
rect 4220 68570 4276 68572
rect 4300 68570 4356 68572
rect 4380 68570 4436 68572
rect 4460 68570 4516 68572
rect 4220 68518 4246 68570
rect 4246 68518 4276 68570
rect 4300 68518 4310 68570
rect 4310 68518 4356 68570
rect 4380 68518 4426 68570
rect 4426 68518 4436 68570
rect 4460 68518 4490 68570
rect 4490 68518 4516 68570
rect 4220 68516 4276 68518
rect 4300 68516 4356 68518
rect 4380 68516 4436 68518
rect 4460 68516 4516 68518
rect 19580 68026 19636 68028
rect 19660 68026 19716 68028
rect 19740 68026 19796 68028
rect 19820 68026 19876 68028
rect 19580 67974 19606 68026
rect 19606 67974 19636 68026
rect 19660 67974 19670 68026
rect 19670 67974 19716 68026
rect 19740 67974 19786 68026
rect 19786 67974 19796 68026
rect 19820 67974 19850 68026
rect 19850 67974 19876 68026
rect 19580 67972 19636 67974
rect 19660 67972 19716 67974
rect 19740 67972 19796 67974
rect 19820 67972 19876 67974
rect 4220 67482 4276 67484
rect 4300 67482 4356 67484
rect 4380 67482 4436 67484
rect 4460 67482 4516 67484
rect 4220 67430 4246 67482
rect 4246 67430 4276 67482
rect 4300 67430 4310 67482
rect 4310 67430 4356 67482
rect 4380 67430 4426 67482
rect 4426 67430 4436 67482
rect 4460 67430 4490 67482
rect 4490 67430 4516 67482
rect 4220 67428 4276 67430
rect 4300 67428 4356 67430
rect 4380 67428 4436 67430
rect 4460 67428 4516 67430
rect 19580 66938 19636 66940
rect 19660 66938 19716 66940
rect 19740 66938 19796 66940
rect 19820 66938 19876 66940
rect 19580 66886 19606 66938
rect 19606 66886 19636 66938
rect 19660 66886 19670 66938
rect 19670 66886 19716 66938
rect 19740 66886 19786 66938
rect 19786 66886 19796 66938
rect 19820 66886 19850 66938
rect 19850 66886 19876 66938
rect 19580 66884 19636 66886
rect 19660 66884 19716 66886
rect 19740 66884 19796 66886
rect 19820 66884 19876 66886
rect 4220 66394 4276 66396
rect 4300 66394 4356 66396
rect 4380 66394 4436 66396
rect 4460 66394 4516 66396
rect 4220 66342 4246 66394
rect 4246 66342 4276 66394
rect 4300 66342 4310 66394
rect 4310 66342 4356 66394
rect 4380 66342 4426 66394
rect 4426 66342 4436 66394
rect 4460 66342 4490 66394
rect 4490 66342 4516 66394
rect 4220 66340 4276 66342
rect 4300 66340 4356 66342
rect 4380 66340 4436 66342
rect 4460 66340 4516 66342
rect 19580 65850 19636 65852
rect 19660 65850 19716 65852
rect 19740 65850 19796 65852
rect 19820 65850 19876 65852
rect 19580 65798 19606 65850
rect 19606 65798 19636 65850
rect 19660 65798 19670 65850
rect 19670 65798 19716 65850
rect 19740 65798 19786 65850
rect 19786 65798 19796 65850
rect 19820 65798 19850 65850
rect 19850 65798 19876 65850
rect 19580 65796 19636 65798
rect 19660 65796 19716 65798
rect 19740 65796 19796 65798
rect 19820 65796 19876 65798
rect 4220 65306 4276 65308
rect 4300 65306 4356 65308
rect 4380 65306 4436 65308
rect 4460 65306 4516 65308
rect 4220 65254 4246 65306
rect 4246 65254 4276 65306
rect 4300 65254 4310 65306
rect 4310 65254 4356 65306
rect 4380 65254 4426 65306
rect 4426 65254 4436 65306
rect 4460 65254 4490 65306
rect 4490 65254 4516 65306
rect 4220 65252 4276 65254
rect 4300 65252 4356 65254
rect 4380 65252 4436 65254
rect 4460 65252 4516 65254
rect 19580 64762 19636 64764
rect 19660 64762 19716 64764
rect 19740 64762 19796 64764
rect 19820 64762 19876 64764
rect 19580 64710 19606 64762
rect 19606 64710 19636 64762
rect 19660 64710 19670 64762
rect 19670 64710 19716 64762
rect 19740 64710 19786 64762
rect 19786 64710 19796 64762
rect 19820 64710 19850 64762
rect 19850 64710 19876 64762
rect 19580 64708 19636 64710
rect 19660 64708 19716 64710
rect 19740 64708 19796 64710
rect 19820 64708 19876 64710
rect 4220 64218 4276 64220
rect 4300 64218 4356 64220
rect 4380 64218 4436 64220
rect 4460 64218 4516 64220
rect 4220 64166 4246 64218
rect 4246 64166 4276 64218
rect 4300 64166 4310 64218
rect 4310 64166 4356 64218
rect 4380 64166 4426 64218
rect 4426 64166 4436 64218
rect 4460 64166 4490 64218
rect 4490 64166 4516 64218
rect 4220 64164 4276 64166
rect 4300 64164 4356 64166
rect 4380 64164 4436 64166
rect 4460 64164 4516 64166
rect 19580 63674 19636 63676
rect 19660 63674 19716 63676
rect 19740 63674 19796 63676
rect 19820 63674 19876 63676
rect 19580 63622 19606 63674
rect 19606 63622 19636 63674
rect 19660 63622 19670 63674
rect 19670 63622 19716 63674
rect 19740 63622 19786 63674
rect 19786 63622 19796 63674
rect 19820 63622 19850 63674
rect 19850 63622 19876 63674
rect 19580 63620 19636 63622
rect 19660 63620 19716 63622
rect 19740 63620 19796 63622
rect 19820 63620 19876 63622
rect 4220 63130 4276 63132
rect 4300 63130 4356 63132
rect 4380 63130 4436 63132
rect 4460 63130 4516 63132
rect 4220 63078 4246 63130
rect 4246 63078 4276 63130
rect 4300 63078 4310 63130
rect 4310 63078 4356 63130
rect 4380 63078 4426 63130
rect 4426 63078 4436 63130
rect 4460 63078 4490 63130
rect 4490 63078 4516 63130
rect 4220 63076 4276 63078
rect 4300 63076 4356 63078
rect 4380 63076 4436 63078
rect 4460 63076 4516 63078
rect 19580 62586 19636 62588
rect 19660 62586 19716 62588
rect 19740 62586 19796 62588
rect 19820 62586 19876 62588
rect 19580 62534 19606 62586
rect 19606 62534 19636 62586
rect 19660 62534 19670 62586
rect 19670 62534 19716 62586
rect 19740 62534 19786 62586
rect 19786 62534 19796 62586
rect 19820 62534 19850 62586
rect 19850 62534 19876 62586
rect 19580 62532 19636 62534
rect 19660 62532 19716 62534
rect 19740 62532 19796 62534
rect 19820 62532 19876 62534
rect 4220 62042 4276 62044
rect 4300 62042 4356 62044
rect 4380 62042 4436 62044
rect 4460 62042 4516 62044
rect 4220 61990 4246 62042
rect 4246 61990 4276 62042
rect 4300 61990 4310 62042
rect 4310 61990 4356 62042
rect 4380 61990 4426 62042
rect 4426 61990 4436 62042
rect 4460 61990 4490 62042
rect 4490 61990 4516 62042
rect 4220 61988 4276 61990
rect 4300 61988 4356 61990
rect 4380 61988 4436 61990
rect 4460 61988 4516 61990
rect 19580 61498 19636 61500
rect 19660 61498 19716 61500
rect 19740 61498 19796 61500
rect 19820 61498 19876 61500
rect 19580 61446 19606 61498
rect 19606 61446 19636 61498
rect 19660 61446 19670 61498
rect 19670 61446 19716 61498
rect 19740 61446 19786 61498
rect 19786 61446 19796 61498
rect 19820 61446 19850 61498
rect 19850 61446 19876 61498
rect 19580 61444 19636 61446
rect 19660 61444 19716 61446
rect 19740 61444 19796 61446
rect 19820 61444 19876 61446
rect 4220 60954 4276 60956
rect 4300 60954 4356 60956
rect 4380 60954 4436 60956
rect 4460 60954 4516 60956
rect 4220 60902 4246 60954
rect 4246 60902 4276 60954
rect 4300 60902 4310 60954
rect 4310 60902 4356 60954
rect 4380 60902 4426 60954
rect 4426 60902 4436 60954
rect 4460 60902 4490 60954
rect 4490 60902 4516 60954
rect 4220 60900 4276 60902
rect 4300 60900 4356 60902
rect 4380 60900 4436 60902
rect 4460 60900 4516 60902
rect 19580 60410 19636 60412
rect 19660 60410 19716 60412
rect 19740 60410 19796 60412
rect 19820 60410 19876 60412
rect 19580 60358 19606 60410
rect 19606 60358 19636 60410
rect 19660 60358 19670 60410
rect 19670 60358 19716 60410
rect 19740 60358 19786 60410
rect 19786 60358 19796 60410
rect 19820 60358 19850 60410
rect 19850 60358 19876 60410
rect 19580 60356 19636 60358
rect 19660 60356 19716 60358
rect 19740 60356 19796 60358
rect 19820 60356 19876 60358
rect 2042 60036 2098 60072
rect 2042 60016 2044 60036
rect 2044 60016 2096 60036
rect 2096 60016 2098 60036
rect 4220 59866 4276 59868
rect 4300 59866 4356 59868
rect 4380 59866 4436 59868
rect 4460 59866 4516 59868
rect 4220 59814 4246 59866
rect 4246 59814 4276 59866
rect 4300 59814 4310 59866
rect 4310 59814 4356 59866
rect 4380 59814 4426 59866
rect 4426 59814 4436 59866
rect 4460 59814 4490 59866
rect 4490 59814 4516 59866
rect 4220 59812 4276 59814
rect 4300 59812 4356 59814
rect 4380 59812 4436 59814
rect 4460 59812 4516 59814
rect 19580 59322 19636 59324
rect 19660 59322 19716 59324
rect 19740 59322 19796 59324
rect 19820 59322 19876 59324
rect 19580 59270 19606 59322
rect 19606 59270 19636 59322
rect 19660 59270 19670 59322
rect 19670 59270 19716 59322
rect 19740 59270 19786 59322
rect 19786 59270 19796 59322
rect 19820 59270 19850 59322
rect 19850 59270 19876 59322
rect 19580 59268 19636 59270
rect 19660 59268 19716 59270
rect 19740 59268 19796 59270
rect 19820 59268 19876 59270
rect 4220 58778 4276 58780
rect 4300 58778 4356 58780
rect 4380 58778 4436 58780
rect 4460 58778 4516 58780
rect 4220 58726 4246 58778
rect 4246 58726 4276 58778
rect 4300 58726 4310 58778
rect 4310 58726 4356 58778
rect 4380 58726 4426 58778
rect 4426 58726 4436 58778
rect 4460 58726 4490 58778
rect 4490 58726 4516 58778
rect 4220 58724 4276 58726
rect 4300 58724 4356 58726
rect 4380 58724 4436 58726
rect 4460 58724 4516 58726
rect 19580 58234 19636 58236
rect 19660 58234 19716 58236
rect 19740 58234 19796 58236
rect 19820 58234 19876 58236
rect 19580 58182 19606 58234
rect 19606 58182 19636 58234
rect 19660 58182 19670 58234
rect 19670 58182 19716 58234
rect 19740 58182 19786 58234
rect 19786 58182 19796 58234
rect 19820 58182 19850 58234
rect 19850 58182 19876 58234
rect 19580 58180 19636 58182
rect 19660 58180 19716 58182
rect 19740 58180 19796 58182
rect 19820 58180 19876 58182
rect 4220 57690 4276 57692
rect 4300 57690 4356 57692
rect 4380 57690 4436 57692
rect 4460 57690 4516 57692
rect 4220 57638 4246 57690
rect 4246 57638 4276 57690
rect 4300 57638 4310 57690
rect 4310 57638 4356 57690
rect 4380 57638 4426 57690
rect 4426 57638 4436 57690
rect 4460 57638 4490 57690
rect 4490 57638 4516 57690
rect 4220 57636 4276 57638
rect 4300 57636 4356 57638
rect 4380 57636 4436 57638
rect 4460 57636 4516 57638
rect 19580 57146 19636 57148
rect 19660 57146 19716 57148
rect 19740 57146 19796 57148
rect 19820 57146 19876 57148
rect 19580 57094 19606 57146
rect 19606 57094 19636 57146
rect 19660 57094 19670 57146
rect 19670 57094 19716 57146
rect 19740 57094 19786 57146
rect 19786 57094 19796 57146
rect 19820 57094 19850 57146
rect 19850 57094 19876 57146
rect 19580 57092 19636 57094
rect 19660 57092 19716 57094
rect 19740 57092 19796 57094
rect 19820 57092 19876 57094
rect 4220 56602 4276 56604
rect 4300 56602 4356 56604
rect 4380 56602 4436 56604
rect 4460 56602 4516 56604
rect 4220 56550 4246 56602
rect 4246 56550 4276 56602
rect 4300 56550 4310 56602
rect 4310 56550 4356 56602
rect 4380 56550 4426 56602
rect 4426 56550 4436 56602
rect 4460 56550 4490 56602
rect 4490 56550 4516 56602
rect 4220 56548 4276 56550
rect 4300 56548 4356 56550
rect 4380 56548 4436 56550
rect 4460 56548 4516 56550
rect 19580 56058 19636 56060
rect 19660 56058 19716 56060
rect 19740 56058 19796 56060
rect 19820 56058 19876 56060
rect 19580 56006 19606 56058
rect 19606 56006 19636 56058
rect 19660 56006 19670 56058
rect 19670 56006 19716 56058
rect 19740 56006 19786 56058
rect 19786 56006 19796 56058
rect 19820 56006 19850 56058
rect 19850 56006 19876 56058
rect 19580 56004 19636 56006
rect 19660 56004 19716 56006
rect 19740 56004 19796 56006
rect 19820 56004 19876 56006
rect 4220 55514 4276 55516
rect 4300 55514 4356 55516
rect 4380 55514 4436 55516
rect 4460 55514 4516 55516
rect 4220 55462 4246 55514
rect 4246 55462 4276 55514
rect 4300 55462 4310 55514
rect 4310 55462 4356 55514
rect 4380 55462 4426 55514
rect 4426 55462 4436 55514
rect 4460 55462 4490 55514
rect 4490 55462 4516 55514
rect 4220 55460 4276 55462
rect 4300 55460 4356 55462
rect 4380 55460 4436 55462
rect 4460 55460 4516 55462
rect 19580 54970 19636 54972
rect 19660 54970 19716 54972
rect 19740 54970 19796 54972
rect 19820 54970 19876 54972
rect 19580 54918 19606 54970
rect 19606 54918 19636 54970
rect 19660 54918 19670 54970
rect 19670 54918 19716 54970
rect 19740 54918 19786 54970
rect 19786 54918 19796 54970
rect 19820 54918 19850 54970
rect 19850 54918 19876 54970
rect 19580 54916 19636 54918
rect 19660 54916 19716 54918
rect 19740 54916 19796 54918
rect 19820 54916 19876 54918
rect 4220 54426 4276 54428
rect 4300 54426 4356 54428
rect 4380 54426 4436 54428
rect 4460 54426 4516 54428
rect 4220 54374 4246 54426
rect 4246 54374 4276 54426
rect 4300 54374 4310 54426
rect 4310 54374 4356 54426
rect 4380 54374 4426 54426
rect 4426 54374 4436 54426
rect 4460 54374 4490 54426
rect 4490 54374 4516 54426
rect 4220 54372 4276 54374
rect 4300 54372 4356 54374
rect 4380 54372 4436 54374
rect 4460 54372 4516 54374
rect 19580 53882 19636 53884
rect 19660 53882 19716 53884
rect 19740 53882 19796 53884
rect 19820 53882 19876 53884
rect 19580 53830 19606 53882
rect 19606 53830 19636 53882
rect 19660 53830 19670 53882
rect 19670 53830 19716 53882
rect 19740 53830 19786 53882
rect 19786 53830 19796 53882
rect 19820 53830 19850 53882
rect 19850 53830 19876 53882
rect 19580 53828 19636 53830
rect 19660 53828 19716 53830
rect 19740 53828 19796 53830
rect 19820 53828 19876 53830
rect 4220 53338 4276 53340
rect 4300 53338 4356 53340
rect 4380 53338 4436 53340
rect 4460 53338 4516 53340
rect 4220 53286 4246 53338
rect 4246 53286 4276 53338
rect 4300 53286 4310 53338
rect 4310 53286 4356 53338
rect 4380 53286 4426 53338
rect 4426 53286 4436 53338
rect 4460 53286 4490 53338
rect 4490 53286 4516 53338
rect 4220 53284 4276 53286
rect 4300 53284 4356 53286
rect 4380 53284 4436 53286
rect 4460 53284 4516 53286
rect 19580 52794 19636 52796
rect 19660 52794 19716 52796
rect 19740 52794 19796 52796
rect 19820 52794 19876 52796
rect 19580 52742 19606 52794
rect 19606 52742 19636 52794
rect 19660 52742 19670 52794
rect 19670 52742 19716 52794
rect 19740 52742 19786 52794
rect 19786 52742 19796 52794
rect 19820 52742 19850 52794
rect 19850 52742 19876 52794
rect 19580 52740 19636 52742
rect 19660 52740 19716 52742
rect 19740 52740 19796 52742
rect 19820 52740 19876 52742
rect 4220 52250 4276 52252
rect 4300 52250 4356 52252
rect 4380 52250 4436 52252
rect 4460 52250 4516 52252
rect 4220 52198 4246 52250
rect 4246 52198 4276 52250
rect 4300 52198 4310 52250
rect 4310 52198 4356 52250
rect 4380 52198 4426 52250
rect 4426 52198 4436 52250
rect 4460 52198 4490 52250
rect 4490 52198 4516 52250
rect 4220 52196 4276 52198
rect 4300 52196 4356 52198
rect 4380 52196 4436 52198
rect 4460 52196 4516 52198
rect 19580 51706 19636 51708
rect 19660 51706 19716 51708
rect 19740 51706 19796 51708
rect 19820 51706 19876 51708
rect 19580 51654 19606 51706
rect 19606 51654 19636 51706
rect 19660 51654 19670 51706
rect 19670 51654 19716 51706
rect 19740 51654 19786 51706
rect 19786 51654 19796 51706
rect 19820 51654 19850 51706
rect 19850 51654 19876 51706
rect 19580 51652 19636 51654
rect 19660 51652 19716 51654
rect 19740 51652 19796 51654
rect 19820 51652 19876 51654
rect 4220 51162 4276 51164
rect 4300 51162 4356 51164
rect 4380 51162 4436 51164
rect 4460 51162 4516 51164
rect 4220 51110 4246 51162
rect 4246 51110 4276 51162
rect 4300 51110 4310 51162
rect 4310 51110 4356 51162
rect 4380 51110 4426 51162
rect 4426 51110 4436 51162
rect 4460 51110 4490 51162
rect 4490 51110 4516 51162
rect 4220 51108 4276 51110
rect 4300 51108 4356 51110
rect 4380 51108 4436 51110
rect 4460 51108 4516 51110
rect 19580 50618 19636 50620
rect 19660 50618 19716 50620
rect 19740 50618 19796 50620
rect 19820 50618 19876 50620
rect 19580 50566 19606 50618
rect 19606 50566 19636 50618
rect 19660 50566 19670 50618
rect 19670 50566 19716 50618
rect 19740 50566 19786 50618
rect 19786 50566 19796 50618
rect 19820 50566 19850 50618
rect 19850 50566 19876 50618
rect 19580 50564 19636 50566
rect 19660 50564 19716 50566
rect 19740 50564 19796 50566
rect 19820 50564 19876 50566
rect 4220 50074 4276 50076
rect 4300 50074 4356 50076
rect 4380 50074 4436 50076
rect 4460 50074 4516 50076
rect 4220 50022 4246 50074
rect 4246 50022 4276 50074
rect 4300 50022 4310 50074
rect 4310 50022 4356 50074
rect 4380 50022 4426 50074
rect 4426 50022 4436 50074
rect 4460 50022 4490 50074
rect 4490 50022 4516 50074
rect 4220 50020 4276 50022
rect 4300 50020 4356 50022
rect 4380 50020 4436 50022
rect 4460 50020 4516 50022
rect 19580 49530 19636 49532
rect 19660 49530 19716 49532
rect 19740 49530 19796 49532
rect 19820 49530 19876 49532
rect 19580 49478 19606 49530
rect 19606 49478 19636 49530
rect 19660 49478 19670 49530
rect 19670 49478 19716 49530
rect 19740 49478 19786 49530
rect 19786 49478 19796 49530
rect 19820 49478 19850 49530
rect 19850 49478 19876 49530
rect 19580 49476 19636 49478
rect 19660 49476 19716 49478
rect 19740 49476 19796 49478
rect 19820 49476 19876 49478
rect 4220 48986 4276 48988
rect 4300 48986 4356 48988
rect 4380 48986 4436 48988
rect 4460 48986 4516 48988
rect 4220 48934 4246 48986
rect 4246 48934 4276 48986
rect 4300 48934 4310 48986
rect 4310 48934 4356 48986
rect 4380 48934 4426 48986
rect 4426 48934 4436 48986
rect 4460 48934 4490 48986
rect 4490 48934 4516 48986
rect 4220 48932 4276 48934
rect 4300 48932 4356 48934
rect 4380 48932 4436 48934
rect 4460 48932 4516 48934
rect 19580 48442 19636 48444
rect 19660 48442 19716 48444
rect 19740 48442 19796 48444
rect 19820 48442 19876 48444
rect 19580 48390 19606 48442
rect 19606 48390 19636 48442
rect 19660 48390 19670 48442
rect 19670 48390 19716 48442
rect 19740 48390 19786 48442
rect 19786 48390 19796 48442
rect 19820 48390 19850 48442
rect 19850 48390 19876 48442
rect 19580 48388 19636 48390
rect 19660 48388 19716 48390
rect 19740 48388 19796 48390
rect 19820 48388 19876 48390
rect 4220 47898 4276 47900
rect 4300 47898 4356 47900
rect 4380 47898 4436 47900
rect 4460 47898 4516 47900
rect 4220 47846 4246 47898
rect 4246 47846 4276 47898
rect 4300 47846 4310 47898
rect 4310 47846 4356 47898
rect 4380 47846 4426 47898
rect 4426 47846 4436 47898
rect 4460 47846 4490 47898
rect 4490 47846 4516 47898
rect 4220 47844 4276 47846
rect 4300 47844 4356 47846
rect 4380 47844 4436 47846
rect 4460 47844 4516 47846
rect 19580 47354 19636 47356
rect 19660 47354 19716 47356
rect 19740 47354 19796 47356
rect 19820 47354 19876 47356
rect 19580 47302 19606 47354
rect 19606 47302 19636 47354
rect 19660 47302 19670 47354
rect 19670 47302 19716 47354
rect 19740 47302 19786 47354
rect 19786 47302 19796 47354
rect 19820 47302 19850 47354
rect 19850 47302 19876 47354
rect 19580 47300 19636 47302
rect 19660 47300 19716 47302
rect 19740 47300 19796 47302
rect 19820 47300 19876 47302
rect 4220 46810 4276 46812
rect 4300 46810 4356 46812
rect 4380 46810 4436 46812
rect 4460 46810 4516 46812
rect 4220 46758 4246 46810
rect 4246 46758 4276 46810
rect 4300 46758 4310 46810
rect 4310 46758 4356 46810
rect 4380 46758 4426 46810
rect 4426 46758 4436 46810
rect 4460 46758 4490 46810
rect 4490 46758 4516 46810
rect 4220 46756 4276 46758
rect 4300 46756 4356 46758
rect 4380 46756 4436 46758
rect 4460 46756 4516 46758
rect 19580 46266 19636 46268
rect 19660 46266 19716 46268
rect 19740 46266 19796 46268
rect 19820 46266 19876 46268
rect 19580 46214 19606 46266
rect 19606 46214 19636 46266
rect 19660 46214 19670 46266
rect 19670 46214 19716 46266
rect 19740 46214 19786 46266
rect 19786 46214 19796 46266
rect 19820 46214 19850 46266
rect 19850 46214 19876 46266
rect 19580 46212 19636 46214
rect 19660 46212 19716 46214
rect 19740 46212 19796 46214
rect 19820 46212 19876 46214
rect 4220 45722 4276 45724
rect 4300 45722 4356 45724
rect 4380 45722 4436 45724
rect 4460 45722 4516 45724
rect 4220 45670 4246 45722
rect 4246 45670 4276 45722
rect 4300 45670 4310 45722
rect 4310 45670 4356 45722
rect 4380 45670 4426 45722
rect 4426 45670 4436 45722
rect 4460 45670 4490 45722
rect 4490 45670 4516 45722
rect 4220 45668 4276 45670
rect 4300 45668 4356 45670
rect 4380 45668 4436 45670
rect 4460 45668 4516 45670
rect 19580 45178 19636 45180
rect 19660 45178 19716 45180
rect 19740 45178 19796 45180
rect 19820 45178 19876 45180
rect 19580 45126 19606 45178
rect 19606 45126 19636 45178
rect 19660 45126 19670 45178
rect 19670 45126 19716 45178
rect 19740 45126 19786 45178
rect 19786 45126 19796 45178
rect 19820 45126 19850 45178
rect 19850 45126 19876 45178
rect 19580 45124 19636 45126
rect 19660 45124 19716 45126
rect 19740 45124 19796 45126
rect 19820 45124 19876 45126
rect 4220 44634 4276 44636
rect 4300 44634 4356 44636
rect 4380 44634 4436 44636
rect 4460 44634 4516 44636
rect 4220 44582 4246 44634
rect 4246 44582 4276 44634
rect 4300 44582 4310 44634
rect 4310 44582 4356 44634
rect 4380 44582 4426 44634
rect 4426 44582 4436 44634
rect 4460 44582 4490 44634
rect 4490 44582 4516 44634
rect 4220 44580 4276 44582
rect 4300 44580 4356 44582
rect 4380 44580 4436 44582
rect 4460 44580 4516 44582
rect 19580 44090 19636 44092
rect 19660 44090 19716 44092
rect 19740 44090 19796 44092
rect 19820 44090 19876 44092
rect 19580 44038 19606 44090
rect 19606 44038 19636 44090
rect 19660 44038 19670 44090
rect 19670 44038 19716 44090
rect 19740 44038 19786 44090
rect 19786 44038 19796 44090
rect 19820 44038 19850 44090
rect 19850 44038 19876 44090
rect 19580 44036 19636 44038
rect 19660 44036 19716 44038
rect 19740 44036 19796 44038
rect 19820 44036 19876 44038
rect 4220 43546 4276 43548
rect 4300 43546 4356 43548
rect 4380 43546 4436 43548
rect 4460 43546 4516 43548
rect 4220 43494 4246 43546
rect 4246 43494 4276 43546
rect 4300 43494 4310 43546
rect 4310 43494 4356 43546
rect 4380 43494 4426 43546
rect 4426 43494 4436 43546
rect 4460 43494 4490 43546
rect 4490 43494 4516 43546
rect 4220 43492 4276 43494
rect 4300 43492 4356 43494
rect 4380 43492 4436 43494
rect 4460 43492 4516 43494
rect 19580 43002 19636 43004
rect 19660 43002 19716 43004
rect 19740 43002 19796 43004
rect 19820 43002 19876 43004
rect 19580 42950 19606 43002
rect 19606 42950 19636 43002
rect 19660 42950 19670 43002
rect 19670 42950 19716 43002
rect 19740 42950 19786 43002
rect 19786 42950 19796 43002
rect 19820 42950 19850 43002
rect 19850 42950 19876 43002
rect 19580 42948 19636 42950
rect 19660 42948 19716 42950
rect 19740 42948 19796 42950
rect 19820 42948 19876 42950
rect 4220 42458 4276 42460
rect 4300 42458 4356 42460
rect 4380 42458 4436 42460
rect 4460 42458 4516 42460
rect 4220 42406 4246 42458
rect 4246 42406 4276 42458
rect 4300 42406 4310 42458
rect 4310 42406 4356 42458
rect 4380 42406 4426 42458
rect 4426 42406 4436 42458
rect 4460 42406 4490 42458
rect 4490 42406 4516 42458
rect 4220 42404 4276 42406
rect 4300 42404 4356 42406
rect 4380 42404 4436 42406
rect 4460 42404 4516 42406
rect 19580 41914 19636 41916
rect 19660 41914 19716 41916
rect 19740 41914 19796 41916
rect 19820 41914 19876 41916
rect 19580 41862 19606 41914
rect 19606 41862 19636 41914
rect 19660 41862 19670 41914
rect 19670 41862 19716 41914
rect 19740 41862 19786 41914
rect 19786 41862 19796 41914
rect 19820 41862 19850 41914
rect 19850 41862 19876 41914
rect 19580 41860 19636 41862
rect 19660 41860 19716 41862
rect 19740 41860 19796 41862
rect 19820 41860 19876 41862
rect 4220 41370 4276 41372
rect 4300 41370 4356 41372
rect 4380 41370 4436 41372
rect 4460 41370 4516 41372
rect 4220 41318 4246 41370
rect 4246 41318 4276 41370
rect 4300 41318 4310 41370
rect 4310 41318 4356 41370
rect 4380 41318 4426 41370
rect 4426 41318 4436 41370
rect 4460 41318 4490 41370
rect 4490 41318 4516 41370
rect 4220 41316 4276 41318
rect 4300 41316 4356 41318
rect 4380 41316 4436 41318
rect 4460 41316 4516 41318
rect 19580 40826 19636 40828
rect 19660 40826 19716 40828
rect 19740 40826 19796 40828
rect 19820 40826 19876 40828
rect 19580 40774 19606 40826
rect 19606 40774 19636 40826
rect 19660 40774 19670 40826
rect 19670 40774 19716 40826
rect 19740 40774 19786 40826
rect 19786 40774 19796 40826
rect 19820 40774 19850 40826
rect 19850 40774 19876 40826
rect 19580 40772 19636 40774
rect 19660 40772 19716 40774
rect 19740 40772 19796 40774
rect 19820 40772 19876 40774
rect 4220 40282 4276 40284
rect 4300 40282 4356 40284
rect 4380 40282 4436 40284
rect 4460 40282 4516 40284
rect 4220 40230 4246 40282
rect 4246 40230 4276 40282
rect 4300 40230 4310 40282
rect 4310 40230 4356 40282
rect 4380 40230 4426 40282
rect 4426 40230 4436 40282
rect 4460 40230 4490 40282
rect 4490 40230 4516 40282
rect 4220 40228 4276 40230
rect 4300 40228 4356 40230
rect 4380 40228 4436 40230
rect 4460 40228 4516 40230
rect 19580 39738 19636 39740
rect 19660 39738 19716 39740
rect 19740 39738 19796 39740
rect 19820 39738 19876 39740
rect 19580 39686 19606 39738
rect 19606 39686 19636 39738
rect 19660 39686 19670 39738
rect 19670 39686 19716 39738
rect 19740 39686 19786 39738
rect 19786 39686 19796 39738
rect 19820 39686 19850 39738
rect 19850 39686 19876 39738
rect 19580 39684 19636 39686
rect 19660 39684 19716 39686
rect 19740 39684 19796 39686
rect 19820 39684 19876 39686
rect 4220 39194 4276 39196
rect 4300 39194 4356 39196
rect 4380 39194 4436 39196
rect 4460 39194 4516 39196
rect 4220 39142 4246 39194
rect 4246 39142 4276 39194
rect 4300 39142 4310 39194
rect 4310 39142 4356 39194
rect 4380 39142 4426 39194
rect 4426 39142 4436 39194
rect 4460 39142 4490 39194
rect 4490 39142 4516 39194
rect 4220 39140 4276 39142
rect 4300 39140 4356 39142
rect 4380 39140 4436 39142
rect 4460 39140 4516 39142
rect 19580 38650 19636 38652
rect 19660 38650 19716 38652
rect 19740 38650 19796 38652
rect 19820 38650 19876 38652
rect 19580 38598 19606 38650
rect 19606 38598 19636 38650
rect 19660 38598 19670 38650
rect 19670 38598 19716 38650
rect 19740 38598 19786 38650
rect 19786 38598 19796 38650
rect 19820 38598 19850 38650
rect 19850 38598 19876 38650
rect 19580 38596 19636 38598
rect 19660 38596 19716 38598
rect 19740 38596 19796 38598
rect 19820 38596 19876 38598
rect 4220 38106 4276 38108
rect 4300 38106 4356 38108
rect 4380 38106 4436 38108
rect 4460 38106 4516 38108
rect 4220 38054 4246 38106
rect 4246 38054 4276 38106
rect 4300 38054 4310 38106
rect 4310 38054 4356 38106
rect 4380 38054 4426 38106
rect 4426 38054 4436 38106
rect 4460 38054 4490 38106
rect 4490 38054 4516 38106
rect 4220 38052 4276 38054
rect 4300 38052 4356 38054
rect 4380 38052 4436 38054
rect 4460 38052 4516 38054
rect 19580 37562 19636 37564
rect 19660 37562 19716 37564
rect 19740 37562 19796 37564
rect 19820 37562 19876 37564
rect 19580 37510 19606 37562
rect 19606 37510 19636 37562
rect 19660 37510 19670 37562
rect 19670 37510 19716 37562
rect 19740 37510 19786 37562
rect 19786 37510 19796 37562
rect 19820 37510 19850 37562
rect 19850 37510 19876 37562
rect 19580 37508 19636 37510
rect 19660 37508 19716 37510
rect 19740 37508 19796 37510
rect 19820 37508 19876 37510
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4246 37018
rect 4246 36966 4276 37018
rect 4300 36966 4310 37018
rect 4310 36966 4356 37018
rect 4380 36966 4426 37018
rect 4426 36966 4436 37018
rect 4460 36966 4490 37018
rect 4490 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 19580 36474 19636 36476
rect 19660 36474 19716 36476
rect 19740 36474 19796 36476
rect 19820 36474 19876 36476
rect 19580 36422 19606 36474
rect 19606 36422 19636 36474
rect 19660 36422 19670 36474
rect 19670 36422 19716 36474
rect 19740 36422 19786 36474
rect 19786 36422 19796 36474
rect 19820 36422 19850 36474
rect 19850 36422 19876 36474
rect 19580 36420 19636 36422
rect 19660 36420 19716 36422
rect 19740 36420 19796 36422
rect 19820 36420 19876 36422
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4246 35930
rect 4246 35878 4276 35930
rect 4300 35878 4310 35930
rect 4310 35878 4356 35930
rect 4380 35878 4426 35930
rect 4426 35878 4436 35930
rect 4460 35878 4490 35930
rect 4490 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 19580 35386 19636 35388
rect 19660 35386 19716 35388
rect 19740 35386 19796 35388
rect 19820 35386 19876 35388
rect 19580 35334 19606 35386
rect 19606 35334 19636 35386
rect 19660 35334 19670 35386
rect 19670 35334 19716 35386
rect 19740 35334 19786 35386
rect 19786 35334 19796 35386
rect 19820 35334 19850 35386
rect 19850 35334 19876 35386
rect 19580 35332 19636 35334
rect 19660 35332 19716 35334
rect 19740 35332 19796 35334
rect 19820 35332 19876 35334
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4246 34842
rect 4246 34790 4276 34842
rect 4300 34790 4310 34842
rect 4310 34790 4356 34842
rect 4380 34790 4426 34842
rect 4426 34790 4436 34842
rect 4460 34790 4490 34842
rect 4490 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 19580 34298 19636 34300
rect 19660 34298 19716 34300
rect 19740 34298 19796 34300
rect 19820 34298 19876 34300
rect 19580 34246 19606 34298
rect 19606 34246 19636 34298
rect 19660 34246 19670 34298
rect 19670 34246 19716 34298
rect 19740 34246 19786 34298
rect 19786 34246 19796 34298
rect 19820 34246 19850 34298
rect 19850 34246 19876 34298
rect 19580 34244 19636 34246
rect 19660 34244 19716 34246
rect 19740 34244 19796 34246
rect 19820 34244 19876 34246
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4246 33754
rect 4246 33702 4276 33754
rect 4300 33702 4310 33754
rect 4310 33702 4356 33754
rect 4380 33702 4426 33754
rect 4426 33702 4436 33754
rect 4460 33702 4490 33754
rect 4490 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 19580 33210 19636 33212
rect 19660 33210 19716 33212
rect 19740 33210 19796 33212
rect 19820 33210 19876 33212
rect 19580 33158 19606 33210
rect 19606 33158 19636 33210
rect 19660 33158 19670 33210
rect 19670 33158 19716 33210
rect 19740 33158 19786 33210
rect 19786 33158 19796 33210
rect 19820 33158 19850 33210
rect 19850 33158 19876 33210
rect 19580 33156 19636 33158
rect 19660 33156 19716 33158
rect 19740 33156 19796 33158
rect 19820 33156 19876 33158
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4246 32666
rect 4246 32614 4276 32666
rect 4300 32614 4310 32666
rect 4310 32614 4356 32666
rect 4380 32614 4426 32666
rect 4426 32614 4436 32666
rect 4460 32614 4490 32666
rect 4490 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 19580 32122 19636 32124
rect 19660 32122 19716 32124
rect 19740 32122 19796 32124
rect 19820 32122 19876 32124
rect 19580 32070 19606 32122
rect 19606 32070 19636 32122
rect 19660 32070 19670 32122
rect 19670 32070 19716 32122
rect 19740 32070 19786 32122
rect 19786 32070 19796 32122
rect 19820 32070 19850 32122
rect 19850 32070 19876 32122
rect 19580 32068 19636 32070
rect 19660 32068 19716 32070
rect 19740 32068 19796 32070
rect 19820 32068 19876 32070
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4246 31578
rect 4246 31526 4276 31578
rect 4300 31526 4310 31578
rect 4310 31526 4356 31578
rect 4380 31526 4426 31578
rect 4426 31526 4436 31578
rect 4460 31526 4490 31578
rect 4490 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 19580 31034 19636 31036
rect 19660 31034 19716 31036
rect 19740 31034 19796 31036
rect 19820 31034 19876 31036
rect 19580 30982 19606 31034
rect 19606 30982 19636 31034
rect 19660 30982 19670 31034
rect 19670 30982 19716 31034
rect 19740 30982 19786 31034
rect 19786 30982 19796 31034
rect 19820 30982 19850 31034
rect 19850 30982 19876 31034
rect 19580 30980 19636 30982
rect 19660 30980 19716 30982
rect 19740 30980 19796 30982
rect 19820 30980 19876 30982
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4246 30490
rect 4246 30438 4276 30490
rect 4300 30438 4310 30490
rect 4310 30438 4356 30490
rect 4380 30438 4426 30490
rect 4426 30438 4436 30490
rect 4460 30438 4490 30490
rect 4490 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 19580 29946 19636 29948
rect 19660 29946 19716 29948
rect 19740 29946 19796 29948
rect 19820 29946 19876 29948
rect 19580 29894 19606 29946
rect 19606 29894 19636 29946
rect 19660 29894 19670 29946
rect 19670 29894 19716 29946
rect 19740 29894 19786 29946
rect 19786 29894 19796 29946
rect 19820 29894 19850 29946
rect 19850 29894 19876 29946
rect 19580 29892 19636 29894
rect 19660 29892 19716 29894
rect 19740 29892 19796 29894
rect 19820 29892 19876 29894
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4246 29402
rect 4246 29350 4276 29402
rect 4300 29350 4310 29402
rect 4310 29350 4356 29402
rect 4380 29350 4426 29402
rect 4426 29350 4436 29402
rect 4460 29350 4490 29402
rect 4490 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 19580 28858 19636 28860
rect 19660 28858 19716 28860
rect 19740 28858 19796 28860
rect 19820 28858 19876 28860
rect 19580 28806 19606 28858
rect 19606 28806 19636 28858
rect 19660 28806 19670 28858
rect 19670 28806 19716 28858
rect 19740 28806 19786 28858
rect 19786 28806 19796 28858
rect 19820 28806 19850 28858
rect 19850 28806 19876 28858
rect 19580 28804 19636 28806
rect 19660 28804 19716 28806
rect 19740 28804 19796 28806
rect 19820 28804 19876 28806
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4246 28314
rect 4246 28262 4276 28314
rect 4300 28262 4310 28314
rect 4310 28262 4356 28314
rect 4380 28262 4426 28314
rect 4426 28262 4436 28314
rect 4460 28262 4490 28314
rect 4490 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 19580 27770 19636 27772
rect 19660 27770 19716 27772
rect 19740 27770 19796 27772
rect 19820 27770 19876 27772
rect 19580 27718 19606 27770
rect 19606 27718 19636 27770
rect 19660 27718 19670 27770
rect 19670 27718 19716 27770
rect 19740 27718 19786 27770
rect 19786 27718 19796 27770
rect 19820 27718 19850 27770
rect 19850 27718 19876 27770
rect 19580 27716 19636 27718
rect 19660 27716 19716 27718
rect 19740 27716 19796 27718
rect 19820 27716 19876 27718
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4246 27226
rect 4246 27174 4276 27226
rect 4300 27174 4310 27226
rect 4310 27174 4356 27226
rect 4380 27174 4426 27226
rect 4426 27174 4436 27226
rect 4460 27174 4490 27226
rect 4490 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 19580 26682 19636 26684
rect 19660 26682 19716 26684
rect 19740 26682 19796 26684
rect 19820 26682 19876 26684
rect 19580 26630 19606 26682
rect 19606 26630 19636 26682
rect 19660 26630 19670 26682
rect 19670 26630 19716 26682
rect 19740 26630 19786 26682
rect 19786 26630 19796 26682
rect 19820 26630 19850 26682
rect 19850 26630 19876 26682
rect 19580 26628 19636 26630
rect 19660 26628 19716 26630
rect 19740 26628 19796 26630
rect 19820 26628 19876 26630
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4246 26138
rect 4246 26086 4276 26138
rect 4300 26086 4310 26138
rect 4310 26086 4356 26138
rect 4380 26086 4426 26138
rect 4426 26086 4436 26138
rect 4460 26086 4490 26138
rect 4490 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 19580 25594 19636 25596
rect 19660 25594 19716 25596
rect 19740 25594 19796 25596
rect 19820 25594 19876 25596
rect 19580 25542 19606 25594
rect 19606 25542 19636 25594
rect 19660 25542 19670 25594
rect 19670 25542 19716 25594
rect 19740 25542 19786 25594
rect 19786 25542 19796 25594
rect 19820 25542 19850 25594
rect 19850 25542 19876 25594
rect 19580 25540 19636 25542
rect 19660 25540 19716 25542
rect 19740 25540 19796 25542
rect 19820 25540 19876 25542
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 19580 24506 19636 24508
rect 19660 24506 19716 24508
rect 19740 24506 19796 24508
rect 19820 24506 19876 24508
rect 19580 24454 19606 24506
rect 19606 24454 19636 24506
rect 19660 24454 19670 24506
rect 19670 24454 19716 24506
rect 19740 24454 19786 24506
rect 19786 24454 19796 24506
rect 19820 24454 19850 24506
rect 19850 24454 19876 24506
rect 19580 24452 19636 24454
rect 19660 24452 19716 24454
rect 19740 24452 19796 24454
rect 19820 24452 19876 24454
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 19580 23418 19636 23420
rect 19660 23418 19716 23420
rect 19740 23418 19796 23420
rect 19820 23418 19876 23420
rect 19580 23366 19606 23418
rect 19606 23366 19636 23418
rect 19660 23366 19670 23418
rect 19670 23366 19716 23418
rect 19740 23366 19786 23418
rect 19786 23366 19796 23418
rect 19820 23366 19850 23418
rect 19850 23366 19876 23418
rect 19580 23364 19636 23366
rect 19660 23364 19716 23366
rect 19740 23364 19796 23366
rect 19820 23364 19876 23366
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 19580 22330 19636 22332
rect 19660 22330 19716 22332
rect 19740 22330 19796 22332
rect 19820 22330 19876 22332
rect 19580 22278 19606 22330
rect 19606 22278 19636 22330
rect 19660 22278 19670 22330
rect 19670 22278 19716 22330
rect 19740 22278 19786 22330
rect 19786 22278 19796 22330
rect 19820 22278 19850 22330
rect 19850 22278 19876 22330
rect 19580 22276 19636 22278
rect 19660 22276 19716 22278
rect 19740 22276 19796 22278
rect 19820 22276 19876 22278
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 19580 21242 19636 21244
rect 19660 21242 19716 21244
rect 19740 21242 19796 21244
rect 19820 21242 19876 21244
rect 19580 21190 19606 21242
rect 19606 21190 19636 21242
rect 19660 21190 19670 21242
rect 19670 21190 19716 21242
rect 19740 21190 19786 21242
rect 19786 21190 19796 21242
rect 19820 21190 19850 21242
rect 19850 21190 19876 21242
rect 19580 21188 19636 21190
rect 19660 21188 19716 21190
rect 19740 21188 19796 21190
rect 19820 21188 19876 21190
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 19580 20154 19636 20156
rect 19660 20154 19716 20156
rect 19740 20154 19796 20156
rect 19820 20154 19876 20156
rect 19580 20102 19606 20154
rect 19606 20102 19636 20154
rect 19660 20102 19670 20154
rect 19670 20102 19716 20154
rect 19740 20102 19786 20154
rect 19786 20102 19796 20154
rect 19820 20102 19850 20154
rect 19850 20102 19876 20154
rect 19580 20100 19636 20102
rect 19660 20100 19716 20102
rect 19740 20100 19796 20102
rect 19820 20100 19876 20102
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 19580 19066 19636 19068
rect 19660 19066 19716 19068
rect 19740 19066 19796 19068
rect 19820 19066 19876 19068
rect 19580 19014 19606 19066
rect 19606 19014 19636 19066
rect 19660 19014 19670 19066
rect 19670 19014 19716 19066
rect 19740 19014 19786 19066
rect 19786 19014 19796 19066
rect 19820 19014 19850 19066
rect 19850 19014 19876 19066
rect 19580 19012 19636 19014
rect 19660 19012 19716 19014
rect 19740 19012 19796 19014
rect 19820 19012 19876 19014
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 19580 17978 19636 17980
rect 19660 17978 19716 17980
rect 19740 17978 19796 17980
rect 19820 17978 19876 17980
rect 19580 17926 19606 17978
rect 19606 17926 19636 17978
rect 19660 17926 19670 17978
rect 19670 17926 19716 17978
rect 19740 17926 19786 17978
rect 19786 17926 19796 17978
rect 19820 17926 19850 17978
rect 19850 17926 19876 17978
rect 19580 17924 19636 17926
rect 19660 17924 19716 17926
rect 19740 17924 19796 17926
rect 19820 17924 19876 17926
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 19580 16890 19636 16892
rect 19660 16890 19716 16892
rect 19740 16890 19796 16892
rect 19820 16890 19876 16892
rect 19580 16838 19606 16890
rect 19606 16838 19636 16890
rect 19660 16838 19670 16890
rect 19670 16838 19716 16890
rect 19740 16838 19786 16890
rect 19786 16838 19796 16890
rect 19820 16838 19850 16890
rect 19850 16838 19876 16890
rect 19580 16836 19636 16838
rect 19660 16836 19716 16838
rect 19740 16836 19796 16838
rect 19820 16836 19876 16838
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 19580 15802 19636 15804
rect 19660 15802 19716 15804
rect 19740 15802 19796 15804
rect 19820 15802 19876 15804
rect 19580 15750 19606 15802
rect 19606 15750 19636 15802
rect 19660 15750 19670 15802
rect 19670 15750 19716 15802
rect 19740 15750 19786 15802
rect 19786 15750 19796 15802
rect 19820 15750 19850 15802
rect 19850 15750 19876 15802
rect 19580 15748 19636 15750
rect 19660 15748 19716 15750
rect 19740 15748 19796 15750
rect 19820 15748 19876 15750
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 19580 14714 19636 14716
rect 19660 14714 19716 14716
rect 19740 14714 19796 14716
rect 19820 14714 19876 14716
rect 19580 14662 19606 14714
rect 19606 14662 19636 14714
rect 19660 14662 19670 14714
rect 19670 14662 19716 14714
rect 19740 14662 19786 14714
rect 19786 14662 19796 14714
rect 19820 14662 19850 14714
rect 19850 14662 19876 14714
rect 19580 14660 19636 14662
rect 19660 14660 19716 14662
rect 19740 14660 19796 14662
rect 19820 14660 19876 14662
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 19580 13626 19636 13628
rect 19660 13626 19716 13628
rect 19740 13626 19796 13628
rect 19820 13626 19876 13628
rect 19580 13574 19606 13626
rect 19606 13574 19636 13626
rect 19660 13574 19670 13626
rect 19670 13574 19716 13626
rect 19740 13574 19786 13626
rect 19786 13574 19796 13626
rect 19820 13574 19850 13626
rect 19850 13574 19876 13626
rect 19580 13572 19636 13574
rect 19660 13572 19716 13574
rect 19740 13572 19796 13574
rect 19820 13572 19876 13574
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 19580 12538 19636 12540
rect 19660 12538 19716 12540
rect 19740 12538 19796 12540
rect 19820 12538 19876 12540
rect 19580 12486 19606 12538
rect 19606 12486 19636 12538
rect 19660 12486 19670 12538
rect 19670 12486 19716 12538
rect 19740 12486 19786 12538
rect 19786 12486 19796 12538
rect 19820 12486 19850 12538
rect 19850 12486 19876 12538
rect 19580 12484 19636 12486
rect 19660 12484 19716 12486
rect 19740 12484 19796 12486
rect 19820 12484 19876 12486
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 19580 11450 19636 11452
rect 19660 11450 19716 11452
rect 19740 11450 19796 11452
rect 19820 11450 19876 11452
rect 19580 11398 19606 11450
rect 19606 11398 19636 11450
rect 19660 11398 19670 11450
rect 19670 11398 19716 11450
rect 19740 11398 19786 11450
rect 19786 11398 19796 11450
rect 19820 11398 19850 11450
rect 19850 11398 19876 11450
rect 19580 11396 19636 11398
rect 19660 11396 19716 11398
rect 19740 11396 19796 11398
rect 19820 11396 19876 11398
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 19580 10362 19636 10364
rect 19660 10362 19716 10364
rect 19740 10362 19796 10364
rect 19820 10362 19876 10364
rect 19580 10310 19606 10362
rect 19606 10310 19636 10362
rect 19660 10310 19670 10362
rect 19670 10310 19716 10362
rect 19740 10310 19786 10362
rect 19786 10310 19796 10362
rect 19820 10310 19850 10362
rect 19850 10310 19876 10362
rect 19580 10308 19636 10310
rect 19660 10308 19716 10310
rect 19740 10308 19796 10310
rect 19820 10308 19876 10310
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 19580 9274 19636 9276
rect 19660 9274 19716 9276
rect 19740 9274 19796 9276
rect 19820 9274 19876 9276
rect 19580 9222 19606 9274
rect 19606 9222 19636 9274
rect 19660 9222 19670 9274
rect 19670 9222 19716 9274
rect 19740 9222 19786 9274
rect 19786 9222 19796 9274
rect 19820 9222 19850 9274
rect 19850 9222 19876 9274
rect 19580 9220 19636 9222
rect 19660 9220 19716 9222
rect 19740 9220 19796 9222
rect 19820 9220 19876 9222
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 19580 8186 19636 8188
rect 19660 8186 19716 8188
rect 19740 8186 19796 8188
rect 19820 8186 19876 8188
rect 19580 8134 19606 8186
rect 19606 8134 19636 8186
rect 19660 8134 19670 8186
rect 19670 8134 19716 8186
rect 19740 8134 19786 8186
rect 19786 8134 19796 8186
rect 19820 8134 19850 8186
rect 19850 8134 19876 8186
rect 19580 8132 19636 8134
rect 19660 8132 19716 8134
rect 19740 8132 19796 8134
rect 19820 8132 19876 8134
rect 20994 7964 20996 7984
rect 20996 7964 21048 7984
rect 21048 7964 21050 7984
rect 20994 7928 21050 7964
rect 28170 7964 28172 7984
rect 28172 7964 28224 7984
rect 28224 7964 28226 7984
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 19580 7098 19636 7100
rect 19660 7098 19716 7100
rect 19740 7098 19796 7100
rect 19820 7098 19876 7100
rect 19580 7046 19606 7098
rect 19606 7046 19636 7098
rect 19660 7046 19670 7098
rect 19670 7046 19716 7098
rect 19740 7046 19786 7098
rect 19786 7046 19796 7098
rect 19820 7046 19850 7098
rect 19850 7046 19876 7098
rect 19580 7044 19636 7046
rect 19660 7044 19716 7046
rect 19740 7044 19796 7046
rect 19820 7044 19876 7046
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 1674 3052 1730 3088
rect 1674 3032 1676 3052
rect 1676 3032 1728 3052
rect 1728 3032 1730 3052
rect 1674 2508 1730 2544
rect 1674 2488 1676 2508
rect 1676 2488 1728 2508
rect 1728 2488 1730 2508
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 10138 3476 10140 3496
rect 10140 3476 10192 3496
rect 10192 3476 10194 3496
rect 10138 3440 10194 3476
rect 11886 3712 11942 3768
rect 11978 3032 12034 3088
rect 12438 4004 12494 4040
rect 12438 3984 12440 4004
rect 12440 3984 12492 4004
rect 12492 3984 12494 4004
rect 12622 3712 12678 3768
rect 12530 3068 12532 3088
rect 12532 3068 12584 3088
rect 12584 3068 12586 3088
rect 12530 3032 12586 3068
rect 15198 2896 15254 2952
rect 15658 3440 15714 3496
rect 17682 3168 17738 3224
rect 17498 2932 17500 2952
rect 17500 2932 17552 2952
rect 17552 2932 17554 2952
rect 17498 2896 17554 2932
rect 17682 2760 17738 2816
rect 18510 2760 18566 2816
rect 20534 6860 20590 6896
rect 20534 6840 20536 6860
rect 20536 6840 20588 6860
rect 20588 6840 20590 6860
rect 19580 6010 19636 6012
rect 19660 6010 19716 6012
rect 19740 6010 19796 6012
rect 19820 6010 19876 6012
rect 19580 5958 19606 6010
rect 19606 5958 19636 6010
rect 19660 5958 19670 6010
rect 19670 5958 19716 6010
rect 19740 5958 19786 6010
rect 19786 5958 19796 6010
rect 19820 5958 19850 6010
rect 19850 5958 19876 6010
rect 19580 5956 19636 5958
rect 19660 5956 19716 5958
rect 19740 5956 19796 5958
rect 19820 5956 19876 5958
rect 20994 6704 21050 6760
rect 20626 5652 20628 5672
rect 20628 5652 20680 5672
rect 20680 5652 20682 5672
rect 20626 5616 20682 5652
rect 22190 7540 22246 7576
rect 22190 7520 22192 7540
rect 22192 7520 22244 7540
rect 22244 7520 22246 7540
rect 21546 6704 21602 6760
rect 21638 5652 21640 5672
rect 21640 5652 21692 5672
rect 21692 5652 21694 5672
rect 21638 5616 21694 5652
rect 19580 4922 19636 4924
rect 19660 4922 19716 4924
rect 19740 4922 19796 4924
rect 19820 4922 19876 4924
rect 19580 4870 19606 4922
rect 19606 4870 19636 4922
rect 19660 4870 19670 4922
rect 19670 4870 19716 4922
rect 19740 4870 19786 4922
rect 19786 4870 19796 4922
rect 19820 4870 19850 4922
rect 19850 4870 19876 4922
rect 19580 4868 19636 4870
rect 19660 4868 19716 4870
rect 19740 4868 19796 4870
rect 19820 4868 19876 4870
rect 19580 3834 19636 3836
rect 19660 3834 19716 3836
rect 19740 3834 19796 3836
rect 19820 3834 19876 3836
rect 19580 3782 19606 3834
rect 19606 3782 19636 3834
rect 19660 3782 19670 3834
rect 19670 3782 19716 3834
rect 19740 3782 19786 3834
rect 19786 3782 19796 3834
rect 19820 3782 19850 3834
rect 19850 3782 19876 3834
rect 19580 3780 19636 3782
rect 19660 3780 19716 3782
rect 19740 3780 19796 3782
rect 19820 3780 19876 3782
rect 19062 3168 19118 3224
rect 19580 2746 19636 2748
rect 19660 2746 19716 2748
rect 19740 2746 19796 2748
rect 19820 2746 19876 2748
rect 19580 2694 19606 2746
rect 19606 2694 19636 2746
rect 19660 2694 19670 2746
rect 19670 2694 19716 2746
rect 19740 2694 19786 2746
rect 19786 2694 19796 2746
rect 19820 2694 19850 2746
rect 19850 2694 19876 2746
rect 19580 2692 19636 2694
rect 19660 2692 19716 2694
rect 19740 2692 19796 2694
rect 19820 2692 19876 2694
rect 20902 3576 20958 3632
rect 21270 3440 21326 3496
rect 21086 3168 21142 3224
rect 23018 6840 23074 6896
rect 28170 7928 28226 7964
rect 26514 7384 26570 7440
rect 21638 3984 21694 4040
rect 22098 3984 22154 4040
rect 22282 3476 22284 3496
rect 22284 3476 22336 3496
rect 22336 3476 22338 3496
rect 22282 3440 22338 3476
rect 22374 3068 22376 3088
rect 22376 3068 22428 3088
rect 22428 3068 22430 3088
rect 22374 3032 22430 3068
rect 28538 7656 28594 7712
rect 28446 7284 28448 7304
rect 28448 7284 28500 7304
rect 28500 7284 28502 7304
rect 28446 7248 28502 7284
rect 28906 7520 28962 7576
rect 28630 7112 28686 7168
rect 28538 6704 28594 6760
rect 28906 7112 28962 7168
rect 29642 7248 29698 7304
rect 30286 6740 30288 6760
rect 30288 6740 30340 6760
rect 30340 6740 30342 6760
rect 30286 6704 30342 6740
rect 30470 7248 30526 7304
rect 28170 3168 28226 3224
rect 28170 3068 28172 3088
rect 28172 3068 28224 3088
rect 28224 3068 28226 3088
rect 28170 3032 28226 3068
rect 28906 3576 28962 3632
rect 30562 3984 30618 4040
rect 31298 7284 31300 7304
rect 31300 7284 31352 7304
rect 31352 7284 31354 7304
rect 31298 7248 31354 7284
rect 34940 116442 34996 116444
rect 35020 116442 35076 116444
rect 35100 116442 35156 116444
rect 35180 116442 35236 116444
rect 34940 116390 34966 116442
rect 34966 116390 34996 116442
rect 35020 116390 35030 116442
rect 35030 116390 35076 116442
rect 35100 116390 35146 116442
rect 35146 116390 35156 116442
rect 35180 116390 35210 116442
rect 35210 116390 35236 116442
rect 34940 116388 34996 116390
rect 35020 116388 35076 116390
rect 35100 116388 35156 116390
rect 35180 116388 35236 116390
rect 34940 115354 34996 115356
rect 35020 115354 35076 115356
rect 35100 115354 35156 115356
rect 35180 115354 35236 115356
rect 34940 115302 34966 115354
rect 34966 115302 34996 115354
rect 35020 115302 35030 115354
rect 35030 115302 35076 115354
rect 35100 115302 35146 115354
rect 35146 115302 35156 115354
rect 35180 115302 35210 115354
rect 35210 115302 35236 115354
rect 34940 115300 34996 115302
rect 35020 115300 35076 115302
rect 35100 115300 35156 115302
rect 35180 115300 35236 115302
rect 34940 114266 34996 114268
rect 35020 114266 35076 114268
rect 35100 114266 35156 114268
rect 35180 114266 35236 114268
rect 34940 114214 34966 114266
rect 34966 114214 34996 114266
rect 35020 114214 35030 114266
rect 35030 114214 35076 114266
rect 35100 114214 35146 114266
rect 35146 114214 35156 114266
rect 35180 114214 35210 114266
rect 35210 114214 35236 114266
rect 34940 114212 34996 114214
rect 35020 114212 35076 114214
rect 35100 114212 35156 114214
rect 35180 114212 35236 114214
rect 34940 113178 34996 113180
rect 35020 113178 35076 113180
rect 35100 113178 35156 113180
rect 35180 113178 35236 113180
rect 34940 113126 34966 113178
rect 34966 113126 34996 113178
rect 35020 113126 35030 113178
rect 35030 113126 35076 113178
rect 35100 113126 35146 113178
rect 35146 113126 35156 113178
rect 35180 113126 35210 113178
rect 35210 113126 35236 113178
rect 34940 113124 34996 113126
rect 35020 113124 35076 113126
rect 35100 113124 35156 113126
rect 35180 113124 35236 113126
rect 34940 112090 34996 112092
rect 35020 112090 35076 112092
rect 35100 112090 35156 112092
rect 35180 112090 35236 112092
rect 34940 112038 34966 112090
rect 34966 112038 34996 112090
rect 35020 112038 35030 112090
rect 35030 112038 35076 112090
rect 35100 112038 35146 112090
rect 35146 112038 35156 112090
rect 35180 112038 35210 112090
rect 35210 112038 35236 112090
rect 34940 112036 34996 112038
rect 35020 112036 35076 112038
rect 35100 112036 35156 112038
rect 35180 112036 35236 112038
rect 34940 111002 34996 111004
rect 35020 111002 35076 111004
rect 35100 111002 35156 111004
rect 35180 111002 35236 111004
rect 34940 110950 34966 111002
rect 34966 110950 34996 111002
rect 35020 110950 35030 111002
rect 35030 110950 35076 111002
rect 35100 110950 35146 111002
rect 35146 110950 35156 111002
rect 35180 110950 35210 111002
rect 35210 110950 35236 111002
rect 34940 110948 34996 110950
rect 35020 110948 35076 110950
rect 35100 110948 35156 110950
rect 35180 110948 35236 110950
rect 34940 109914 34996 109916
rect 35020 109914 35076 109916
rect 35100 109914 35156 109916
rect 35180 109914 35236 109916
rect 34940 109862 34966 109914
rect 34966 109862 34996 109914
rect 35020 109862 35030 109914
rect 35030 109862 35076 109914
rect 35100 109862 35146 109914
rect 35146 109862 35156 109914
rect 35180 109862 35210 109914
rect 35210 109862 35236 109914
rect 34940 109860 34996 109862
rect 35020 109860 35076 109862
rect 35100 109860 35156 109862
rect 35180 109860 35236 109862
rect 34940 108826 34996 108828
rect 35020 108826 35076 108828
rect 35100 108826 35156 108828
rect 35180 108826 35236 108828
rect 34940 108774 34966 108826
rect 34966 108774 34996 108826
rect 35020 108774 35030 108826
rect 35030 108774 35076 108826
rect 35100 108774 35146 108826
rect 35146 108774 35156 108826
rect 35180 108774 35210 108826
rect 35210 108774 35236 108826
rect 34940 108772 34996 108774
rect 35020 108772 35076 108774
rect 35100 108772 35156 108774
rect 35180 108772 35236 108774
rect 34940 107738 34996 107740
rect 35020 107738 35076 107740
rect 35100 107738 35156 107740
rect 35180 107738 35236 107740
rect 34940 107686 34966 107738
rect 34966 107686 34996 107738
rect 35020 107686 35030 107738
rect 35030 107686 35076 107738
rect 35100 107686 35146 107738
rect 35146 107686 35156 107738
rect 35180 107686 35210 107738
rect 35210 107686 35236 107738
rect 34940 107684 34996 107686
rect 35020 107684 35076 107686
rect 35100 107684 35156 107686
rect 35180 107684 35236 107686
rect 34940 106650 34996 106652
rect 35020 106650 35076 106652
rect 35100 106650 35156 106652
rect 35180 106650 35236 106652
rect 34940 106598 34966 106650
rect 34966 106598 34996 106650
rect 35020 106598 35030 106650
rect 35030 106598 35076 106650
rect 35100 106598 35146 106650
rect 35146 106598 35156 106650
rect 35180 106598 35210 106650
rect 35210 106598 35236 106650
rect 34940 106596 34996 106598
rect 35020 106596 35076 106598
rect 35100 106596 35156 106598
rect 35180 106596 35236 106598
rect 34940 105562 34996 105564
rect 35020 105562 35076 105564
rect 35100 105562 35156 105564
rect 35180 105562 35236 105564
rect 34940 105510 34966 105562
rect 34966 105510 34996 105562
rect 35020 105510 35030 105562
rect 35030 105510 35076 105562
rect 35100 105510 35146 105562
rect 35146 105510 35156 105562
rect 35180 105510 35210 105562
rect 35210 105510 35236 105562
rect 34940 105508 34996 105510
rect 35020 105508 35076 105510
rect 35100 105508 35156 105510
rect 35180 105508 35236 105510
rect 34940 104474 34996 104476
rect 35020 104474 35076 104476
rect 35100 104474 35156 104476
rect 35180 104474 35236 104476
rect 34940 104422 34966 104474
rect 34966 104422 34996 104474
rect 35020 104422 35030 104474
rect 35030 104422 35076 104474
rect 35100 104422 35146 104474
rect 35146 104422 35156 104474
rect 35180 104422 35210 104474
rect 35210 104422 35236 104474
rect 34940 104420 34996 104422
rect 35020 104420 35076 104422
rect 35100 104420 35156 104422
rect 35180 104420 35236 104422
rect 34940 103386 34996 103388
rect 35020 103386 35076 103388
rect 35100 103386 35156 103388
rect 35180 103386 35236 103388
rect 34940 103334 34966 103386
rect 34966 103334 34996 103386
rect 35020 103334 35030 103386
rect 35030 103334 35076 103386
rect 35100 103334 35146 103386
rect 35146 103334 35156 103386
rect 35180 103334 35210 103386
rect 35210 103334 35236 103386
rect 34940 103332 34996 103334
rect 35020 103332 35076 103334
rect 35100 103332 35156 103334
rect 35180 103332 35236 103334
rect 34940 102298 34996 102300
rect 35020 102298 35076 102300
rect 35100 102298 35156 102300
rect 35180 102298 35236 102300
rect 34940 102246 34966 102298
rect 34966 102246 34996 102298
rect 35020 102246 35030 102298
rect 35030 102246 35076 102298
rect 35100 102246 35146 102298
rect 35146 102246 35156 102298
rect 35180 102246 35210 102298
rect 35210 102246 35236 102298
rect 34940 102244 34996 102246
rect 35020 102244 35076 102246
rect 35100 102244 35156 102246
rect 35180 102244 35236 102246
rect 34940 101210 34996 101212
rect 35020 101210 35076 101212
rect 35100 101210 35156 101212
rect 35180 101210 35236 101212
rect 34940 101158 34966 101210
rect 34966 101158 34996 101210
rect 35020 101158 35030 101210
rect 35030 101158 35076 101210
rect 35100 101158 35146 101210
rect 35146 101158 35156 101210
rect 35180 101158 35210 101210
rect 35210 101158 35236 101210
rect 34940 101156 34996 101158
rect 35020 101156 35076 101158
rect 35100 101156 35156 101158
rect 35180 101156 35236 101158
rect 34940 100122 34996 100124
rect 35020 100122 35076 100124
rect 35100 100122 35156 100124
rect 35180 100122 35236 100124
rect 34940 100070 34966 100122
rect 34966 100070 34996 100122
rect 35020 100070 35030 100122
rect 35030 100070 35076 100122
rect 35100 100070 35146 100122
rect 35146 100070 35156 100122
rect 35180 100070 35210 100122
rect 35210 100070 35236 100122
rect 34940 100068 34996 100070
rect 35020 100068 35076 100070
rect 35100 100068 35156 100070
rect 35180 100068 35236 100070
rect 34940 99034 34996 99036
rect 35020 99034 35076 99036
rect 35100 99034 35156 99036
rect 35180 99034 35236 99036
rect 34940 98982 34966 99034
rect 34966 98982 34996 99034
rect 35020 98982 35030 99034
rect 35030 98982 35076 99034
rect 35100 98982 35146 99034
rect 35146 98982 35156 99034
rect 35180 98982 35210 99034
rect 35210 98982 35236 99034
rect 34940 98980 34996 98982
rect 35020 98980 35076 98982
rect 35100 98980 35156 98982
rect 35180 98980 35236 98982
rect 34940 97946 34996 97948
rect 35020 97946 35076 97948
rect 35100 97946 35156 97948
rect 35180 97946 35236 97948
rect 34940 97894 34966 97946
rect 34966 97894 34996 97946
rect 35020 97894 35030 97946
rect 35030 97894 35076 97946
rect 35100 97894 35146 97946
rect 35146 97894 35156 97946
rect 35180 97894 35210 97946
rect 35210 97894 35236 97946
rect 34940 97892 34996 97894
rect 35020 97892 35076 97894
rect 35100 97892 35156 97894
rect 35180 97892 35236 97894
rect 34940 96858 34996 96860
rect 35020 96858 35076 96860
rect 35100 96858 35156 96860
rect 35180 96858 35236 96860
rect 34940 96806 34966 96858
rect 34966 96806 34996 96858
rect 35020 96806 35030 96858
rect 35030 96806 35076 96858
rect 35100 96806 35146 96858
rect 35146 96806 35156 96858
rect 35180 96806 35210 96858
rect 35210 96806 35236 96858
rect 34940 96804 34996 96806
rect 35020 96804 35076 96806
rect 35100 96804 35156 96806
rect 35180 96804 35236 96806
rect 34940 95770 34996 95772
rect 35020 95770 35076 95772
rect 35100 95770 35156 95772
rect 35180 95770 35236 95772
rect 34940 95718 34966 95770
rect 34966 95718 34996 95770
rect 35020 95718 35030 95770
rect 35030 95718 35076 95770
rect 35100 95718 35146 95770
rect 35146 95718 35156 95770
rect 35180 95718 35210 95770
rect 35210 95718 35236 95770
rect 34940 95716 34996 95718
rect 35020 95716 35076 95718
rect 35100 95716 35156 95718
rect 35180 95716 35236 95718
rect 34940 94682 34996 94684
rect 35020 94682 35076 94684
rect 35100 94682 35156 94684
rect 35180 94682 35236 94684
rect 34940 94630 34966 94682
rect 34966 94630 34996 94682
rect 35020 94630 35030 94682
rect 35030 94630 35076 94682
rect 35100 94630 35146 94682
rect 35146 94630 35156 94682
rect 35180 94630 35210 94682
rect 35210 94630 35236 94682
rect 34940 94628 34996 94630
rect 35020 94628 35076 94630
rect 35100 94628 35156 94630
rect 35180 94628 35236 94630
rect 34940 93594 34996 93596
rect 35020 93594 35076 93596
rect 35100 93594 35156 93596
rect 35180 93594 35236 93596
rect 34940 93542 34966 93594
rect 34966 93542 34996 93594
rect 35020 93542 35030 93594
rect 35030 93542 35076 93594
rect 35100 93542 35146 93594
rect 35146 93542 35156 93594
rect 35180 93542 35210 93594
rect 35210 93542 35236 93594
rect 34940 93540 34996 93542
rect 35020 93540 35076 93542
rect 35100 93540 35156 93542
rect 35180 93540 35236 93542
rect 34940 92506 34996 92508
rect 35020 92506 35076 92508
rect 35100 92506 35156 92508
rect 35180 92506 35236 92508
rect 34940 92454 34966 92506
rect 34966 92454 34996 92506
rect 35020 92454 35030 92506
rect 35030 92454 35076 92506
rect 35100 92454 35146 92506
rect 35146 92454 35156 92506
rect 35180 92454 35210 92506
rect 35210 92454 35236 92506
rect 34940 92452 34996 92454
rect 35020 92452 35076 92454
rect 35100 92452 35156 92454
rect 35180 92452 35236 92454
rect 34940 91418 34996 91420
rect 35020 91418 35076 91420
rect 35100 91418 35156 91420
rect 35180 91418 35236 91420
rect 34940 91366 34966 91418
rect 34966 91366 34996 91418
rect 35020 91366 35030 91418
rect 35030 91366 35076 91418
rect 35100 91366 35146 91418
rect 35146 91366 35156 91418
rect 35180 91366 35210 91418
rect 35210 91366 35236 91418
rect 34940 91364 34996 91366
rect 35020 91364 35076 91366
rect 35100 91364 35156 91366
rect 35180 91364 35236 91366
rect 34940 90330 34996 90332
rect 35020 90330 35076 90332
rect 35100 90330 35156 90332
rect 35180 90330 35236 90332
rect 34940 90278 34966 90330
rect 34966 90278 34996 90330
rect 35020 90278 35030 90330
rect 35030 90278 35076 90330
rect 35100 90278 35146 90330
rect 35146 90278 35156 90330
rect 35180 90278 35210 90330
rect 35210 90278 35236 90330
rect 34940 90276 34996 90278
rect 35020 90276 35076 90278
rect 35100 90276 35156 90278
rect 35180 90276 35236 90278
rect 34940 89242 34996 89244
rect 35020 89242 35076 89244
rect 35100 89242 35156 89244
rect 35180 89242 35236 89244
rect 34940 89190 34966 89242
rect 34966 89190 34996 89242
rect 35020 89190 35030 89242
rect 35030 89190 35076 89242
rect 35100 89190 35146 89242
rect 35146 89190 35156 89242
rect 35180 89190 35210 89242
rect 35210 89190 35236 89242
rect 34940 89188 34996 89190
rect 35020 89188 35076 89190
rect 35100 89188 35156 89190
rect 35180 89188 35236 89190
rect 34940 88154 34996 88156
rect 35020 88154 35076 88156
rect 35100 88154 35156 88156
rect 35180 88154 35236 88156
rect 34940 88102 34966 88154
rect 34966 88102 34996 88154
rect 35020 88102 35030 88154
rect 35030 88102 35076 88154
rect 35100 88102 35146 88154
rect 35146 88102 35156 88154
rect 35180 88102 35210 88154
rect 35210 88102 35236 88154
rect 34940 88100 34996 88102
rect 35020 88100 35076 88102
rect 35100 88100 35156 88102
rect 35180 88100 35236 88102
rect 34940 87066 34996 87068
rect 35020 87066 35076 87068
rect 35100 87066 35156 87068
rect 35180 87066 35236 87068
rect 34940 87014 34966 87066
rect 34966 87014 34996 87066
rect 35020 87014 35030 87066
rect 35030 87014 35076 87066
rect 35100 87014 35146 87066
rect 35146 87014 35156 87066
rect 35180 87014 35210 87066
rect 35210 87014 35236 87066
rect 34940 87012 34996 87014
rect 35020 87012 35076 87014
rect 35100 87012 35156 87014
rect 35180 87012 35236 87014
rect 34940 85978 34996 85980
rect 35020 85978 35076 85980
rect 35100 85978 35156 85980
rect 35180 85978 35236 85980
rect 34940 85926 34966 85978
rect 34966 85926 34996 85978
rect 35020 85926 35030 85978
rect 35030 85926 35076 85978
rect 35100 85926 35146 85978
rect 35146 85926 35156 85978
rect 35180 85926 35210 85978
rect 35210 85926 35236 85978
rect 34940 85924 34996 85926
rect 35020 85924 35076 85926
rect 35100 85924 35156 85926
rect 35180 85924 35236 85926
rect 34940 84890 34996 84892
rect 35020 84890 35076 84892
rect 35100 84890 35156 84892
rect 35180 84890 35236 84892
rect 34940 84838 34966 84890
rect 34966 84838 34996 84890
rect 35020 84838 35030 84890
rect 35030 84838 35076 84890
rect 35100 84838 35146 84890
rect 35146 84838 35156 84890
rect 35180 84838 35210 84890
rect 35210 84838 35236 84890
rect 34940 84836 34996 84838
rect 35020 84836 35076 84838
rect 35100 84836 35156 84838
rect 35180 84836 35236 84838
rect 34940 83802 34996 83804
rect 35020 83802 35076 83804
rect 35100 83802 35156 83804
rect 35180 83802 35236 83804
rect 34940 83750 34966 83802
rect 34966 83750 34996 83802
rect 35020 83750 35030 83802
rect 35030 83750 35076 83802
rect 35100 83750 35146 83802
rect 35146 83750 35156 83802
rect 35180 83750 35210 83802
rect 35210 83750 35236 83802
rect 34940 83748 34996 83750
rect 35020 83748 35076 83750
rect 35100 83748 35156 83750
rect 35180 83748 35236 83750
rect 34940 82714 34996 82716
rect 35020 82714 35076 82716
rect 35100 82714 35156 82716
rect 35180 82714 35236 82716
rect 34940 82662 34966 82714
rect 34966 82662 34996 82714
rect 35020 82662 35030 82714
rect 35030 82662 35076 82714
rect 35100 82662 35146 82714
rect 35146 82662 35156 82714
rect 35180 82662 35210 82714
rect 35210 82662 35236 82714
rect 34940 82660 34996 82662
rect 35020 82660 35076 82662
rect 35100 82660 35156 82662
rect 35180 82660 35236 82662
rect 34940 81626 34996 81628
rect 35020 81626 35076 81628
rect 35100 81626 35156 81628
rect 35180 81626 35236 81628
rect 34940 81574 34966 81626
rect 34966 81574 34996 81626
rect 35020 81574 35030 81626
rect 35030 81574 35076 81626
rect 35100 81574 35146 81626
rect 35146 81574 35156 81626
rect 35180 81574 35210 81626
rect 35210 81574 35236 81626
rect 34940 81572 34996 81574
rect 35020 81572 35076 81574
rect 35100 81572 35156 81574
rect 35180 81572 35236 81574
rect 34940 80538 34996 80540
rect 35020 80538 35076 80540
rect 35100 80538 35156 80540
rect 35180 80538 35236 80540
rect 34940 80486 34966 80538
rect 34966 80486 34996 80538
rect 35020 80486 35030 80538
rect 35030 80486 35076 80538
rect 35100 80486 35146 80538
rect 35146 80486 35156 80538
rect 35180 80486 35210 80538
rect 35210 80486 35236 80538
rect 34940 80484 34996 80486
rect 35020 80484 35076 80486
rect 35100 80484 35156 80486
rect 35180 80484 35236 80486
rect 34940 79450 34996 79452
rect 35020 79450 35076 79452
rect 35100 79450 35156 79452
rect 35180 79450 35236 79452
rect 34940 79398 34966 79450
rect 34966 79398 34996 79450
rect 35020 79398 35030 79450
rect 35030 79398 35076 79450
rect 35100 79398 35146 79450
rect 35146 79398 35156 79450
rect 35180 79398 35210 79450
rect 35210 79398 35236 79450
rect 34940 79396 34996 79398
rect 35020 79396 35076 79398
rect 35100 79396 35156 79398
rect 35180 79396 35236 79398
rect 34940 78362 34996 78364
rect 35020 78362 35076 78364
rect 35100 78362 35156 78364
rect 35180 78362 35236 78364
rect 34940 78310 34966 78362
rect 34966 78310 34996 78362
rect 35020 78310 35030 78362
rect 35030 78310 35076 78362
rect 35100 78310 35146 78362
rect 35146 78310 35156 78362
rect 35180 78310 35210 78362
rect 35210 78310 35236 78362
rect 34940 78308 34996 78310
rect 35020 78308 35076 78310
rect 35100 78308 35156 78310
rect 35180 78308 35236 78310
rect 34940 77274 34996 77276
rect 35020 77274 35076 77276
rect 35100 77274 35156 77276
rect 35180 77274 35236 77276
rect 34940 77222 34966 77274
rect 34966 77222 34996 77274
rect 35020 77222 35030 77274
rect 35030 77222 35076 77274
rect 35100 77222 35146 77274
rect 35146 77222 35156 77274
rect 35180 77222 35210 77274
rect 35210 77222 35236 77274
rect 34940 77220 34996 77222
rect 35020 77220 35076 77222
rect 35100 77220 35156 77222
rect 35180 77220 35236 77222
rect 34940 76186 34996 76188
rect 35020 76186 35076 76188
rect 35100 76186 35156 76188
rect 35180 76186 35236 76188
rect 34940 76134 34966 76186
rect 34966 76134 34996 76186
rect 35020 76134 35030 76186
rect 35030 76134 35076 76186
rect 35100 76134 35146 76186
rect 35146 76134 35156 76186
rect 35180 76134 35210 76186
rect 35210 76134 35236 76186
rect 34940 76132 34996 76134
rect 35020 76132 35076 76134
rect 35100 76132 35156 76134
rect 35180 76132 35236 76134
rect 34940 75098 34996 75100
rect 35020 75098 35076 75100
rect 35100 75098 35156 75100
rect 35180 75098 35236 75100
rect 34940 75046 34966 75098
rect 34966 75046 34996 75098
rect 35020 75046 35030 75098
rect 35030 75046 35076 75098
rect 35100 75046 35146 75098
rect 35146 75046 35156 75098
rect 35180 75046 35210 75098
rect 35210 75046 35236 75098
rect 34940 75044 34996 75046
rect 35020 75044 35076 75046
rect 35100 75044 35156 75046
rect 35180 75044 35236 75046
rect 34940 74010 34996 74012
rect 35020 74010 35076 74012
rect 35100 74010 35156 74012
rect 35180 74010 35236 74012
rect 34940 73958 34966 74010
rect 34966 73958 34996 74010
rect 35020 73958 35030 74010
rect 35030 73958 35076 74010
rect 35100 73958 35146 74010
rect 35146 73958 35156 74010
rect 35180 73958 35210 74010
rect 35210 73958 35236 74010
rect 34940 73956 34996 73958
rect 35020 73956 35076 73958
rect 35100 73956 35156 73958
rect 35180 73956 35236 73958
rect 34940 72922 34996 72924
rect 35020 72922 35076 72924
rect 35100 72922 35156 72924
rect 35180 72922 35236 72924
rect 34940 72870 34966 72922
rect 34966 72870 34996 72922
rect 35020 72870 35030 72922
rect 35030 72870 35076 72922
rect 35100 72870 35146 72922
rect 35146 72870 35156 72922
rect 35180 72870 35210 72922
rect 35210 72870 35236 72922
rect 34940 72868 34996 72870
rect 35020 72868 35076 72870
rect 35100 72868 35156 72870
rect 35180 72868 35236 72870
rect 34940 71834 34996 71836
rect 35020 71834 35076 71836
rect 35100 71834 35156 71836
rect 35180 71834 35236 71836
rect 34940 71782 34966 71834
rect 34966 71782 34996 71834
rect 35020 71782 35030 71834
rect 35030 71782 35076 71834
rect 35100 71782 35146 71834
rect 35146 71782 35156 71834
rect 35180 71782 35210 71834
rect 35210 71782 35236 71834
rect 34940 71780 34996 71782
rect 35020 71780 35076 71782
rect 35100 71780 35156 71782
rect 35180 71780 35236 71782
rect 34940 70746 34996 70748
rect 35020 70746 35076 70748
rect 35100 70746 35156 70748
rect 35180 70746 35236 70748
rect 34940 70694 34966 70746
rect 34966 70694 34996 70746
rect 35020 70694 35030 70746
rect 35030 70694 35076 70746
rect 35100 70694 35146 70746
rect 35146 70694 35156 70746
rect 35180 70694 35210 70746
rect 35210 70694 35236 70746
rect 34940 70692 34996 70694
rect 35020 70692 35076 70694
rect 35100 70692 35156 70694
rect 35180 70692 35236 70694
rect 34940 69658 34996 69660
rect 35020 69658 35076 69660
rect 35100 69658 35156 69660
rect 35180 69658 35236 69660
rect 34940 69606 34966 69658
rect 34966 69606 34996 69658
rect 35020 69606 35030 69658
rect 35030 69606 35076 69658
rect 35100 69606 35146 69658
rect 35146 69606 35156 69658
rect 35180 69606 35210 69658
rect 35210 69606 35236 69658
rect 34940 69604 34996 69606
rect 35020 69604 35076 69606
rect 35100 69604 35156 69606
rect 35180 69604 35236 69606
rect 34940 68570 34996 68572
rect 35020 68570 35076 68572
rect 35100 68570 35156 68572
rect 35180 68570 35236 68572
rect 34940 68518 34966 68570
rect 34966 68518 34996 68570
rect 35020 68518 35030 68570
rect 35030 68518 35076 68570
rect 35100 68518 35146 68570
rect 35146 68518 35156 68570
rect 35180 68518 35210 68570
rect 35210 68518 35236 68570
rect 34940 68516 34996 68518
rect 35020 68516 35076 68518
rect 35100 68516 35156 68518
rect 35180 68516 35236 68518
rect 34940 67482 34996 67484
rect 35020 67482 35076 67484
rect 35100 67482 35156 67484
rect 35180 67482 35236 67484
rect 34940 67430 34966 67482
rect 34966 67430 34996 67482
rect 35020 67430 35030 67482
rect 35030 67430 35076 67482
rect 35100 67430 35146 67482
rect 35146 67430 35156 67482
rect 35180 67430 35210 67482
rect 35210 67430 35236 67482
rect 34940 67428 34996 67430
rect 35020 67428 35076 67430
rect 35100 67428 35156 67430
rect 35180 67428 35236 67430
rect 34940 66394 34996 66396
rect 35020 66394 35076 66396
rect 35100 66394 35156 66396
rect 35180 66394 35236 66396
rect 34940 66342 34966 66394
rect 34966 66342 34996 66394
rect 35020 66342 35030 66394
rect 35030 66342 35076 66394
rect 35100 66342 35146 66394
rect 35146 66342 35156 66394
rect 35180 66342 35210 66394
rect 35210 66342 35236 66394
rect 34940 66340 34996 66342
rect 35020 66340 35076 66342
rect 35100 66340 35156 66342
rect 35180 66340 35236 66342
rect 34940 65306 34996 65308
rect 35020 65306 35076 65308
rect 35100 65306 35156 65308
rect 35180 65306 35236 65308
rect 34940 65254 34966 65306
rect 34966 65254 34996 65306
rect 35020 65254 35030 65306
rect 35030 65254 35076 65306
rect 35100 65254 35146 65306
rect 35146 65254 35156 65306
rect 35180 65254 35210 65306
rect 35210 65254 35236 65306
rect 34940 65252 34996 65254
rect 35020 65252 35076 65254
rect 35100 65252 35156 65254
rect 35180 65252 35236 65254
rect 34940 64218 34996 64220
rect 35020 64218 35076 64220
rect 35100 64218 35156 64220
rect 35180 64218 35236 64220
rect 34940 64166 34966 64218
rect 34966 64166 34996 64218
rect 35020 64166 35030 64218
rect 35030 64166 35076 64218
rect 35100 64166 35146 64218
rect 35146 64166 35156 64218
rect 35180 64166 35210 64218
rect 35210 64166 35236 64218
rect 34940 64164 34996 64166
rect 35020 64164 35076 64166
rect 35100 64164 35156 64166
rect 35180 64164 35236 64166
rect 34940 63130 34996 63132
rect 35020 63130 35076 63132
rect 35100 63130 35156 63132
rect 35180 63130 35236 63132
rect 34940 63078 34966 63130
rect 34966 63078 34996 63130
rect 35020 63078 35030 63130
rect 35030 63078 35076 63130
rect 35100 63078 35146 63130
rect 35146 63078 35156 63130
rect 35180 63078 35210 63130
rect 35210 63078 35236 63130
rect 34940 63076 34996 63078
rect 35020 63076 35076 63078
rect 35100 63076 35156 63078
rect 35180 63076 35236 63078
rect 34940 62042 34996 62044
rect 35020 62042 35076 62044
rect 35100 62042 35156 62044
rect 35180 62042 35236 62044
rect 34940 61990 34966 62042
rect 34966 61990 34996 62042
rect 35020 61990 35030 62042
rect 35030 61990 35076 62042
rect 35100 61990 35146 62042
rect 35146 61990 35156 62042
rect 35180 61990 35210 62042
rect 35210 61990 35236 62042
rect 34940 61988 34996 61990
rect 35020 61988 35076 61990
rect 35100 61988 35156 61990
rect 35180 61988 35236 61990
rect 34940 60954 34996 60956
rect 35020 60954 35076 60956
rect 35100 60954 35156 60956
rect 35180 60954 35236 60956
rect 34940 60902 34966 60954
rect 34966 60902 34996 60954
rect 35020 60902 35030 60954
rect 35030 60902 35076 60954
rect 35100 60902 35146 60954
rect 35146 60902 35156 60954
rect 35180 60902 35210 60954
rect 35210 60902 35236 60954
rect 34940 60900 34996 60902
rect 35020 60900 35076 60902
rect 35100 60900 35156 60902
rect 35180 60900 35236 60902
rect 34940 59866 34996 59868
rect 35020 59866 35076 59868
rect 35100 59866 35156 59868
rect 35180 59866 35236 59868
rect 34940 59814 34966 59866
rect 34966 59814 34996 59866
rect 35020 59814 35030 59866
rect 35030 59814 35076 59866
rect 35100 59814 35146 59866
rect 35146 59814 35156 59866
rect 35180 59814 35210 59866
rect 35210 59814 35236 59866
rect 34940 59812 34996 59814
rect 35020 59812 35076 59814
rect 35100 59812 35156 59814
rect 35180 59812 35236 59814
rect 34940 58778 34996 58780
rect 35020 58778 35076 58780
rect 35100 58778 35156 58780
rect 35180 58778 35236 58780
rect 34940 58726 34966 58778
rect 34966 58726 34996 58778
rect 35020 58726 35030 58778
rect 35030 58726 35076 58778
rect 35100 58726 35146 58778
rect 35146 58726 35156 58778
rect 35180 58726 35210 58778
rect 35210 58726 35236 58778
rect 34940 58724 34996 58726
rect 35020 58724 35076 58726
rect 35100 58724 35156 58726
rect 35180 58724 35236 58726
rect 34940 57690 34996 57692
rect 35020 57690 35076 57692
rect 35100 57690 35156 57692
rect 35180 57690 35236 57692
rect 34940 57638 34966 57690
rect 34966 57638 34996 57690
rect 35020 57638 35030 57690
rect 35030 57638 35076 57690
rect 35100 57638 35146 57690
rect 35146 57638 35156 57690
rect 35180 57638 35210 57690
rect 35210 57638 35236 57690
rect 34940 57636 34996 57638
rect 35020 57636 35076 57638
rect 35100 57636 35156 57638
rect 35180 57636 35236 57638
rect 34940 56602 34996 56604
rect 35020 56602 35076 56604
rect 35100 56602 35156 56604
rect 35180 56602 35236 56604
rect 34940 56550 34966 56602
rect 34966 56550 34996 56602
rect 35020 56550 35030 56602
rect 35030 56550 35076 56602
rect 35100 56550 35146 56602
rect 35146 56550 35156 56602
rect 35180 56550 35210 56602
rect 35210 56550 35236 56602
rect 34940 56548 34996 56550
rect 35020 56548 35076 56550
rect 35100 56548 35156 56550
rect 35180 56548 35236 56550
rect 34940 55514 34996 55516
rect 35020 55514 35076 55516
rect 35100 55514 35156 55516
rect 35180 55514 35236 55516
rect 34940 55462 34966 55514
rect 34966 55462 34996 55514
rect 35020 55462 35030 55514
rect 35030 55462 35076 55514
rect 35100 55462 35146 55514
rect 35146 55462 35156 55514
rect 35180 55462 35210 55514
rect 35210 55462 35236 55514
rect 34940 55460 34996 55462
rect 35020 55460 35076 55462
rect 35100 55460 35156 55462
rect 35180 55460 35236 55462
rect 34940 54426 34996 54428
rect 35020 54426 35076 54428
rect 35100 54426 35156 54428
rect 35180 54426 35236 54428
rect 34940 54374 34966 54426
rect 34966 54374 34996 54426
rect 35020 54374 35030 54426
rect 35030 54374 35076 54426
rect 35100 54374 35146 54426
rect 35146 54374 35156 54426
rect 35180 54374 35210 54426
rect 35210 54374 35236 54426
rect 34940 54372 34996 54374
rect 35020 54372 35076 54374
rect 35100 54372 35156 54374
rect 35180 54372 35236 54374
rect 34940 53338 34996 53340
rect 35020 53338 35076 53340
rect 35100 53338 35156 53340
rect 35180 53338 35236 53340
rect 34940 53286 34966 53338
rect 34966 53286 34996 53338
rect 35020 53286 35030 53338
rect 35030 53286 35076 53338
rect 35100 53286 35146 53338
rect 35146 53286 35156 53338
rect 35180 53286 35210 53338
rect 35210 53286 35236 53338
rect 34940 53284 34996 53286
rect 35020 53284 35076 53286
rect 35100 53284 35156 53286
rect 35180 53284 35236 53286
rect 34940 52250 34996 52252
rect 35020 52250 35076 52252
rect 35100 52250 35156 52252
rect 35180 52250 35236 52252
rect 34940 52198 34966 52250
rect 34966 52198 34996 52250
rect 35020 52198 35030 52250
rect 35030 52198 35076 52250
rect 35100 52198 35146 52250
rect 35146 52198 35156 52250
rect 35180 52198 35210 52250
rect 35210 52198 35236 52250
rect 34940 52196 34996 52198
rect 35020 52196 35076 52198
rect 35100 52196 35156 52198
rect 35180 52196 35236 52198
rect 34940 51162 34996 51164
rect 35020 51162 35076 51164
rect 35100 51162 35156 51164
rect 35180 51162 35236 51164
rect 34940 51110 34966 51162
rect 34966 51110 34996 51162
rect 35020 51110 35030 51162
rect 35030 51110 35076 51162
rect 35100 51110 35146 51162
rect 35146 51110 35156 51162
rect 35180 51110 35210 51162
rect 35210 51110 35236 51162
rect 34940 51108 34996 51110
rect 35020 51108 35076 51110
rect 35100 51108 35156 51110
rect 35180 51108 35236 51110
rect 34940 50074 34996 50076
rect 35020 50074 35076 50076
rect 35100 50074 35156 50076
rect 35180 50074 35236 50076
rect 34940 50022 34966 50074
rect 34966 50022 34996 50074
rect 35020 50022 35030 50074
rect 35030 50022 35076 50074
rect 35100 50022 35146 50074
rect 35146 50022 35156 50074
rect 35180 50022 35210 50074
rect 35210 50022 35236 50074
rect 34940 50020 34996 50022
rect 35020 50020 35076 50022
rect 35100 50020 35156 50022
rect 35180 50020 35236 50022
rect 34940 48986 34996 48988
rect 35020 48986 35076 48988
rect 35100 48986 35156 48988
rect 35180 48986 35236 48988
rect 34940 48934 34966 48986
rect 34966 48934 34996 48986
rect 35020 48934 35030 48986
rect 35030 48934 35076 48986
rect 35100 48934 35146 48986
rect 35146 48934 35156 48986
rect 35180 48934 35210 48986
rect 35210 48934 35236 48986
rect 34940 48932 34996 48934
rect 35020 48932 35076 48934
rect 35100 48932 35156 48934
rect 35180 48932 35236 48934
rect 34940 47898 34996 47900
rect 35020 47898 35076 47900
rect 35100 47898 35156 47900
rect 35180 47898 35236 47900
rect 34940 47846 34966 47898
rect 34966 47846 34996 47898
rect 35020 47846 35030 47898
rect 35030 47846 35076 47898
rect 35100 47846 35146 47898
rect 35146 47846 35156 47898
rect 35180 47846 35210 47898
rect 35210 47846 35236 47898
rect 34940 47844 34996 47846
rect 35020 47844 35076 47846
rect 35100 47844 35156 47846
rect 35180 47844 35236 47846
rect 34940 46810 34996 46812
rect 35020 46810 35076 46812
rect 35100 46810 35156 46812
rect 35180 46810 35236 46812
rect 34940 46758 34966 46810
rect 34966 46758 34996 46810
rect 35020 46758 35030 46810
rect 35030 46758 35076 46810
rect 35100 46758 35146 46810
rect 35146 46758 35156 46810
rect 35180 46758 35210 46810
rect 35210 46758 35236 46810
rect 34940 46756 34996 46758
rect 35020 46756 35076 46758
rect 35100 46756 35156 46758
rect 35180 46756 35236 46758
rect 34940 45722 34996 45724
rect 35020 45722 35076 45724
rect 35100 45722 35156 45724
rect 35180 45722 35236 45724
rect 34940 45670 34966 45722
rect 34966 45670 34996 45722
rect 35020 45670 35030 45722
rect 35030 45670 35076 45722
rect 35100 45670 35146 45722
rect 35146 45670 35156 45722
rect 35180 45670 35210 45722
rect 35210 45670 35236 45722
rect 34940 45668 34996 45670
rect 35020 45668 35076 45670
rect 35100 45668 35156 45670
rect 35180 45668 35236 45670
rect 34940 44634 34996 44636
rect 35020 44634 35076 44636
rect 35100 44634 35156 44636
rect 35180 44634 35236 44636
rect 34940 44582 34966 44634
rect 34966 44582 34996 44634
rect 35020 44582 35030 44634
rect 35030 44582 35076 44634
rect 35100 44582 35146 44634
rect 35146 44582 35156 44634
rect 35180 44582 35210 44634
rect 35210 44582 35236 44634
rect 34940 44580 34996 44582
rect 35020 44580 35076 44582
rect 35100 44580 35156 44582
rect 35180 44580 35236 44582
rect 34940 43546 34996 43548
rect 35020 43546 35076 43548
rect 35100 43546 35156 43548
rect 35180 43546 35236 43548
rect 34940 43494 34966 43546
rect 34966 43494 34996 43546
rect 35020 43494 35030 43546
rect 35030 43494 35076 43546
rect 35100 43494 35146 43546
rect 35146 43494 35156 43546
rect 35180 43494 35210 43546
rect 35210 43494 35236 43546
rect 34940 43492 34996 43494
rect 35020 43492 35076 43494
rect 35100 43492 35156 43494
rect 35180 43492 35236 43494
rect 34940 42458 34996 42460
rect 35020 42458 35076 42460
rect 35100 42458 35156 42460
rect 35180 42458 35236 42460
rect 34940 42406 34966 42458
rect 34966 42406 34996 42458
rect 35020 42406 35030 42458
rect 35030 42406 35076 42458
rect 35100 42406 35146 42458
rect 35146 42406 35156 42458
rect 35180 42406 35210 42458
rect 35210 42406 35236 42458
rect 34940 42404 34996 42406
rect 35020 42404 35076 42406
rect 35100 42404 35156 42406
rect 35180 42404 35236 42406
rect 34940 41370 34996 41372
rect 35020 41370 35076 41372
rect 35100 41370 35156 41372
rect 35180 41370 35236 41372
rect 34940 41318 34966 41370
rect 34966 41318 34996 41370
rect 35020 41318 35030 41370
rect 35030 41318 35076 41370
rect 35100 41318 35146 41370
rect 35146 41318 35156 41370
rect 35180 41318 35210 41370
rect 35210 41318 35236 41370
rect 34940 41316 34996 41318
rect 35020 41316 35076 41318
rect 35100 41316 35156 41318
rect 35180 41316 35236 41318
rect 34940 40282 34996 40284
rect 35020 40282 35076 40284
rect 35100 40282 35156 40284
rect 35180 40282 35236 40284
rect 34940 40230 34966 40282
rect 34966 40230 34996 40282
rect 35020 40230 35030 40282
rect 35030 40230 35076 40282
rect 35100 40230 35146 40282
rect 35146 40230 35156 40282
rect 35180 40230 35210 40282
rect 35210 40230 35236 40282
rect 34940 40228 34996 40230
rect 35020 40228 35076 40230
rect 35100 40228 35156 40230
rect 35180 40228 35236 40230
rect 34940 39194 34996 39196
rect 35020 39194 35076 39196
rect 35100 39194 35156 39196
rect 35180 39194 35236 39196
rect 34940 39142 34966 39194
rect 34966 39142 34996 39194
rect 35020 39142 35030 39194
rect 35030 39142 35076 39194
rect 35100 39142 35146 39194
rect 35146 39142 35156 39194
rect 35180 39142 35210 39194
rect 35210 39142 35236 39194
rect 34940 39140 34996 39142
rect 35020 39140 35076 39142
rect 35100 39140 35156 39142
rect 35180 39140 35236 39142
rect 34940 38106 34996 38108
rect 35020 38106 35076 38108
rect 35100 38106 35156 38108
rect 35180 38106 35236 38108
rect 34940 38054 34966 38106
rect 34966 38054 34996 38106
rect 35020 38054 35030 38106
rect 35030 38054 35076 38106
rect 35100 38054 35146 38106
rect 35146 38054 35156 38106
rect 35180 38054 35210 38106
rect 35210 38054 35236 38106
rect 34940 38052 34996 38054
rect 35020 38052 35076 38054
rect 35100 38052 35156 38054
rect 35180 38052 35236 38054
rect 34940 37018 34996 37020
rect 35020 37018 35076 37020
rect 35100 37018 35156 37020
rect 35180 37018 35236 37020
rect 34940 36966 34966 37018
rect 34966 36966 34996 37018
rect 35020 36966 35030 37018
rect 35030 36966 35076 37018
rect 35100 36966 35146 37018
rect 35146 36966 35156 37018
rect 35180 36966 35210 37018
rect 35210 36966 35236 37018
rect 34940 36964 34996 36966
rect 35020 36964 35076 36966
rect 35100 36964 35156 36966
rect 35180 36964 35236 36966
rect 34940 35930 34996 35932
rect 35020 35930 35076 35932
rect 35100 35930 35156 35932
rect 35180 35930 35236 35932
rect 34940 35878 34966 35930
rect 34966 35878 34996 35930
rect 35020 35878 35030 35930
rect 35030 35878 35076 35930
rect 35100 35878 35146 35930
rect 35146 35878 35156 35930
rect 35180 35878 35210 35930
rect 35210 35878 35236 35930
rect 34940 35876 34996 35878
rect 35020 35876 35076 35878
rect 35100 35876 35156 35878
rect 35180 35876 35236 35878
rect 34940 34842 34996 34844
rect 35020 34842 35076 34844
rect 35100 34842 35156 34844
rect 35180 34842 35236 34844
rect 34940 34790 34966 34842
rect 34966 34790 34996 34842
rect 35020 34790 35030 34842
rect 35030 34790 35076 34842
rect 35100 34790 35146 34842
rect 35146 34790 35156 34842
rect 35180 34790 35210 34842
rect 35210 34790 35236 34842
rect 34940 34788 34996 34790
rect 35020 34788 35076 34790
rect 35100 34788 35156 34790
rect 35180 34788 35236 34790
rect 34940 33754 34996 33756
rect 35020 33754 35076 33756
rect 35100 33754 35156 33756
rect 35180 33754 35236 33756
rect 34940 33702 34966 33754
rect 34966 33702 34996 33754
rect 35020 33702 35030 33754
rect 35030 33702 35076 33754
rect 35100 33702 35146 33754
rect 35146 33702 35156 33754
rect 35180 33702 35210 33754
rect 35210 33702 35236 33754
rect 34940 33700 34996 33702
rect 35020 33700 35076 33702
rect 35100 33700 35156 33702
rect 35180 33700 35236 33702
rect 34940 32666 34996 32668
rect 35020 32666 35076 32668
rect 35100 32666 35156 32668
rect 35180 32666 35236 32668
rect 34940 32614 34966 32666
rect 34966 32614 34996 32666
rect 35020 32614 35030 32666
rect 35030 32614 35076 32666
rect 35100 32614 35146 32666
rect 35146 32614 35156 32666
rect 35180 32614 35210 32666
rect 35210 32614 35236 32666
rect 34940 32612 34996 32614
rect 35020 32612 35076 32614
rect 35100 32612 35156 32614
rect 35180 32612 35236 32614
rect 34940 31578 34996 31580
rect 35020 31578 35076 31580
rect 35100 31578 35156 31580
rect 35180 31578 35236 31580
rect 34940 31526 34966 31578
rect 34966 31526 34996 31578
rect 35020 31526 35030 31578
rect 35030 31526 35076 31578
rect 35100 31526 35146 31578
rect 35146 31526 35156 31578
rect 35180 31526 35210 31578
rect 35210 31526 35236 31578
rect 34940 31524 34996 31526
rect 35020 31524 35076 31526
rect 35100 31524 35156 31526
rect 35180 31524 35236 31526
rect 34940 30490 34996 30492
rect 35020 30490 35076 30492
rect 35100 30490 35156 30492
rect 35180 30490 35236 30492
rect 34940 30438 34966 30490
rect 34966 30438 34996 30490
rect 35020 30438 35030 30490
rect 35030 30438 35076 30490
rect 35100 30438 35146 30490
rect 35146 30438 35156 30490
rect 35180 30438 35210 30490
rect 35210 30438 35236 30490
rect 34940 30436 34996 30438
rect 35020 30436 35076 30438
rect 35100 30436 35156 30438
rect 35180 30436 35236 30438
rect 34940 29402 34996 29404
rect 35020 29402 35076 29404
rect 35100 29402 35156 29404
rect 35180 29402 35236 29404
rect 34940 29350 34966 29402
rect 34966 29350 34996 29402
rect 35020 29350 35030 29402
rect 35030 29350 35076 29402
rect 35100 29350 35146 29402
rect 35146 29350 35156 29402
rect 35180 29350 35210 29402
rect 35210 29350 35236 29402
rect 34940 29348 34996 29350
rect 35020 29348 35076 29350
rect 35100 29348 35156 29350
rect 35180 29348 35236 29350
rect 34940 28314 34996 28316
rect 35020 28314 35076 28316
rect 35100 28314 35156 28316
rect 35180 28314 35236 28316
rect 34940 28262 34966 28314
rect 34966 28262 34996 28314
rect 35020 28262 35030 28314
rect 35030 28262 35076 28314
rect 35100 28262 35146 28314
rect 35146 28262 35156 28314
rect 35180 28262 35210 28314
rect 35210 28262 35236 28314
rect 34940 28260 34996 28262
rect 35020 28260 35076 28262
rect 35100 28260 35156 28262
rect 35180 28260 35236 28262
rect 34940 27226 34996 27228
rect 35020 27226 35076 27228
rect 35100 27226 35156 27228
rect 35180 27226 35236 27228
rect 34940 27174 34966 27226
rect 34966 27174 34996 27226
rect 35020 27174 35030 27226
rect 35030 27174 35076 27226
rect 35100 27174 35146 27226
rect 35146 27174 35156 27226
rect 35180 27174 35210 27226
rect 35210 27174 35236 27226
rect 34940 27172 34996 27174
rect 35020 27172 35076 27174
rect 35100 27172 35156 27174
rect 35180 27172 35236 27174
rect 34940 26138 34996 26140
rect 35020 26138 35076 26140
rect 35100 26138 35156 26140
rect 35180 26138 35236 26140
rect 34940 26086 34966 26138
rect 34966 26086 34996 26138
rect 35020 26086 35030 26138
rect 35030 26086 35076 26138
rect 35100 26086 35146 26138
rect 35146 26086 35156 26138
rect 35180 26086 35210 26138
rect 35210 26086 35236 26138
rect 34940 26084 34996 26086
rect 35020 26084 35076 26086
rect 35100 26084 35156 26086
rect 35180 26084 35236 26086
rect 34940 25050 34996 25052
rect 35020 25050 35076 25052
rect 35100 25050 35156 25052
rect 35180 25050 35236 25052
rect 34940 24998 34966 25050
rect 34966 24998 34996 25050
rect 35020 24998 35030 25050
rect 35030 24998 35076 25050
rect 35100 24998 35146 25050
rect 35146 24998 35156 25050
rect 35180 24998 35210 25050
rect 35210 24998 35236 25050
rect 34940 24996 34996 24998
rect 35020 24996 35076 24998
rect 35100 24996 35156 24998
rect 35180 24996 35236 24998
rect 34940 23962 34996 23964
rect 35020 23962 35076 23964
rect 35100 23962 35156 23964
rect 35180 23962 35236 23964
rect 34940 23910 34966 23962
rect 34966 23910 34996 23962
rect 35020 23910 35030 23962
rect 35030 23910 35076 23962
rect 35100 23910 35146 23962
rect 35146 23910 35156 23962
rect 35180 23910 35210 23962
rect 35210 23910 35236 23962
rect 34940 23908 34996 23910
rect 35020 23908 35076 23910
rect 35100 23908 35156 23910
rect 35180 23908 35236 23910
rect 34940 22874 34996 22876
rect 35020 22874 35076 22876
rect 35100 22874 35156 22876
rect 35180 22874 35236 22876
rect 34940 22822 34966 22874
rect 34966 22822 34996 22874
rect 35020 22822 35030 22874
rect 35030 22822 35076 22874
rect 35100 22822 35146 22874
rect 35146 22822 35156 22874
rect 35180 22822 35210 22874
rect 35210 22822 35236 22874
rect 34940 22820 34996 22822
rect 35020 22820 35076 22822
rect 35100 22820 35156 22822
rect 35180 22820 35236 22822
rect 31298 6976 31354 7032
rect 31758 6704 31814 6760
rect 31666 6024 31722 6080
rect 32494 8064 32550 8120
rect 32126 6296 32182 6352
rect 31850 5652 31852 5672
rect 31852 5652 31904 5672
rect 31904 5652 31906 5672
rect 31850 5616 31906 5652
rect 31758 4800 31814 4856
rect 31666 4392 31722 4448
rect 31850 4392 31906 4448
rect 32954 8064 33010 8120
rect 32770 7928 32826 7984
rect 32862 6024 32918 6080
rect 34940 21786 34996 21788
rect 35020 21786 35076 21788
rect 35100 21786 35156 21788
rect 35180 21786 35236 21788
rect 34940 21734 34966 21786
rect 34966 21734 34996 21786
rect 35020 21734 35030 21786
rect 35030 21734 35076 21786
rect 35100 21734 35146 21786
rect 35146 21734 35156 21786
rect 35180 21734 35210 21786
rect 35210 21734 35236 21786
rect 34940 21732 34996 21734
rect 35020 21732 35076 21734
rect 35100 21732 35156 21734
rect 35180 21732 35236 21734
rect 34940 20698 34996 20700
rect 35020 20698 35076 20700
rect 35100 20698 35156 20700
rect 35180 20698 35236 20700
rect 34940 20646 34966 20698
rect 34966 20646 34996 20698
rect 35020 20646 35030 20698
rect 35030 20646 35076 20698
rect 35100 20646 35146 20698
rect 35146 20646 35156 20698
rect 35180 20646 35210 20698
rect 35210 20646 35236 20698
rect 34940 20644 34996 20646
rect 35020 20644 35076 20646
rect 35100 20644 35156 20646
rect 35180 20644 35236 20646
rect 34940 19610 34996 19612
rect 35020 19610 35076 19612
rect 35100 19610 35156 19612
rect 35180 19610 35236 19612
rect 34940 19558 34966 19610
rect 34966 19558 34996 19610
rect 35020 19558 35030 19610
rect 35030 19558 35076 19610
rect 35100 19558 35146 19610
rect 35146 19558 35156 19610
rect 35180 19558 35210 19610
rect 35210 19558 35236 19610
rect 34940 19556 34996 19558
rect 35020 19556 35076 19558
rect 35100 19556 35156 19558
rect 35180 19556 35236 19558
rect 34940 18522 34996 18524
rect 35020 18522 35076 18524
rect 35100 18522 35156 18524
rect 35180 18522 35236 18524
rect 34940 18470 34966 18522
rect 34966 18470 34996 18522
rect 35020 18470 35030 18522
rect 35030 18470 35076 18522
rect 35100 18470 35146 18522
rect 35146 18470 35156 18522
rect 35180 18470 35210 18522
rect 35210 18470 35236 18522
rect 34940 18468 34996 18470
rect 35020 18468 35076 18470
rect 35100 18468 35156 18470
rect 35180 18468 35236 18470
rect 34940 17434 34996 17436
rect 35020 17434 35076 17436
rect 35100 17434 35156 17436
rect 35180 17434 35236 17436
rect 34940 17382 34966 17434
rect 34966 17382 34996 17434
rect 35020 17382 35030 17434
rect 35030 17382 35076 17434
rect 35100 17382 35146 17434
rect 35146 17382 35156 17434
rect 35180 17382 35210 17434
rect 35210 17382 35236 17434
rect 34940 17380 34996 17382
rect 35020 17380 35076 17382
rect 35100 17380 35156 17382
rect 35180 17380 35236 17382
rect 34940 16346 34996 16348
rect 35020 16346 35076 16348
rect 35100 16346 35156 16348
rect 35180 16346 35236 16348
rect 34940 16294 34966 16346
rect 34966 16294 34996 16346
rect 35020 16294 35030 16346
rect 35030 16294 35076 16346
rect 35100 16294 35146 16346
rect 35146 16294 35156 16346
rect 35180 16294 35210 16346
rect 35210 16294 35236 16346
rect 34940 16292 34996 16294
rect 35020 16292 35076 16294
rect 35100 16292 35156 16294
rect 35180 16292 35236 16294
rect 33138 6196 33140 6216
rect 33140 6196 33192 6216
rect 33192 6196 33194 6216
rect 33138 6160 33194 6196
rect 33046 5072 33102 5128
rect 33322 6840 33378 6896
rect 34940 15258 34996 15260
rect 35020 15258 35076 15260
rect 35100 15258 35156 15260
rect 35180 15258 35236 15260
rect 34940 15206 34966 15258
rect 34966 15206 34996 15258
rect 35020 15206 35030 15258
rect 35030 15206 35076 15258
rect 35100 15206 35146 15258
rect 35146 15206 35156 15258
rect 35180 15206 35210 15258
rect 35210 15206 35236 15258
rect 34940 15204 34996 15206
rect 35020 15204 35076 15206
rect 35100 15204 35156 15206
rect 35180 15204 35236 15206
rect 50300 116986 50356 116988
rect 50380 116986 50436 116988
rect 50460 116986 50516 116988
rect 50540 116986 50596 116988
rect 50300 116934 50326 116986
rect 50326 116934 50356 116986
rect 50380 116934 50390 116986
rect 50390 116934 50436 116986
rect 50460 116934 50506 116986
rect 50506 116934 50516 116986
rect 50540 116934 50570 116986
rect 50570 116934 50596 116986
rect 50300 116932 50356 116934
rect 50380 116932 50436 116934
rect 50460 116932 50516 116934
rect 50540 116932 50596 116934
rect 50300 115898 50356 115900
rect 50380 115898 50436 115900
rect 50460 115898 50516 115900
rect 50540 115898 50596 115900
rect 50300 115846 50326 115898
rect 50326 115846 50356 115898
rect 50380 115846 50390 115898
rect 50390 115846 50436 115898
rect 50460 115846 50506 115898
rect 50506 115846 50516 115898
rect 50540 115846 50570 115898
rect 50570 115846 50596 115898
rect 50300 115844 50356 115846
rect 50380 115844 50436 115846
rect 50460 115844 50516 115846
rect 50540 115844 50596 115846
rect 50300 114810 50356 114812
rect 50380 114810 50436 114812
rect 50460 114810 50516 114812
rect 50540 114810 50596 114812
rect 50300 114758 50326 114810
rect 50326 114758 50356 114810
rect 50380 114758 50390 114810
rect 50390 114758 50436 114810
rect 50460 114758 50506 114810
rect 50506 114758 50516 114810
rect 50540 114758 50570 114810
rect 50570 114758 50596 114810
rect 50300 114756 50356 114758
rect 50380 114756 50436 114758
rect 50460 114756 50516 114758
rect 50540 114756 50596 114758
rect 50300 113722 50356 113724
rect 50380 113722 50436 113724
rect 50460 113722 50516 113724
rect 50540 113722 50596 113724
rect 50300 113670 50326 113722
rect 50326 113670 50356 113722
rect 50380 113670 50390 113722
rect 50390 113670 50436 113722
rect 50460 113670 50506 113722
rect 50506 113670 50516 113722
rect 50540 113670 50570 113722
rect 50570 113670 50596 113722
rect 50300 113668 50356 113670
rect 50380 113668 50436 113670
rect 50460 113668 50516 113670
rect 50540 113668 50596 113670
rect 50300 112634 50356 112636
rect 50380 112634 50436 112636
rect 50460 112634 50516 112636
rect 50540 112634 50596 112636
rect 50300 112582 50326 112634
rect 50326 112582 50356 112634
rect 50380 112582 50390 112634
rect 50390 112582 50436 112634
rect 50460 112582 50506 112634
rect 50506 112582 50516 112634
rect 50540 112582 50570 112634
rect 50570 112582 50596 112634
rect 50300 112580 50356 112582
rect 50380 112580 50436 112582
rect 50460 112580 50516 112582
rect 50540 112580 50596 112582
rect 50300 111546 50356 111548
rect 50380 111546 50436 111548
rect 50460 111546 50516 111548
rect 50540 111546 50596 111548
rect 50300 111494 50326 111546
rect 50326 111494 50356 111546
rect 50380 111494 50390 111546
rect 50390 111494 50436 111546
rect 50460 111494 50506 111546
rect 50506 111494 50516 111546
rect 50540 111494 50570 111546
rect 50570 111494 50596 111546
rect 50300 111492 50356 111494
rect 50380 111492 50436 111494
rect 50460 111492 50516 111494
rect 50540 111492 50596 111494
rect 50300 110458 50356 110460
rect 50380 110458 50436 110460
rect 50460 110458 50516 110460
rect 50540 110458 50596 110460
rect 50300 110406 50326 110458
rect 50326 110406 50356 110458
rect 50380 110406 50390 110458
rect 50390 110406 50436 110458
rect 50460 110406 50506 110458
rect 50506 110406 50516 110458
rect 50540 110406 50570 110458
rect 50570 110406 50596 110458
rect 50300 110404 50356 110406
rect 50380 110404 50436 110406
rect 50460 110404 50516 110406
rect 50540 110404 50596 110406
rect 50300 109370 50356 109372
rect 50380 109370 50436 109372
rect 50460 109370 50516 109372
rect 50540 109370 50596 109372
rect 50300 109318 50326 109370
rect 50326 109318 50356 109370
rect 50380 109318 50390 109370
rect 50390 109318 50436 109370
rect 50460 109318 50506 109370
rect 50506 109318 50516 109370
rect 50540 109318 50570 109370
rect 50570 109318 50596 109370
rect 50300 109316 50356 109318
rect 50380 109316 50436 109318
rect 50460 109316 50516 109318
rect 50540 109316 50596 109318
rect 50300 108282 50356 108284
rect 50380 108282 50436 108284
rect 50460 108282 50516 108284
rect 50540 108282 50596 108284
rect 50300 108230 50326 108282
rect 50326 108230 50356 108282
rect 50380 108230 50390 108282
rect 50390 108230 50436 108282
rect 50460 108230 50506 108282
rect 50506 108230 50516 108282
rect 50540 108230 50570 108282
rect 50570 108230 50596 108282
rect 50300 108228 50356 108230
rect 50380 108228 50436 108230
rect 50460 108228 50516 108230
rect 50540 108228 50596 108230
rect 50300 107194 50356 107196
rect 50380 107194 50436 107196
rect 50460 107194 50516 107196
rect 50540 107194 50596 107196
rect 50300 107142 50326 107194
rect 50326 107142 50356 107194
rect 50380 107142 50390 107194
rect 50390 107142 50436 107194
rect 50460 107142 50506 107194
rect 50506 107142 50516 107194
rect 50540 107142 50570 107194
rect 50570 107142 50596 107194
rect 50300 107140 50356 107142
rect 50380 107140 50436 107142
rect 50460 107140 50516 107142
rect 50540 107140 50596 107142
rect 50300 106106 50356 106108
rect 50380 106106 50436 106108
rect 50460 106106 50516 106108
rect 50540 106106 50596 106108
rect 50300 106054 50326 106106
rect 50326 106054 50356 106106
rect 50380 106054 50390 106106
rect 50390 106054 50436 106106
rect 50460 106054 50506 106106
rect 50506 106054 50516 106106
rect 50540 106054 50570 106106
rect 50570 106054 50596 106106
rect 50300 106052 50356 106054
rect 50380 106052 50436 106054
rect 50460 106052 50516 106054
rect 50540 106052 50596 106054
rect 50300 105018 50356 105020
rect 50380 105018 50436 105020
rect 50460 105018 50516 105020
rect 50540 105018 50596 105020
rect 50300 104966 50326 105018
rect 50326 104966 50356 105018
rect 50380 104966 50390 105018
rect 50390 104966 50436 105018
rect 50460 104966 50506 105018
rect 50506 104966 50516 105018
rect 50540 104966 50570 105018
rect 50570 104966 50596 105018
rect 50300 104964 50356 104966
rect 50380 104964 50436 104966
rect 50460 104964 50516 104966
rect 50540 104964 50596 104966
rect 50300 103930 50356 103932
rect 50380 103930 50436 103932
rect 50460 103930 50516 103932
rect 50540 103930 50596 103932
rect 50300 103878 50326 103930
rect 50326 103878 50356 103930
rect 50380 103878 50390 103930
rect 50390 103878 50436 103930
rect 50460 103878 50506 103930
rect 50506 103878 50516 103930
rect 50540 103878 50570 103930
rect 50570 103878 50596 103930
rect 50300 103876 50356 103878
rect 50380 103876 50436 103878
rect 50460 103876 50516 103878
rect 50540 103876 50596 103878
rect 50300 102842 50356 102844
rect 50380 102842 50436 102844
rect 50460 102842 50516 102844
rect 50540 102842 50596 102844
rect 50300 102790 50326 102842
rect 50326 102790 50356 102842
rect 50380 102790 50390 102842
rect 50390 102790 50436 102842
rect 50460 102790 50506 102842
rect 50506 102790 50516 102842
rect 50540 102790 50570 102842
rect 50570 102790 50596 102842
rect 50300 102788 50356 102790
rect 50380 102788 50436 102790
rect 50460 102788 50516 102790
rect 50540 102788 50596 102790
rect 50300 101754 50356 101756
rect 50380 101754 50436 101756
rect 50460 101754 50516 101756
rect 50540 101754 50596 101756
rect 50300 101702 50326 101754
rect 50326 101702 50356 101754
rect 50380 101702 50390 101754
rect 50390 101702 50436 101754
rect 50460 101702 50506 101754
rect 50506 101702 50516 101754
rect 50540 101702 50570 101754
rect 50570 101702 50596 101754
rect 50300 101700 50356 101702
rect 50380 101700 50436 101702
rect 50460 101700 50516 101702
rect 50540 101700 50596 101702
rect 50300 100666 50356 100668
rect 50380 100666 50436 100668
rect 50460 100666 50516 100668
rect 50540 100666 50596 100668
rect 50300 100614 50326 100666
rect 50326 100614 50356 100666
rect 50380 100614 50390 100666
rect 50390 100614 50436 100666
rect 50460 100614 50506 100666
rect 50506 100614 50516 100666
rect 50540 100614 50570 100666
rect 50570 100614 50596 100666
rect 50300 100612 50356 100614
rect 50380 100612 50436 100614
rect 50460 100612 50516 100614
rect 50540 100612 50596 100614
rect 50300 99578 50356 99580
rect 50380 99578 50436 99580
rect 50460 99578 50516 99580
rect 50540 99578 50596 99580
rect 50300 99526 50326 99578
rect 50326 99526 50356 99578
rect 50380 99526 50390 99578
rect 50390 99526 50436 99578
rect 50460 99526 50506 99578
rect 50506 99526 50516 99578
rect 50540 99526 50570 99578
rect 50570 99526 50596 99578
rect 50300 99524 50356 99526
rect 50380 99524 50436 99526
rect 50460 99524 50516 99526
rect 50540 99524 50596 99526
rect 50300 98490 50356 98492
rect 50380 98490 50436 98492
rect 50460 98490 50516 98492
rect 50540 98490 50596 98492
rect 50300 98438 50326 98490
rect 50326 98438 50356 98490
rect 50380 98438 50390 98490
rect 50390 98438 50436 98490
rect 50460 98438 50506 98490
rect 50506 98438 50516 98490
rect 50540 98438 50570 98490
rect 50570 98438 50596 98490
rect 50300 98436 50356 98438
rect 50380 98436 50436 98438
rect 50460 98436 50516 98438
rect 50540 98436 50596 98438
rect 50300 97402 50356 97404
rect 50380 97402 50436 97404
rect 50460 97402 50516 97404
rect 50540 97402 50596 97404
rect 50300 97350 50326 97402
rect 50326 97350 50356 97402
rect 50380 97350 50390 97402
rect 50390 97350 50436 97402
rect 50460 97350 50506 97402
rect 50506 97350 50516 97402
rect 50540 97350 50570 97402
rect 50570 97350 50596 97402
rect 50300 97348 50356 97350
rect 50380 97348 50436 97350
rect 50460 97348 50516 97350
rect 50540 97348 50596 97350
rect 50300 96314 50356 96316
rect 50380 96314 50436 96316
rect 50460 96314 50516 96316
rect 50540 96314 50596 96316
rect 50300 96262 50326 96314
rect 50326 96262 50356 96314
rect 50380 96262 50390 96314
rect 50390 96262 50436 96314
rect 50460 96262 50506 96314
rect 50506 96262 50516 96314
rect 50540 96262 50570 96314
rect 50570 96262 50596 96314
rect 50300 96260 50356 96262
rect 50380 96260 50436 96262
rect 50460 96260 50516 96262
rect 50540 96260 50596 96262
rect 50300 95226 50356 95228
rect 50380 95226 50436 95228
rect 50460 95226 50516 95228
rect 50540 95226 50596 95228
rect 50300 95174 50326 95226
rect 50326 95174 50356 95226
rect 50380 95174 50390 95226
rect 50390 95174 50436 95226
rect 50460 95174 50506 95226
rect 50506 95174 50516 95226
rect 50540 95174 50570 95226
rect 50570 95174 50596 95226
rect 50300 95172 50356 95174
rect 50380 95172 50436 95174
rect 50460 95172 50516 95174
rect 50540 95172 50596 95174
rect 50300 94138 50356 94140
rect 50380 94138 50436 94140
rect 50460 94138 50516 94140
rect 50540 94138 50596 94140
rect 50300 94086 50326 94138
rect 50326 94086 50356 94138
rect 50380 94086 50390 94138
rect 50390 94086 50436 94138
rect 50460 94086 50506 94138
rect 50506 94086 50516 94138
rect 50540 94086 50570 94138
rect 50570 94086 50596 94138
rect 50300 94084 50356 94086
rect 50380 94084 50436 94086
rect 50460 94084 50516 94086
rect 50540 94084 50596 94086
rect 50300 93050 50356 93052
rect 50380 93050 50436 93052
rect 50460 93050 50516 93052
rect 50540 93050 50596 93052
rect 50300 92998 50326 93050
rect 50326 92998 50356 93050
rect 50380 92998 50390 93050
rect 50390 92998 50436 93050
rect 50460 92998 50506 93050
rect 50506 92998 50516 93050
rect 50540 92998 50570 93050
rect 50570 92998 50596 93050
rect 50300 92996 50356 92998
rect 50380 92996 50436 92998
rect 50460 92996 50516 92998
rect 50540 92996 50596 92998
rect 50300 91962 50356 91964
rect 50380 91962 50436 91964
rect 50460 91962 50516 91964
rect 50540 91962 50596 91964
rect 50300 91910 50326 91962
rect 50326 91910 50356 91962
rect 50380 91910 50390 91962
rect 50390 91910 50436 91962
rect 50460 91910 50506 91962
rect 50506 91910 50516 91962
rect 50540 91910 50570 91962
rect 50570 91910 50596 91962
rect 50300 91908 50356 91910
rect 50380 91908 50436 91910
rect 50460 91908 50516 91910
rect 50540 91908 50596 91910
rect 50300 90874 50356 90876
rect 50380 90874 50436 90876
rect 50460 90874 50516 90876
rect 50540 90874 50596 90876
rect 50300 90822 50326 90874
rect 50326 90822 50356 90874
rect 50380 90822 50390 90874
rect 50390 90822 50436 90874
rect 50460 90822 50506 90874
rect 50506 90822 50516 90874
rect 50540 90822 50570 90874
rect 50570 90822 50596 90874
rect 50300 90820 50356 90822
rect 50380 90820 50436 90822
rect 50460 90820 50516 90822
rect 50540 90820 50596 90822
rect 50300 89786 50356 89788
rect 50380 89786 50436 89788
rect 50460 89786 50516 89788
rect 50540 89786 50596 89788
rect 50300 89734 50326 89786
rect 50326 89734 50356 89786
rect 50380 89734 50390 89786
rect 50390 89734 50436 89786
rect 50460 89734 50506 89786
rect 50506 89734 50516 89786
rect 50540 89734 50570 89786
rect 50570 89734 50596 89786
rect 50300 89732 50356 89734
rect 50380 89732 50436 89734
rect 50460 89732 50516 89734
rect 50540 89732 50596 89734
rect 50300 88698 50356 88700
rect 50380 88698 50436 88700
rect 50460 88698 50516 88700
rect 50540 88698 50596 88700
rect 50300 88646 50326 88698
rect 50326 88646 50356 88698
rect 50380 88646 50390 88698
rect 50390 88646 50436 88698
rect 50460 88646 50506 88698
rect 50506 88646 50516 88698
rect 50540 88646 50570 88698
rect 50570 88646 50596 88698
rect 50300 88644 50356 88646
rect 50380 88644 50436 88646
rect 50460 88644 50516 88646
rect 50540 88644 50596 88646
rect 50300 87610 50356 87612
rect 50380 87610 50436 87612
rect 50460 87610 50516 87612
rect 50540 87610 50596 87612
rect 50300 87558 50326 87610
rect 50326 87558 50356 87610
rect 50380 87558 50390 87610
rect 50390 87558 50436 87610
rect 50460 87558 50506 87610
rect 50506 87558 50516 87610
rect 50540 87558 50570 87610
rect 50570 87558 50596 87610
rect 50300 87556 50356 87558
rect 50380 87556 50436 87558
rect 50460 87556 50516 87558
rect 50540 87556 50596 87558
rect 50300 86522 50356 86524
rect 50380 86522 50436 86524
rect 50460 86522 50516 86524
rect 50540 86522 50596 86524
rect 50300 86470 50326 86522
rect 50326 86470 50356 86522
rect 50380 86470 50390 86522
rect 50390 86470 50436 86522
rect 50460 86470 50506 86522
rect 50506 86470 50516 86522
rect 50540 86470 50570 86522
rect 50570 86470 50596 86522
rect 50300 86468 50356 86470
rect 50380 86468 50436 86470
rect 50460 86468 50516 86470
rect 50540 86468 50596 86470
rect 50300 85434 50356 85436
rect 50380 85434 50436 85436
rect 50460 85434 50516 85436
rect 50540 85434 50596 85436
rect 50300 85382 50326 85434
rect 50326 85382 50356 85434
rect 50380 85382 50390 85434
rect 50390 85382 50436 85434
rect 50460 85382 50506 85434
rect 50506 85382 50516 85434
rect 50540 85382 50570 85434
rect 50570 85382 50596 85434
rect 50300 85380 50356 85382
rect 50380 85380 50436 85382
rect 50460 85380 50516 85382
rect 50540 85380 50596 85382
rect 50300 84346 50356 84348
rect 50380 84346 50436 84348
rect 50460 84346 50516 84348
rect 50540 84346 50596 84348
rect 50300 84294 50326 84346
rect 50326 84294 50356 84346
rect 50380 84294 50390 84346
rect 50390 84294 50436 84346
rect 50460 84294 50506 84346
rect 50506 84294 50516 84346
rect 50540 84294 50570 84346
rect 50570 84294 50596 84346
rect 50300 84292 50356 84294
rect 50380 84292 50436 84294
rect 50460 84292 50516 84294
rect 50540 84292 50596 84294
rect 50300 83258 50356 83260
rect 50380 83258 50436 83260
rect 50460 83258 50516 83260
rect 50540 83258 50596 83260
rect 50300 83206 50326 83258
rect 50326 83206 50356 83258
rect 50380 83206 50390 83258
rect 50390 83206 50436 83258
rect 50460 83206 50506 83258
rect 50506 83206 50516 83258
rect 50540 83206 50570 83258
rect 50570 83206 50596 83258
rect 50300 83204 50356 83206
rect 50380 83204 50436 83206
rect 50460 83204 50516 83206
rect 50540 83204 50596 83206
rect 50300 82170 50356 82172
rect 50380 82170 50436 82172
rect 50460 82170 50516 82172
rect 50540 82170 50596 82172
rect 50300 82118 50326 82170
rect 50326 82118 50356 82170
rect 50380 82118 50390 82170
rect 50390 82118 50436 82170
rect 50460 82118 50506 82170
rect 50506 82118 50516 82170
rect 50540 82118 50570 82170
rect 50570 82118 50596 82170
rect 50300 82116 50356 82118
rect 50380 82116 50436 82118
rect 50460 82116 50516 82118
rect 50540 82116 50596 82118
rect 50300 81082 50356 81084
rect 50380 81082 50436 81084
rect 50460 81082 50516 81084
rect 50540 81082 50596 81084
rect 50300 81030 50326 81082
rect 50326 81030 50356 81082
rect 50380 81030 50390 81082
rect 50390 81030 50436 81082
rect 50460 81030 50506 81082
rect 50506 81030 50516 81082
rect 50540 81030 50570 81082
rect 50570 81030 50596 81082
rect 50300 81028 50356 81030
rect 50380 81028 50436 81030
rect 50460 81028 50516 81030
rect 50540 81028 50596 81030
rect 50300 79994 50356 79996
rect 50380 79994 50436 79996
rect 50460 79994 50516 79996
rect 50540 79994 50596 79996
rect 50300 79942 50326 79994
rect 50326 79942 50356 79994
rect 50380 79942 50390 79994
rect 50390 79942 50436 79994
rect 50460 79942 50506 79994
rect 50506 79942 50516 79994
rect 50540 79942 50570 79994
rect 50570 79942 50596 79994
rect 50300 79940 50356 79942
rect 50380 79940 50436 79942
rect 50460 79940 50516 79942
rect 50540 79940 50596 79942
rect 50300 78906 50356 78908
rect 50380 78906 50436 78908
rect 50460 78906 50516 78908
rect 50540 78906 50596 78908
rect 50300 78854 50326 78906
rect 50326 78854 50356 78906
rect 50380 78854 50390 78906
rect 50390 78854 50436 78906
rect 50460 78854 50506 78906
rect 50506 78854 50516 78906
rect 50540 78854 50570 78906
rect 50570 78854 50596 78906
rect 50300 78852 50356 78854
rect 50380 78852 50436 78854
rect 50460 78852 50516 78854
rect 50540 78852 50596 78854
rect 50300 77818 50356 77820
rect 50380 77818 50436 77820
rect 50460 77818 50516 77820
rect 50540 77818 50596 77820
rect 50300 77766 50326 77818
rect 50326 77766 50356 77818
rect 50380 77766 50390 77818
rect 50390 77766 50436 77818
rect 50460 77766 50506 77818
rect 50506 77766 50516 77818
rect 50540 77766 50570 77818
rect 50570 77766 50596 77818
rect 50300 77764 50356 77766
rect 50380 77764 50436 77766
rect 50460 77764 50516 77766
rect 50540 77764 50596 77766
rect 50300 76730 50356 76732
rect 50380 76730 50436 76732
rect 50460 76730 50516 76732
rect 50540 76730 50596 76732
rect 50300 76678 50326 76730
rect 50326 76678 50356 76730
rect 50380 76678 50390 76730
rect 50390 76678 50436 76730
rect 50460 76678 50506 76730
rect 50506 76678 50516 76730
rect 50540 76678 50570 76730
rect 50570 76678 50596 76730
rect 50300 76676 50356 76678
rect 50380 76676 50436 76678
rect 50460 76676 50516 76678
rect 50540 76676 50596 76678
rect 50300 75642 50356 75644
rect 50380 75642 50436 75644
rect 50460 75642 50516 75644
rect 50540 75642 50596 75644
rect 50300 75590 50326 75642
rect 50326 75590 50356 75642
rect 50380 75590 50390 75642
rect 50390 75590 50436 75642
rect 50460 75590 50506 75642
rect 50506 75590 50516 75642
rect 50540 75590 50570 75642
rect 50570 75590 50596 75642
rect 50300 75588 50356 75590
rect 50380 75588 50436 75590
rect 50460 75588 50516 75590
rect 50540 75588 50596 75590
rect 50300 74554 50356 74556
rect 50380 74554 50436 74556
rect 50460 74554 50516 74556
rect 50540 74554 50596 74556
rect 50300 74502 50326 74554
rect 50326 74502 50356 74554
rect 50380 74502 50390 74554
rect 50390 74502 50436 74554
rect 50460 74502 50506 74554
rect 50506 74502 50516 74554
rect 50540 74502 50570 74554
rect 50570 74502 50596 74554
rect 50300 74500 50356 74502
rect 50380 74500 50436 74502
rect 50460 74500 50516 74502
rect 50540 74500 50596 74502
rect 50300 73466 50356 73468
rect 50380 73466 50436 73468
rect 50460 73466 50516 73468
rect 50540 73466 50596 73468
rect 50300 73414 50326 73466
rect 50326 73414 50356 73466
rect 50380 73414 50390 73466
rect 50390 73414 50436 73466
rect 50460 73414 50506 73466
rect 50506 73414 50516 73466
rect 50540 73414 50570 73466
rect 50570 73414 50596 73466
rect 50300 73412 50356 73414
rect 50380 73412 50436 73414
rect 50460 73412 50516 73414
rect 50540 73412 50596 73414
rect 50300 72378 50356 72380
rect 50380 72378 50436 72380
rect 50460 72378 50516 72380
rect 50540 72378 50596 72380
rect 50300 72326 50326 72378
rect 50326 72326 50356 72378
rect 50380 72326 50390 72378
rect 50390 72326 50436 72378
rect 50460 72326 50506 72378
rect 50506 72326 50516 72378
rect 50540 72326 50570 72378
rect 50570 72326 50596 72378
rect 50300 72324 50356 72326
rect 50380 72324 50436 72326
rect 50460 72324 50516 72326
rect 50540 72324 50596 72326
rect 50300 71290 50356 71292
rect 50380 71290 50436 71292
rect 50460 71290 50516 71292
rect 50540 71290 50596 71292
rect 50300 71238 50326 71290
rect 50326 71238 50356 71290
rect 50380 71238 50390 71290
rect 50390 71238 50436 71290
rect 50460 71238 50506 71290
rect 50506 71238 50516 71290
rect 50540 71238 50570 71290
rect 50570 71238 50596 71290
rect 50300 71236 50356 71238
rect 50380 71236 50436 71238
rect 50460 71236 50516 71238
rect 50540 71236 50596 71238
rect 50300 70202 50356 70204
rect 50380 70202 50436 70204
rect 50460 70202 50516 70204
rect 50540 70202 50596 70204
rect 50300 70150 50326 70202
rect 50326 70150 50356 70202
rect 50380 70150 50390 70202
rect 50390 70150 50436 70202
rect 50460 70150 50506 70202
rect 50506 70150 50516 70202
rect 50540 70150 50570 70202
rect 50570 70150 50596 70202
rect 50300 70148 50356 70150
rect 50380 70148 50436 70150
rect 50460 70148 50516 70150
rect 50540 70148 50596 70150
rect 50300 69114 50356 69116
rect 50380 69114 50436 69116
rect 50460 69114 50516 69116
rect 50540 69114 50596 69116
rect 50300 69062 50326 69114
rect 50326 69062 50356 69114
rect 50380 69062 50390 69114
rect 50390 69062 50436 69114
rect 50460 69062 50506 69114
rect 50506 69062 50516 69114
rect 50540 69062 50570 69114
rect 50570 69062 50596 69114
rect 50300 69060 50356 69062
rect 50380 69060 50436 69062
rect 50460 69060 50516 69062
rect 50540 69060 50596 69062
rect 50300 68026 50356 68028
rect 50380 68026 50436 68028
rect 50460 68026 50516 68028
rect 50540 68026 50596 68028
rect 50300 67974 50326 68026
rect 50326 67974 50356 68026
rect 50380 67974 50390 68026
rect 50390 67974 50436 68026
rect 50460 67974 50506 68026
rect 50506 67974 50516 68026
rect 50540 67974 50570 68026
rect 50570 67974 50596 68026
rect 50300 67972 50356 67974
rect 50380 67972 50436 67974
rect 50460 67972 50516 67974
rect 50540 67972 50596 67974
rect 50300 66938 50356 66940
rect 50380 66938 50436 66940
rect 50460 66938 50516 66940
rect 50540 66938 50596 66940
rect 50300 66886 50326 66938
rect 50326 66886 50356 66938
rect 50380 66886 50390 66938
rect 50390 66886 50436 66938
rect 50460 66886 50506 66938
rect 50506 66886 50516 66938
rect 50540 66886 50570 66938
rect 50570 66886 50596 66938
rect 50300 66884 50356 66886
rect 50380 66884 50436 66886
rect 50460 66884 50516 66886
rect 50540 66884 50596 66886
rect 50300 65850 50356 65852
rect 50380 65850 50436 65852
rect 50460 65850 50516 65852
rect 50540 65850 50596 65852
rect 50300 65798 50326 65850
rect 50326 65798 50356 65850
rect 50380 65798 50390 65850
rect 50390 65798 50436 65850
rect 50460 65798 50506 65850
rect 50506 65798 50516 65850
rect 50540 65798 50570 65850
rect 50570 65798 50596 65850
rect 50300 65796 50356 65798
rect 50380 65796 50436 65798
rect 50460 65796 50516 65798
rect 50540 65796 50596 65798
rect 50300 64762 50356 64764
rect 50380 64762 50436 64764
rect 50460 64762 50516 64764
rect 50540 64762 50596 64764
rect 50300 64710 50326 64762
rect 50326 64710 50356 64762
rect 50380 64710 50390 64762
rect 50390 64710 50436 64762
rect 50460 64710 50506 64762
rect 50506 64710 50516 64762
rect 50540 64710 50570 64762
rect 50570 64710 50596 64762
rect 50300 64708 50356 64710
rect 50380 64708 50436 64710
rect 50460 64708 50516 64710
rect 50540 64708 50596 64710
rect 50300 63674 50356 63676
rect 50380 63674 50436 63676
rect 50460 63674 50516 63676
rect 50540 63674 50596 63676
rect 50300 63622 50326 63674
rect 50326 63622 50356 63674
rect 50380 63622 50390 63674
rect 50390 63622 50436 63674
rect 50460 63622 50506 63674
rect 50506 63622 50516 63674
rect 50540 63622 50570 63674
rect 50570 63622 50596 63674
rect 50300 63620 50356 63622
rect 50380 63620 50436 63622
rect 50460 63620 50516 63622
rect 50540 63620 50596 63622
rect 50300 62586 50356 62588
rect 50380 62586 50436 62588
rect 50460 62586 50516 62588
rect 50540 62586 50596 62588
rect 50300 62534 50326 62586
rect 50326 62534 50356 62586
rect 50380 62534 50390 62586
rect 50390 62534 50436 62586
rect 50460 62534 50506 62586
rect 50506 62534 50516 62586
rect 50540 62534 50570 62586
rect 50570 62534 50596 62586
rect 50300 62532 50356 62534
rect 50380 62532 50436 62534
rect 50460 62532 50516 62534
rect 50540 62532 50596 62534
rect 50300 61498 50356 61500
rect 50380 61498 50436 61500
rect 50460 61498 50516 61500
rect 50540 61498 50596 61500
rect 50300 61446 50326 61498
rect 50326 61446 50356 61498
rect 50380 61446 50390 61498
rect 50390 61446 50436 61498
rect 50460 61446 50506 61498
rect 50506 61446 50516 61498
rect 50540 61446 50570 61498
rect 50570 61446 50596 61498
rect 50300 61444 50356 61446
rect 50380 61444 50436 61446
rect 50460 61444 50516 61446
rect 50540 61444 50596 61446
rect 50300 60410 50356 60412
rect 50380 60410 50436 60412
rect 50460 60410 50516 60412
rect 50540 60410 50596 60412
rect 50300 60358 50326 60410
rect 50326 60358 50356 60410
rect 50380 60358 50390 60410
rect 50390 60358 50436 60410
rect 50460 60358 50506 60410
rect 50506 60358 50516 60410
rect 50540 60358 50570 60410
rect 50570 60358 50596 60410
rect 50300 60356 50356 60358
rect 50380 60356 50436 60358
rect 50460 60356 50516 60358
rect 50540 60356 50596 60358
rect 50300 59322 50356 59324
rect 50380 59322 50436 59324
rect 50460 59322 50516 59324
rect 50540 59322 50596 59324
rect 50300 59270 50326 59322
rect 50326 59270 50356 59322
rect 50380 59270 50390 59322
rect 50390 59270 50436 59322
rect 50460 59270 50506 59322
rect 50506 59270 50516 59322
rect 50540 59270 50570 59322
rect 50570 59270 50596 59322
rect 50300 59268 50356 59270
rect 50380 59268 50436 59270
rect 50460 59268 50516 59270
rect 50540 59268 50596 59270
rect 50300 58234 50356 58236
rect 50380 58234 50436 58236
rect 50460 58234 50516 58236
rect 50540 58234 50596 58236
rect 50300 58182 50326 58234
rect 50326 58182 50356 58234
rect 50380 58182 50390 58234
rect 50390 58182 50436 58234
rect 50460 58182 50506 58234
rect 50506 58182 50516 58234
rect 50540 58182 50570 58234
rect 50570 58182 50596 58234
rect 50300 58180 50356 58182
rect 50380 58180 50436 58182
rect 50460 58180 50516 58182
rect 50540 58180 50596 58182
rect 50300 57146 50356 57148
rect 50380 57146 50436 57148
rect 50460 57146 50516 57148
rect 50540 57146 50596 57148
rect 50300 57094 50326 57146
rect 50326 57094 50356 57146
rect 50380 57094 50390 57146
rect 50390 57094 50436 57146
rect 50460 57094 50506 57146
rect 50506 57094 50516 57146
rect 50540 57094 50570 57146
rect 50570 57094 50596 57146
rect 50300 57092 50356 57094
rect 50380 57092 50436 57094
rect 50460 57092 50516 57094
rect 50540 57092 50596 57094
rect 50300 56058 50356 56060
rect 50380 56058 50436 56060
rect 50460 56058 50516 56060
rect 50540 56058 50596 56060
rect 50300 56006 50326 56058
rect 50326 56006 50356 56058
rect 50380 56006 50390 56058
rect 50390 56006 50436 56058
rect 50460 56006 50506 56058
rect 50506 56006 50516 56058
rect 50540 56006 50570 56058
rect 50570 56006 50596 56058
rect 50300 56004 50356 56006
rect 50380 56004 50436 56006
rect 50460 56004 50516 56006
rect 50540 56004 50596 56006
rect 50300 54970 50356 54972
rect 50380 54970 50436 54972
rect 50460 54970 50516 54972
rect 50540 54970 50596 54972
rect 50300 54918 50326 54970
rect 50326 54918 50356 54970
rect 50380 54918 50390 54970
rect 50390 54918 50436 54970
rect 50460 54918 50506 54970
rect 50506 54918 50516 54970
rect 50540 54918 50570 54970
rect 50570 54918 50596 54970
rect 50300 54916 50356 54918
rect 50380 54916 50436 54918
rect 50460 54916 50516 54918
rect 50540 54916 50596 54918
rect 50300 53882 50356 53884
rect 50380 53882 50436 53884
rect 50460 53882 50516 53884
rect 50540 53882 50596 53884
rect 50300 53830 50326 53882
rect 50326 53830 50356 53882
rect 50380 53830 50390 53882
rect 50390 53830 50436 53882
rect 50460 53830 50506 53882
rect 50506 53830 50516 53882
rect 50540 53830 50570 53882
rect 50570 53830 50596 53882
rect 50300 53828 50356 53830
rect 50380 53828 50436 53830
rect 50460 53828 50516 53830
rect 50540 53828 50596 53830
rect 50300 52794 50356 52796
rect 50380 52794 50436 52796
rect 50460 52794 50516 52796
rect 50540 52794 50596 52796
rect 50300 52742 50326 52794
rect 50326 52742 50356 52794
rect 50380 52742 50390 52794
rect 50390 52742 50436 52794
rect 50460 52742 50506 52794
rect 50506 52742 50516 52794
rect 50540 52742 50570 52794
rect 50570 52742 50596 52794
rect 50300 52740 50356 52742
rect 50380 52740 50436 52742
rect 50460 52740 50516 52742
rect 50540 52740 50596 52742
rect 50300 51706 50356 51708
rect 50380 51706 50436 51708
rect 50460 51706 50516 51708
rect 50540 51706 50596 51708
rect 50300 51654 50326 51706
rect 50326 51654 50356 51706
rect 50380 51654 50390 51706
rect 50390 51654 50436 51706
rect 50460 51654 50506 51706
rect 50506 51654 50516 51706
rect 50540 51654 50570 51706
rect 50570 51654 50596 51706
rect 50300 51652 50356 51654
rect 50380 51652 50436 51654
rect 50460 51652 50516 51654
rect 50540 51652 50596 51654
rect 50300 50618 50356 50620
rect 50380 50618 50436 50620
rect 50460 50618 50516 50620
rect 50540 50618 50596 50620
rect 50300 50566 50326 50618
rect 50326 50566 50356 50618
rect 50380 50566 50390 50618
rect 50390 50566 50436 50618
rect 50460 50566 50506 50618
rect 50506 50566 50516 50618
rect 50540 50566 50570 50618
rect 50570 50566 50596 50618
rect 50300 50564 50356 50566
rect 50380 50564 50436 50566
rect 50460 50564 50516 50566
rect 50540 50564 50596 50566
rect 50300 49530 50356 49532
rect 50380 49530 50436 49532
rect 50460 49530 50516 49532
rect 50540 49530 50596 49532
rect 50300 49478 50326 49530
rect 50326 49478 50356 49530
rect 50380 49478 50390 49530
rect 50390 49478 50436 49530
rect 50460 49478 50506 49530
rect 50506 49478 50516 49530
rect 50540 49478 50570 49530
rect 50570 49478 50596 49530
rect 50300 49476 50356 49478
rect 50380 49476 50436 49478
rect 50460 49476 50516 49478
rect 50540 49476 50596 49478
rect 50300 48442 50356 48444
rect 50380 48442 50436 48444
rect 50460 48442 50516 48444
rect 50540 48442 50596 48444
rect 50300 48390 50326 48442
rect 50326 48390 50356 48442
rect 50380 48390 50390 48442
rect 50390 48390 50436 48442
rect 50460 48390 50506 48442
rect 50506 48390 50516 48442
rect 50540 48390 50570 48442
rect 50570 48390 50596 48442
rect 50300 48388 50356 48390
rect 50380 48388 50436 48390
rect 50460 48388 50516 48390
rect 50540 48388 50596 48390
rect 50300 47354 50356 47356
rect 50380 47354 50436 47356
rect 50460 47354 50516 47356
rect 50540 47354 50596 47356
rect 50300 47302 50326 47354
rect 50326 47302 50356 47354
rect 50380 47302 50390 47354
rect 50390 47302 50436 47354
rect 50460 47302 50506 47354
rect 50506 47302 50516 47354
rect 50540 47302 50570 47354
rect 50570 47302 50596 47354
rect 50300 47300 50356 47302
rect 50380 47300 50436 47302
rect 50460 47300 50516 47302
rect 50540 47300 50596 47302
rect 50300 46266 50356 46268
rect 50380 46266 50436 46268
rect 50460 46266 50516 46268
rect 50540 46266 50596 46268
rect 50300 46214 50326 46266
rect 50326 46214 50356 46266
rect 50380 46214 50390 46266
rect 50390 46214 50436 46266
rect 50460 46214 50506 46266
rect 50506 46214 50516 46266
rect 50540 46214 50570 46266
rect 50570 46214 50596 46266
rect 50300 46212 50356 46214
rect 50380 46212 50436 46214
rect 50460 46212 50516 46214
rect 50540 46212 50596 46214
rect 50300 45178 50356 45180
rect 50380 45178 50436 45180
rect 50460 45178 50516 45180
rect 50540 45178 50596 45180
rect 50300 45126 50326 45178
rect 50326 45126 50356 45178
rect 50380 45126 50390 45178
rect 50390 45126 50436 45178
rect 50460 45126 50506 45178
rect 50506 45126 50516 45178
rect 50540 45126 50570 45178
rect 50570 45126 50596 45178
rect 50300 45124 50356 45126
rect 50380 45124 50436 45126
rect 50460 45124 50516 45126
rect 50540 45124 50596 45126
rect 50300 44090 50356 44092
rect 50380 44090 50436 44092
rect 50460 44090 50516 44092
rect 50540 44090 50596 44092
rect 50300 44038 50326 44090
rect 50326 44038 50356 44090
rect 50380 44038 50390 44090
rect 50390 44038 50436 44090
rect 50460 44038 50506 44090
rect 50506 44038 50516 44090
rect 50540 44038 50570 44090
rect 50570 44038 50596 44090
rect 50300 44036 50356 44038
rect 50380 44036 50436 44038
rect 50460 44036 50516 44038
rect 50540 44036 50596 44038
rect 50300 43002 50356 43004
rect 50380 43002 50436 43004
rect 50460 43002 50516 43004
rect 50540 43002 50596 43004
rect 50300 42950 50326 43002
rect 50326 42950 50356 43002
rect 50380 42950 50390 43002
rect 50390 42950 50436 43002
rect 50460 42950 50506 43002
rect 50506 42950 50516 43002
rect 50540 42950 50570 43002
rect 50570 42950 50596 43002
rect 50300 42948 50356 42950
rect 50380 42948 50436 42950
rect 50460 42948 50516 42950
rect 50540 42948 50596 42950
rect 50300 41914 50356 41916
rect 50380 41914 50436 41916
rect 50460 41914 50516 41916
rect 50540 41914 50596 41916
rect 50300 41862 50326 41914
rect 50326 41862 50356 41914
rect 50380 41862 50390 41914
rect 50390 41862 50436 41914
rect 50460 41862 50506 41914
rect 50506 41862 50516 41914
rect 50540 41862 50570 41914
rect 50570 41862 50596 41914
rect 50300 41860 50356 41862
rect 50380 41860 50436 41862
rect 50460 41860 50516 41862
rect 50540 41860 50596 41862
rect 50300 40826 50356 40828
rect 50380 40826 50436 40828
rect 50460 40826 50516 40828
rect 50540 40826 50596 40828
rect 50300 40774 50326 40826
rect 50326 40774 50356 40826
rect 50380 40774 50390 40826
rect 50390 40774 50436 40826
rect 50460 40774 50506 40826
rect 50506 40774 50516 40826
rect 50540 40774 50570 40826
rect 50570 40774 50596 40826
rect 50300 40772 50356 40774
rect 50380 40772 50436 40774
rect 50460 40772 50516 40774
rect 50540 40772 50596 40774
rect 50300 39738 50356 39740
rect 50380 39738 50436 39740
rect 50460 39738 50516 39740
rect 50540 39738 50596 39740
rect 50300 39686 50326 39738
rect 50326 39686 50356 39738
rect 50380 39686 50390 39738
rect 50390 39686 50436 39738
rect 50460 39686 50506 39738
rect 50506 39686 50516 39738
rect 50540 39686 50570 39738
rect 50570 39686 50596 39738
rect 50300 39684 50356 39686
rect 50380 39684 50436 39686
rect 50460 39684 50516 39686
rect 50540 39684 50596 39686
rect 50300 38650 50356 38652
rect 50380 38650 50436 38652
rect 50460 38650 50516 38652
rect 50540 38650 50596 38652
rect 50300 38598 50326 38650
rect 50326 38598 50356 38650
rect 50380 38598 50390 38650
rect 50390 38598 50436 38650
rect 50460 38598 50506 38650
rect 50506 38598 50516 38650
rect 50540 38598 50570 38650
rect 50570 38598 50596 38650
rect 50300 38596 50356 38598
rect 50380 38596 50436 38598
rect 50460 38596 50516 38598
rect 50540 38596 50596 38598
rect 50300 37562 50356 37564
rect 50380 37562 50436 37564
rect 50460 37562 50516 37564
rect 50540 37562 50596 37564
rect 50300 37510 50326 37562
rect 50326 37510 50356 37562
rect 50380 37510 50390 37562
rect 50390 37510 50436 37562
rect 50460 37510 50506 37562
rect 50506 37510 50516 37562
rect 50540 37510 50570 37562
rect 50570 37510 50596 37562
rect 50300 37508 50356 37510
rect 50380 37508 50436 37510
rect 50460 37508 50516 37510
rect 50540 37508 50596 37510
rect 50300 36474 50356 36476
rect 50380 36474 50436 36476
rect 50460 36474 50516 36476
rect 50540 36474 50596 36476
rect 50300 36422 50326 36474
rect 50326 36422 50356 36474
rect 50380 36422 50390 36474
rect 50390 36422 50436 36474
rect 50460 36422 50506 36474
rect 50506 36422 50516 36474
rect 50540 36422 50570 36474
rect 50570 36422 50596 36474
rect 50300 36420 50356 36422
rect 50380 36420 50436 36422
rect 50460 36420 50516 36422
rect 50540 36420 50596 36422
rect 50300 35386 50356 35388
rect 50380 35386 50436 35388
rect 50460 35386 50516 35388
rect 50540 35386 50596 35388
rect 50300 35334 50326 35386
rect 50326 35334 50356 35386
rect 50380 35334 50390 35386
rect 50390 35334 50436 35386
rect 50460 35334 50506 35386
rect 50506 35334 50516 35386
rect 50540 35334 50570 35386
rect 50570 35334 50596 35386
rect 50300 35332 50356 35334
rect 50380 35332 50436 35334
rect 50460 35332 50516 35334
rect 50540 35332 50596 35334
rect 50300 34298 50356 34300
rect 50380 34298 50436 34300
rect 50460 34298 50516 34300
rect 50540 34298 50596 34300
rect 50300 34246 50326 34298
rect 50326 34246 50356 34298
rect 50380 34246 50390 34298
rect 50390 34246 50436 34298
rect 50460 34246 50506 34298
rect 50506 34246 50516 34298
rect 50540 34246 50570 34298
rect 50570 34246 50596 34298
rect 50300 34244 50356 34246
rect 50380 34244 50436 34246
rect 50460 34244 50516 34246
rect 50540 34244 50596 34246
rect 50300 33210 50356 33212
rect 50380 33210 50436 33212
rect 50460 33210 50516 33212
rect 50540 33210 50596 33212
rect 50300 33158 50326 33210
rect 50326 33158 50356 33210
rect 50380 33158 50390 33210
rect 50390 33158 50436 33210
rect 50460 33158 50506 33210
rect 50506 33158 50516 33210
rect 50540 33158 50570 33210
rect 50570 33158 50596 33210
rect 50300 33156 50356 33158
rect 50380 33156 50436 33158
rect 50460 33156 50516 33158
rect 50540 33156 50596 33158
rect 50300 32122 50356 32124
rect 50380 32122 50436 32124
rect 50460 32122 50516 32124
rect 50540 32122 50596 32124
rect 50300 32070 50326 32122
rect 50326 32070 50356 32122
rect 50380 32070 50390 32122
rect 50390 32070 50436 32122
rect 50460 32070 50506 32122
rect 50506 32070 50516 32122
rect 50540 32070 50570 32122
rect 50570 32070 50596 32122
rect 50300 32068 50356 32070
rect 50380 32068 50436 32070
rect 50460 32068 50516 32070
rect 50540 32068 50596 32070
rect 50300 31034 50356 31036
rect 50380 31034 50436 31036
rect 50460 31034 50516 31036
rect 50540 31034 50596 31036
rect 50300 30982 50326 31034
rect 50326 30982 50356 31034
rect 50380 30982 50390 31034
rect 50390 30982 50436 31034
rect 50460 30982 50506 31034
rect 50506 30982 50516 31034
rect 50540 30982 50570 31034
rect 50570 30982 50596 31034
rect 50300 30980 50356 30982
rect 50380 30980 50436 30982
rect 50460 30980 50516 30982
rect 50540 30980 50596 30982
rect 50300 29946 50356 29948
rect 50380 29946 50436 29948
rect 50460 29946 50516 29948
rect 50540 29946 50596 29948
rect 50300 29894 50326 29946
rect 50326 29894 50356 29946
rect 50380 29894 50390 29946
rect 50390 29894 50436 29946
rect 50460 29894 50506 29946
rect 50506 29894 50516 29946
rect 50540 29894 50570 29946
rect 50570 29894 50596 29946
rect 50300 29892 50356 29894
rect 50380 29892 50436 29894
rect 50460 29892 50516 29894
rect 50540 29892 50596 29894
rect 50300 28858 50356 28860
rect 50380 28858 50436 28860
rect 50460 28858 50516 28860
rect 50540 28858 50596 28860
rect 50300 28806 50326 28858
rect 50326 28806 50356 28858
rect 50380 28806 50390 28858
rect 50390 28806 50436 28858
rect 50460 28806 50506 28858
rect 50506 28806 50516 28858
rect 50540 28806 50570 28858
rect 50570 28806 50596 28858
rect 50300 28804 50356 28806
rect 50380 28804 50436 28806
rect 50460 28804 50516 28806
rect 50540 28804 50596 28806
rect 50300 27770 50356 27772
rect 50380 27770 50436 27772
rect 50460 27770 50516 27772
rect 50540 27770 50596 27772
rect 50300 27718 50326 27770
rect 50326 27718 50356 27770
rect 50380 27718 50390 27770
rect 50390 27718 50436 27770
rect 50460 27718 50506 27770
rect 50506 27718 50516 27770
rect 50540 27718 50570 27770
rect 50570 27718 50596 27770
rect 50300 27716 50356 27718
rect 50380 27716 50436 27718
rect 50460 27716 50516 27718
rect 50540 27716 50596 27718
rect 50300 26682 50356 26684
rect 50380 26682 50436 26684
rect 50460 26682 50516 26684
rect 50540 26682 50596 26684
rect 50300 26630 50326 26682
rect 50326 26630 50356 26682
rect 50380 26630 50390 26682
rect 50390 26630 50436 26682
rect 50460 26630 50506 26682
rect 50506 26630 50516 26682
rect 50540 26630 50570 26682
rect 50570 26630 50596 26682
rect 50300 26628 50356 26630
rect 50380 26628 50436 26630
rect 50460 26628 50516 26630
rect 50540 26628 50596 26630
rect 50300 25594 50356 25596
rect 50380 25594 50436 25596
rect 50460 25594 50516 25596
rect 50540 25594 50596 25596
rect 50300 25542 50326 25594
rect 50326 25542 50356 25594
rect 50380 25542 50390 25594
rect 50390 25542 50436 25594
rect 50460 25542 50506 25594
rect 50506 25542 50516 25594
rect 50540 25542 50570 25594
rect 50570 25542 50596 25594
rect 50300 25540 50356 25542
rect 50380 25540 50436 25542
rect 50460 25540 50516 25542
rect 50540 25540 50596 25542
rect 50300 24506 50356 24508
rect 50380 24506 50436 24508
rect 50460 24506 50516 24508
rect 50540 24506 50596 24508
rect 50300 24454 50326 24506
rect 50326 24454 50356 24506
rect 50380 24454 50390 24506
rect 50390 24454 50436 24506
rect 50460 24454 50506 24506
rect 50506 24454 50516 24506
rect 50540 24454 50570 24506
rect 50570 24454 50596 24506
rect 50300 24452 50356 24454
rect 50380 24452 50436 24454
rect 50460 24452 50516 24454
rect 50540 24452 50596 24454
rect 50300 23418 50356 23420
rect 50380 23418 50436 23420
rect 50460 23418 50516 23420
rect 50540 23418 50596 23420
rect 50300 23366 50326 23418
rect 50326 23366 50356 23418
rect 50380 23366 50390 23418
rect 50390 23366 50436 23418
rect 50460 23366 50506 23418
rect 50506 23366 50516 23418
rect 50540 23366 50570 23418
rect 50570 23366 50596 23418
rect 50300 23364 50356 23366
rect 50380 23364 50436 23366
rect 50460 23364 50516 23366
rect 50540 23364 50596 23366
rect 50300 22330 50356 22332
rect 50380 22330 50436 22332
rect 50460 22330 50516 22332
rect 50540 22330 50596 22332
rect 50300 22278 50326 22330
rect 50326 22278 50356 22330
rect 50380 22278 50390 22330
rect 50390 22278 50436 22330
rect 50460 22278 50506 22330
rect 50506 22278 50516 22330
rect 50540 22278 50570 22330
rect 50570 22278 50596 22330
rect 50300 22276 50356 22278
rect 50380 22276 50436 22278
rect 50460 22276 50516 22278
rect 50540 22276 50596 22278
rect 34940 14170 34996 14172
rect 35020 14170 35076 14172
rect 35100 14170 35156 14172
rect 35180 14170 35236 14172
rect 34940 14118 34966 14170
rect 34966 14118 34996 14170
rect 35020 14118 35030 14170
rect 35030 14118 35076 14170
rect 35100 14118 35146 14170
rect 35146 14118 35156 14170
rect 35180 14118 35210 14170
rect 35210 14118 35236 14170
rect 34940 14116 34996 14118
rect 35020 14116 35076 14118
rect 35100 14116 35156 14118
rect 35180 14116 35236 14118
rect 34940 13082 34996 13084
rect 35020 13082 35076 13084
rect 35100 13082 35156 13084
rect 35180 13082 35236 13084
rect 34940 13030 34966 13082
rect 34966 13030 34996 13082
rect 35020 13030 35030 13082
rect 35030 13030 35076 13082
rect 35100 13030 35146 13082
rect 35146 13030 35156 13082
rect 35180 13030 35210 13082
rect 35210 13030 35236 13082
rect 34940 13028 34996 13030
rect 35020 13028 35076 13030
rect 35100 13028 35156 13030
rect 35180 13028 35236 13030
rect 34940 11994 34996 11996
rect 35020 11994 35076 11996
rect 35100 11994 35156 11996
rect 35180 11994 35236 11996
rect 34940 11942 34966 11994
rect 34966 11942 34996 11994
rect 35020 11942 35030 11994
rect 35030 11942 35076 11994
rect 35100 11942 35146 11994
rect 35146 11942 35156 11994
rect 35180 11942 35210 11994
rect 35210 11942 35236 11994
rect 34940 11940 34996 11942
rect 35020 11940 35076 11942
rect 35100 11940 35156 11942
rect 35180 11940 35236 11942
rect 34940 10906 34996 10908
rect 35020 10906 35076 10908
rect 35100 10906 35156 10908
rect 35180 10906 35236 10908
rect 34940 10854 34966 10906
rect 34966 10854 34996 10906
rect 35020 10854 35030 10906
rect 35030 10854 35076 10906
rect 35100 10854 35146 10906
rect 35146 10854 35156 10906
rect 35180 10854 35210 10906
rect 35210 10854 35236 10906
rect 34940 10852 34996 10854
rect 35020 10852 35076 10854
rect 35100 10852 35156 10854
rect 35180 10852 35236 10854
rect 33966 7656 34022 7712
rect 33782 6024 33838 6080
rect 34242 7248 34298 7304
rect 34150 7148 34152 7168
rect 34152 7148 34204 7168
rect 34204 7148 34206 7168
rect 34150 7112 34206 7148
rect 34940 9818 34996 9820
rect 35020 9818 35076 9820
rect 35100 9818 35156 9820
rect 35180 9818 35236 9820
rect 34940 9766 34966 9818
rect 34966 9766 34996 9818
rect 35020 9766 35030 9818
rect 35030 9766 35076 9818
rect 35100 9766 35146 9818
rect 35146 9766 35156 9818
rect 35180 9766 35210 9818
rect 35210 9766 35236 9818
rect 34940 9764 34996 9766
rect 35020 9764 35076 9766
rect 35100 9764 35156 9766
rect 35180 9764 35236 9766
rect 34940 8730 34996 8732
rect 35020 8730 35076 8732
rect 35100 8730 35156 8732
rect 35180 8730 35236 8732
rect 34940 8678 34966 8730
rect 34966 8678 34996 8730
rect 35020 8678 35030 8730
rect 35030 8678 35076 8730
rect 35100 8678 35146 8730
rect 35146 8678 35156 8730
rect 35180 8678 35210 8730
rect 35210 8678 35236 8730
rect 34940 8676 34996 8678
rect 35020 8676 35076 8678
rect 35100 8676 35156 8678
rect 35180 8676 35236 8678
rect 34940 7642 34996 7644
rect 35020 7642 35076 7644
rect 35100 7642 35156 7644
rect 35180 7642 35236 7644
rect 34940 7590 34966 7642
rect 34966 7590 34996 7642
rect 35020 7590 35030 7642
rect 35030 7590 35076 7642
rect 35100 7590 35146 7642
rect 35146 7590 35156 7642
rect 35180 7590 35210 7642
rect 35210 7590 35236 7642
rect 34940 7588 34996 7590
rect 35020 7588 35076 7590
rect 35100 7588 35156 7590
rect 35180 7588 35236 7590
rect 34794 7112 34850 7168
rect 35254 7284 35256 7304
rect 35256 7284 35308 7304
rect 35308 7284 35310 7304
rect 35254 7248 35310 7284
rect 34940 6554 34996 6556
rect 35020 6554 35076 6556
rect 35100 6554 35156 6556
rect 35180 6554 35236 6556
rect 34940 6502 34966 6554
rect 34966 6502 34996 6554
rect 35020 6502 35030 6554
rect 35030 6502 35076 6554
rect 35100 6502 35146 6554
rect 35146 6502 35156 6554
rect 35180 6502 35210 6554
rect 35210 6502 35236 6554
rect 34940 6500 34996 6502
rect 35020 6500 35076 6502
rect 35100 6500 35156 6502
rect 35180 6500 35236 6502
rect 35254 5616 35310 5672
rect 34940 5466 34996 5468
rect 35020 5466 35076 5468
rect 35100 5466 35156 5468
rect 35180 5466 35236 5468
rect 34940 5414 34966 5466
rect 34966 5414 34996 5466
rect 35020 5414 35030 5466
rect 35030 5414 35076 5466
rect 35100 5414 35146 5466
rect 35146 5414 35156 5466
rect 35180 5414 35210 5466
rect 35210 5414 35236 5466
rect 34940 5412 34996 5414
rect 35020 5412 35076 5414
rect 35100 5412 35156 5414
rect 35180 5412 35236 5414
rect 34518 5092 34574 5128
rect 34518 5072 34520 5092
rect 34520 5072 34572 5092
rect 34572 5072 34574 5092
rect 34940 4378 34996 4380
rect 35020 4378 35076 4380
rect 35100 4378 35156 4380
rect 35180 4378 35236 4380
rect 34940 4326 34966 4378
rect 34966 4326 34996 4378
rect 35020 4326 35030 4378
rect 35030 4326 35076 4378
rect 35100 4326 35146 4378
rect 35146 4326 35156 4378
rect 35180 4326 35210 4378
rect 35210 4326 35236 4378
rect 34940 4324 34996 4326
rect 35020 4324 35076 4326
rect 35100 4324 35156 4326
rect 35180 4324 35236 4326
rect 35898 6976 35954 7032
rect 36174 7384 36230 7440
rect 36082 6840 36138 6896
rect 34940 3290 34996 3292
rect 35020 3290 35076 3292
rect 35100 3290 35156 3292
rect 35180 3290 35236 3292
rect 34940 3238 34966 3290
rect 34966 3238 34996 3290
rect 35020 3238 35030 3290
rect 35030 3238 35076 3290
rect 35100 3238 35146 3290
rect 35146 3238 35156 3290
rect 35180 3238 35210 3290
rect 35210 3238 35236 3290
rect 34940 3236 34996 3238
rect 35020 3236 35076 3238
rect 35100 3236 35156 3238
rect 35180 3236 35236 3238
rect 34940 2202 34996 2204
rect 35020 2202 35076 2204
rect 35100 2202 35156 2204
rect 35180 2202 35236 2204
rect 34940 2150 34966 2202
rect 34966 2150 34996 2202
rect 35020 2150 35030 2202
rect 35030 2150 35076 2202
rect 35100 2150 35146 2202
rect 35146 2150 35156 2202
rect 35180 2150 35210 2202
rect 35210 2150 35236 2202
rect 34940 2148 34996 2150
rect 35020 2148 35076 2150
rect 35100 2148 35156 2150
rect 35180 2148 35236 2150
rect 36174 6160 36230 6216
rect 36634 6860 36690 6896
rect 36634 6840 36636 6860
rect 36636 6840 36688 6860
rect 36688 6840 36690 6860
rect 36082 4120 36138 4176
rect 37186 6160 37242 6216
rect 37278 4820 37334 4856
rect 37278 4800 37280 4820
rect 37280 4800 37332 4820
rect 37332 4800 37334 4820
rect 37646 6860 37702 6896
rect 37646 6840 37648 6860
rect 37648 6840 37700 6860
rect 37700 6840 37702 6860
rect 38290 6160 38346 6216
rect 37738 5752 37794 5808
rect 38106 5616 38162 5672
rect 39118 8200 39174 8256
rect 38658 8064 38714 8120
rect 39210 7928 39266 7984
rect 39486 7520 39542 7576
rect 39394 7384 39450 7440
rect 39486 5772 39542 5808
rect 39486 5752 39488 5772
rect 39488 5752 39540 5772
rect 39540 5752 39542 5772
rect 39946 8064 40002 8120
rect 40038 7112 40094 7168
rect 39946 6976 40002 7032
rect 39854 4120 39910 4176
rect 41050 7792 41106 7848
rect 40866 6740 40868 6760
rect 40868 6740 40920 6760
rect 40920 6740 40922 6760
rect 40866 6704 40922 6740
rect 41234 8064 41290 8120
rect 41602 8064 41658 8120
rect 41510 7520 41566 7576
rect 41878 7656 41934 7712
rect 41694 7284 41696 7304
rect 41696 7284 41748 7304
rect 41748 7284 41750 7304
rect 41694 7248 41750 7284
rect 41694 6976 41750 7032
rect 41142 6840 41198 6896
rect 41142 6160 41198 6216
rect 41878 6860 41934 6896
rect 41878 6840 41880 6860
rect 41880 6840 41932 6860
rect 41932 6840 41934 6860
rect 42338 7384 42394 7440
rect 50300 21242 50356 21244
rect 50380 21242 50436 21244
rect 50460 21242 50516 21244
rect 50540 21242 50596 21244
rect 50300 21190 50326 21242
rect 50326 21190 50356 21242
rect 50380 21190 50390 21242
rect 50390 21190 50436 21242
rect 50460 21190 50506 21242
rect 50506 21190 50516 21242
rect 50540 21190 50570 21242
rect 50570 21190 50596 21242
rect 50300 21188 50356 21190
rect 50380 21188 50436 21190
rect 50460 21188 50516 21190
rect 50540 21188 50596 21190
rect 50300 20154 50356 20156
rect 50380 20154 50436 20156
rect 50460 20154 50516 20156
rect 50540 20154 50596 20156
rect 50300 20102 50326 20154
rect 50326 20102 50356 20154
rect 50380 20102 50390 20154
rect 50390 20102 50436 20154
rect 50460 20102 50506 20154
rect 50506 20102 50516 20154
rect 50540 20102 50570 20154
rect 50570 20102 50596 20154
rect 50300 20100 50356 20102
rect 50380 20100 50436 20102
rect 50460 20100 50516 20102
rect 50540 20100 50596 20102
rect 50300 19066 50356 19068
rect 50380 19066 50436 19068
rect 50460 19066 50516 19068
rect 50540 19066 50596 19068
rect 50300 19014 50326 19066
rect 50326 19014 50356 19066
rect 50380 19014 50390 19066
rect 50390 19014 50436 19066
rect 50460 19014 50506 19066
rect 50506 19014 50516 19066
rect 50540 19014 50570 19066
rect 50570 19014 50596 19066
rect 50300 19012 50356 19014
rect 50380 19012 50436 19014
rect 50460 19012 50516 19014
rect 50540 19012 50596 19014
rect 42798 7792 42854 7848
rect 42614 7384 42670 7440
rect 44178 7948 44234 7984
rect 44178 7928 44180 7948
rect 44180 7928 44232 7948
rect 44232 7928 44234 7948
rect 43626 7284 43628 7304
rect 43628 7284 43680 7304
rect 43680 7284 43682 7304
rect 43626 7248 43682 7284
rect 44086 6724 44142 6760
rect 44086 6704 44088 6724
rect 44088 6704 44140 6724
rect 44140 6704 44142 6724
rect 43810 5772 43866 5808
rect 43810 5752 43812 5772
rect 43812 5752 43864 5772
rect 43864 5752 43866 5772
rect 43718 5208 43774 5264
rect 44638 6976 44694 7032
rect 44270 6160 44326 6216
rect 45006 6976 45062 7032
rect 45558 6160 45614 6216
rect 46018 8200 46074 8256
rect 46018 7928 46074 7984
rect 50300 17978 50356 17980
rect 50380 17978 50436 17980
rect 50460 17978 50516 17980
rect 50540 17978 50596 17980
rect 50300 17926 50326 17978
rect 50326 17926 50356 17978
rect 50380 17926 50390 17978
rect 50390 17926 50436 17978
rect 50460 17926 50506 17978
rect 50506 17926 50516 17978
rect 50540 17926 50570 17978
rect 50570 17926 50596 17978
rect 50300 17924 50356 17926
rect 50380 17924 50436 17926
rect 50460 17924 50516 17926
rect 50540 17924 50596 17926
rect 46386 8200 46442 8256
rect 46294 7792 46350 7848
rect 46478 6452 46534 6488
rect 46478 6432 46480 6452
rect 46480 6432 46532 6452
rect 46532 6432 46534 6452
rect 46018 5888 46074 5944
rect 46018 5480 46074 5536
rect 46662 6860 46718 6896
rect 46938 7656 46994 7712
rect 46938 7384 46994 7440
rect 46662 6840 46664 6860
rect 46664 6840 46716 6860
rect 46716 6840 46718 6860
rect 47306 8200 47362 8256
rect 47398 8064 47454 8120
rect 47214 7520 47270 7576
rect 46846 6568 46902 6624
rect 46938 6432 46994 6488
rect 46846 6024 46902 6080
rect 46662 5652 46664 5672
rect 46664 5652 46716 5672
rect 46716 5652 46718 5672
rect 46662 5616 46718 5652
rect 47214 6704 47270 6760
rect 47398 6840 47454 6896
rect 47490 6432 47546 6488
rect 47674 6976 47730 7032
rect 47582 6024 47638 6080
rect 47490 5908 47546 5944
rect 47490 5888 47492 5908
rect 47492 5888 47544 5908
rect 47544 5888 47546 5908
rect 47490 5636 47546 5672
rect 47490 5616 47492 5636
rect 47492 5616 47544 5636
rect 47544 5616 47546 5636
rect 47398 5208 47454 5264
rect 47950 7964 47952 7984
rect 47952 7964 48004 7984
rect 48004 7964 48006 7984
rect 47950 7928 48006 7964
rect 47858 6568 47914 6624
rect 47858 6180 47914 6216
rect 47858 6160 47860 6180
rect 47860 6160 47912 6180
rect 47912 6160 47914 6180
rect 47858 5516 47860 5536
rect 47860 5516 47912 5536
rect 47912 5516 47914 5536
rect 47858 5480 47914 5516
rect 48502 7964 48504 7984
rect 48504 7964 48556 7984
rect 48556 7964 48558 7984
rect 48502 7928 48558 7964
rect 50300 16890 50356 16892
rect 50380 16890 50436 16892
rect 50460 16890 50516 16892
rect 50540 16890 50596 16892
rect 50300 16838 50326 16890
rect 50326 16838 50356 16890
rect 50380 16838 50390 16890
rect 50390 16838 50436 16890
rect 50460 16838 50506 16890
rect 50506 16838 50516 16890
rect 50540 16838 50570 16890
rect 50570 16838 50596 16890
rect 50300 16836 50356 16838
rect 50380 16836 50436 16838
rect 50460 16836 50516 16838
rect 50540 16836 50596 16838
rect 50300 15802 50356 15804
rect 50380 15802 50436 15804
rect 50460 15802 50516 15804
rect 50540 15802 50596 15804
rect 50300 15750 50326 15802
rect 50326 15750 50356 15802
rect 50380 15750 50390 15802
rect 50390 15750 50436 15802
rect 50460 15750 50506 15802
rect 50506 15750 50516 15802
rect 50540 15750 50570 15802
rect 50570 15750 50596 15802
rect 50300 15748 50356 15750
rect 50380 15748 50436 15750
rect 50460 15748 50516 15750
rect 50540 15748 50596 15750
rect 50300 14714 50356 14716
rect 50380 14714 50436 14716
rect 50460 14714 50516 14716
rect 50540 14714 50596 14716
rect 50300 14662 50326 14714
rect 50326 14662 50356 14714
rect 50380 14662 50390 14714
rect 50390 14662 50436 14714
rect 50460 14662 50506 14714
rect 50506 14662 50516 14714
rect 50540 14662 50570 14714
rect 50570 14662 50596 14714
rect 50300 14660 50356 14662
rect 50380 14660 50436 14662
rect 50460 14660 50516 14662
rect 50540 14660 50596 14662
rect 50300 13626 50356 13628
rect 50380 13626 50436 13628
rect 50460 13626 50516 13628
rect 50540 13626 50596 13628
rect 50300 13574 50326 13626
rect 50326 13574 50356 13626
rect 50380 13574 50390 13626
rect 50390 13574 50436 13626
rect 50460 13574 50506 13626
rect 50506 13574 50516 13626
rect 50540 13574 50570 13626
rect 50570 13574 50596 13626
rect 50300 13572 50356 13574
rect 50380 13572 50436 13574
rect 50460 13572 50516 13574
rect 50540 13572 50596 13574
rect 50300 12538 50356 12540
rect 50380 12538 50436 12540
rect 50460 12538 50516 12540
rect 50540 12538 50596 12540
rect 50300 12486 50326 12538
rect 50326 12486 50356 12538
rect 50380 12486 50390 12538
rect 50390 12486 50436 12538
rect 50460 12486 50506 12538
rect 50506 12486 50516 12538
rect 50540 12486 50570 12538
rect 50570 12486 50596 12538
rect 50300 12484 50356 12486
rect 50380 12484 50436 12486
rect 50460 12484 50516 12486
rect 50540 12484 50596 12486
rect 50300 11450 50356 11452
rect 50380 11450 50436 11452
rect 50460 11450 50516 11452
rect 50540 11450 50596 11452
rect 50300 11398 50326 11450
rect 50326 11398 50356 11450
rect 50380 11398 50390 11450
rect 50390 11398 50436 11450
rect 50460 11398 50506 11450
rect 50506 11398 50516 11450
rect 50540 11398 50570 11450
rect 50570 11398 50596 11450
rect 50300 11396 50356 11398
rect 50380 11396 50436 11398
rect 50460 11396 50516 11398
rect 50540 11396 50596 11398
rect 50300 10362 50356 10364
rect 50380 10362 50436 10364
rect 50460 10362 50516 10364
rect 50540 10362 50596 10364
rect 50300 10310 50326 10362
rect 50326 10310 50356 10362
rect 50380 10310 50390 10362
rect 50390 10310 50436 10362
rect 50460 10310 50506 10362
rect 50506 10310 50516 10362
rect 50540 10310 50570 10362
rect 50570 10310 50596 10362
rect 50300 10308 50356 10310
rect 50380 10308 50436 10310
rect 50460 10308 50516 10310
rect 50540 10308 50596 10310
rect 48686 7792 48742 7848
rect 49330 7520 49386 7576
rect 49238 7420 49240 7440
rect 49240 7420 49292 7440
rect 49292 7420 49294 7440
rect 49238 7384 49294 7420
rect 49146 7112 49202 7168
rect 48962 6568 49018 6624
rect 48686 6024 48742 6080
rect 48962 6180 49018 6216
rect 48962 6160 48964 6180
rect 48964 6160 49016 6180
rect 49016 6160 49018 6180
rect 48778 5752 48834 5808
rect 50300 9274 50356 9276
rect 50380 9274 50436 9276
rect 50460 9274 50516 9276
rect 50540 9274 50596 9276
rect 50300 9222 50326 9274
rect 50326 9222 50356 9274
rect 50380 9222 50390 9274
rect 50390 9222 50436 9274
rect 50460 9222 50506 9274
rect 50506 9222 50516 9274
rect 50540 9222 50570 9274
rect 50570 9222 50596 9274
rect 50300 9220 50356 9222
rect 50380 9220 50436 9222
rect 50460 9220 50516 9222
rect 50540 9220 50596 9222
rect 50300 8186 50356 8188
rect 50380 8186 50436 8188
rect 50460 8186 50516 8188
rect 50540 8186 50596 8188
rect 50300 8134 50326 8186
rect 50326 8134 50356 8186
rect 50380 8134 50390 8186
rect 50390 8134 50436 8186
rect 50460 8134 50506 8186
rect 50506 8134 50516 8186
rect 50540 8134 50570 8186
rect 50570 8134 50596 8186
rect 50300 8132 50356 8134
rect 50380 8132 50436 8134
rect 50460 8132 50516 8134
rect 50540 8132 50596 8134
rect 50894 7384 50950 7440
rect 51078 7384 51134 7440
rect 50158 7112 50214 7168
rect 49790 6432 49846 6488
rect 50300 7098 50356 7100
rect 50380 7098 50436 7100
rect 50460 7098 50516 7100
rect 50540 7098 50596 7100
rect 50300 7046 50326 7098
rect 50326 7046 50356 7098
rect 50380 7046 50390 7098
rect 50390 7046 50436 7098
rect 50460 7046 50506 7098
rect 50506 7046 50516 7098
rect 50540 7046 50570 7098
rect 50570 7046 50596 7098
rect 50300 7044 50356 7046
rect 50380 7044 50436 7046
rect 50460 7044 50516 7046
rect 50540 7044 50596 7046
rect 50066 6432 50122 6488
rect 50066 6024 50122 6080
rect 50300 6010 50356 6012
rect 50380 6010 50436 6012
rect 50460 6010 50516 6012
rect 50540 6010 50596 6012
rect 50300 5958 50326 6010
rect 50326 5958 50356 6010
rect 50380 5958 50390 6010
rect 50390 5958 50436 6010
rect 50460 5958 50506 6010
rect 50506 5958 50516 6010
rect 50540 5958 50570 6010
rect 50570 5958 50596 6010
rect 50300 5956 50356 5958
rect 50380 5956 50436 5958
rect 50460 5956 50516 5958
rect 50540 5956 50596 5958
rect 50300 4922 50356 4924
rect 50380 4922 50436 4924
rect 50460 4922 50516 4924
rect 50540 4922 50596 4924
rect 50300 4870 50326 4922
rect 50326 4870 50356 4922
rect 50380 4870 50390 4922
rect 50390 4870 50436 4922
rect 50460 4870 50506 4922
rect 50506 4870 50516 4922
rect 50540 4870 50570 4922
rect 50570 4870 50596 4922
rect 50300 4868 50356 4870
rect 50380 4868 50436 4870
rect 50460 4868 50516 4870
rect 50540 4868 50596 4870
rect 50300 3834 50356 3836
rect 50380 3834 50436 3836
rect 50460 3834 50516 3836
rect 50540 3834 50596 3836
rect 50300 3782 50326 3834
rect 50326 3782 50356 3834
rect 50380 3782 50390 3834
rect 50390 3782 50436 3834
rect 50460 3782 50506 3834
rect 50506 3782 50516 3834
rect 50540 3782 50570 3834
rect 50570 3782 50596 3834
rect 50300 3780 50356 3782
rect 50380 3780 50436 3782
rect 50460 3780 50516 3782
rect 50540 3780 50596 3782
rect 50300 2746 50356 2748
rect 50380 2746 50436 2748
rect 50460 2746 50516 2748
rect 50540 2746 50596 2748
rect 50300 2694 50326 2746
rect 50326 2694 50356 2746
rect 50380 2694 50390 2746
rect 50390 2694 50436 2746
rect 50460 2694 50506 2746
rect 50506 2694 50516 2746
rect 50540 2694 50570 2746
rect 50570 2694 50596 2746
rect 50300 2692 50356 2694
rect 50380 2692 50436 2694
rect 50460 2692 50516 2694
rect 50540 2692 50596 2694
rect 53194 5772 53250 5808
rect 53194 5752 53196 5772
rect 53196 5752 53248 5772
rect 53248 5752 53250 5772
rect 54206 6432 54262 6488
rect 54298 5772 54354 5808
rect 54298 5752 54300 5772
rect 54300 5752 54352 5772
rect 54352 5752 54354 5772
rect 55862 7928 55918 7984
rect 57886 6568 57942 6624
rect 58070 6704 58126 6760
rect 58346 6432 58402 6488
rect 59174 6704 59230 6760
rect 58714 6296 58770 6352
rect 65660 116442 65716 116444
rect 65740 116442 65796 116444
rect 65820 116442 65876 116444
rect 65900 116442 65956 116444
rect 65660 116390 65686 116442
rect 65686 116390 65716 116442
rect 65740 116390 65750 116442
rect 65750 116390 65796 116442
rect 65820 116390 65866 116442
rect 65866 116390 65876 116442
rect 65900 116390 65930 116442
rect 65930 116390 65956 116442
rect 65660 116388 65716 116390
rect 65740 116388 65796 116390
rect 65820 116388 65876 116390
rect 65900 116388 65956 116390
rect 65660 115354 65716 115356
rect 65740 115354 65796 115356
rect 65820 115354 65876 115356
rect 65900 115354 65956 115356
rect 65660 115302 65686 115354
rect 65686 115302 65716 115354
rect 65740 115302 65750 115354
rect 65750 115302 65796 115354
rect 65820 115302 65866 115354
rect 65866 115302 65876 115354
rect 65900 115302 65930 115354
rect 65930 115302 65956 115354
rect 65660 115300 65716 115302
rect 65740 115300 65796 115302
rect 65820 115300 65876 115302
rect 65900 115300 65956 115302
rect 65660 114266 65716 114268
rect 65740 114266 65796 114268
rect 65820 114266 65876 114268
rect 65900 114266 65956 114268
rect 65660 114214 65686 114266
rect 65686 114214 65716 114266
rect 65740 114214 65750 114266
rect 65750 114214 65796 114266
rect 65820 114214 65866 114266
rect 65866 114214 65876 114266
rect 65900 114214 65930 114266
rect 65930 114214 65956 114266
rect 65660 114212 65716 114214
rect 65740 114212 65796 114214
rect 65820 114212 65876 114214
rect 65900 114212 65956 114214
rect 65660 113178 65716 113180
rect 65740 113178 65796 113180
rect 65820 113178 65876 113180
rect 65900 113178 65956 113180
rect 65660 113126 65686 113178
rect 65686 113126 65716 113178
rect 65740 113126 65750 113178
rect 65750 113126 65796 113178
rect 65820 113126 65866 113178
rect 65866 113126 65876 113178
rect 65900 113126 65930 113178
rect 65930 113126 65956 113178
rect 65660 113124 65716 113126
rect 65740 113124 65796 113126
rect 65820 113124 65876 113126
rect 65900 113124 65956 113126
rect 65660 112090 65716 112092
rect 65740 112090 65796 112092
rect 65820 112090 65876 112092
rect 65900 112090 65956 112092
rect 65660 112038 65686 112090
rect 65686 112038 65716 112090
rect 65740 112038 65750 112090
rect 65750 112038 65796 112090
rect 65820 112038 65866 112090
rect 65866 112038 65876 112090
rect 65900 112038 65930 112090
rect 65930 112038 65956 112090
rect 65660 112036 65716 112038
rect 65740 112036 65796 112038
rect 65820 112036 65876 112038
rect 65900 112036 65956 112038
rect 65660 111002 65716 111004
rect 65740 111002 65796 111004
rect 65820 111002 65876 111004
rect 65900 111002 65956 111004
rect 65660 110950 65686 111002
rect 65686 110950 65716 111002
rect 65740 110950 65750 111002
rect 65750 110950 65796 111002
rect 65820 110950 65866 111002
rect 65866 110950 65876 111002
rect 65900 110950 65930 111002
rect 65930 110950 65956 111002
rect 65660 110948 65716 110950
rect 65740 110948 65796 110950
rect 65820 110948 65876 110950
rect 65900 110948 65956 110950
rect 65660 109914 65716 109916
rect 65740 109914 65796 109916
rect 65820 109914 65876 109916
rect 65900 109914 65956 109916
rect 65660 109862 65686 109914
rect 65686 109862 65716 109914
rect 65740 109862 65750 109914
rect 65750 109862 65796 109914
rect 65820 109862 65866 109914
rect 65866 109862 65876 109914
rect 65900 109862 65930 109914
rect 65930 109862 65956 109914
rect 65660 109860 65716 109862
rect 65740 109860 65796 109862
rect 65820 109860 65876 109862
rect 65900 109860 65956 109862
rect 65660 108826 65716 108828
rect 65740 108826 65796 108828
rect 65820 108826 65876 108828
rect 65900 108826 65956 108828
rect 65660 108774 65686 108826
rect 65686 108774 65716 108826
rect 65740 108774 65750 108826
rect 65750 108774 65796 108826
rect 65820 108774 65866 108826
rect 65866 108774 65876 108826
rect 65900 108774 65930 108826
rect 65930 108774 65956 108826
rect 65660 108772 65716 108774
rect 65740 108772 65796 108774
rect 65820 108772 65876 108774
rect 65900 108772 65956 108774
rect 65660 107738 65716 107740
rect 65740 107738 65796 107740
rect 65820 107738 65876 107740
rect 65900 107738 65956 107740
rect 65660 107686 65686 107738
rect 65686 107686 65716 107738
rect 65740 107686 65750 107738
rect 65750 107686 65796 107738
rect 65820 107686 65866 107738
rect 65866 107686 65876 107738
rect 65900 107686 65930 107738
rect 65930 107686 65956 107738
rect 65660 107684 65716 107686
rect 65740 107684 65796 107686
rect 65820 107684 65876 107686
rect 65900 107684 65956 107686
rect 65660 106650 65716 106652
rect 65740 106650 65796 106652
rect 65820 106650 65876 106652
rect 65900 106650 65956 106652
rect 65660 106598 65686 106650
rect 65686 106598 65716 106650
rect 65740 106598 65750 106650
rect 65750 106598 65796 106650
rect 65820 106598 65866 106650
rect 65866 106598 65876 106650
rect 65900 106598 65930 106650
rect 65930 106598 65956 106650
rect 65660 106596 65716 106598
rect 65740 106596 65796 106598
rect 65820 106596 65876 106598
rect 65900 106596 65956 106598
rect 65660 105562 65716 105564
rect 65740 105562 65796 105564
rect 65820 105562 65876 105564
rect 65900 105562 65956 105564
rect 65660 105510 65686 105562
rect 65686 105510 65716 105562
rect 65740 105510 65750 105562
rect 65750 105510 65796 105562
rect 65820 105510 65866 105562
rect 65866 105510 65876 105562
rect 65900 105510 65930 105562
rect 65930 105510 65956 105562
rect 65660 105508 65716 105510
rect 65740 105508 65796 105510
rect 65820 105508 65876 105510
rect 65900 105508 65956 105510
rect 65660 104474 65716 104476
rect 65740 104474 65796 104476
rect 65820 104474 65876 104476
rect 65900 104474 65956 104476
rect 65660 104422 65686 104474
rect 65686 104422 65716 104474
rect 65740 104422 65750 104474
rect 65750 104422 65796 104474
rect 65820 104422 65866 104474
rect 65866 104422 65876 104474
rect 65900 104422 65930 104474
rect 65930 104422 65956 104474
rect 65660 104420 65716 104422
rect 65740 104420 65796 104422
rect 65820 104420 65876 104422
rect 65900 104420 65956 104422
rect 65660 103386 65716 103388
rect 65740 103386 65796 103388
rect 65820 103386 65876 103388
rect 65900 103386 65956 103388
rect 65660 103334 65686 103386
rect 65686 103334 65716 103386
rect 65740 103334 65750 103386
rect 65750 103334 65796 103386
rect 65820 103334 65866 103386
rect 65866 103334 65876 103386
rect 65900 103334 65930 103386
rect 65930 103334 65956 103386
rect 65660 103332 65716 103334
rect 65740 103332 65796 103334
rect 65820 103332 65876 103334
rect 65900 103332 65956 103334
rect 65660 102298 65716 102300
rect 65740 102298 65796 102300
rect 65820 102298 65876 102300
rect 65900 102298 65956 102300
rect 65660 102246 65686 102298
rect 65686 102246 65716 102298
rect 65740 102246 65750 102298
rect 65750 102246 65796 102298
rect 65820 102246 65866 102298
rect 65866 102246 65876 102298
rect 65900 102246 65930 102298
rect 65930 102246 65956 102298
rect 65660 102244 65716 102246
rect 65740 102244 65796 102246
rect 65820 102244 65876 102246
rect 65900 102244 65956 102246
rect 65660 101210 65716 101212
rect 65740 101210 65796 101212
rect 65820 101210 65876 101212
rect 65900 101210 65956 101212
rect 65660 101158 65686 101210
rect 65686 101158 65716 101210
rect 65740 101158 65750 101210
rect 65750 101158 65796 101210
rect 65820 101158 65866 101210
rect 65866 101158 65876 101210
rect 65900 101158 65930 101210
rect 65930 101158 65956 101210
rect 65660 101156 65716 101158
rect 65740 101156 65796 101158
rect 65820 101156 65876 101158
rect 65900 101156 65956 101158
rect 65660 100122 65716 100124
rect 65740 100122 65796 100124
rect 65820 100122 65876 100124
rect 65900 100122 65956 100124
rect 65660 100070 65686 100122
rect 65686 100070 65716 100122
rect 65740 100070 65750 100122
rect 65750 100070 65796 100122
rect 65820 100070 65866 100122
rect 65866 100070 65876 100122
rect 65900 100070 65930 100122
rect 65930 100070 65956 100122
rect 65660 100068 65716 100070
rect 65740 100068 65796 100070
rect 65820 100068 65876 100070
rect 65900 100068 65956 100070
rect 65660 99034 65716 99036
rect 65740 99034 65796 99036
rect 65820 99034 65876 99036
rect 65900 99034 65956 99036
rect 65660 98982 65686 99034
rect 65686 98982 65716 99034
rect 65740 98982 65750 99034
rect 65750 98982 65796 99034
rect 65820 98982 65866 99034
rect 65866 98982 65876 99034
rect 65900 98982 65930 99034
rect 65930 98982 65956 99034
rect 65660 98980 65716 98982
rect 65740 98980 65796 98982
rect 65820 98980 65876 98982
rect 65900 98980 65956 98982
rect 65660 97946 65716 97948
rect 65740 97946 65796 97948
rect 65820 97946 65876 97948
rect 65900 97946 65956 97948
rect 65660 97894 65686 97946
rect 65686 97894 65716 97946
rect 65740 97894 65750 97946
rect 65750 97894 65796 97946
rect 65820 97894 65866 97946
rect 65866 97894 65876 97946
rect 65900 97894 65930 97946
rect 65930 97894 65956 97946
rect 65660 97892 65716 97894
rect 65740 97892 65796 97894
rect 65820 97892 65876 97894
rect 65900 97892 65956 97894
rect 65660 96858 65716 96860
rect 65740 96858 65796 96860
rect 65820 96858 65876 96860
rect 65900 96858 65956 96860
rect 65660 96806 65686 96858
rect 65686 96806 65716 96858
rect 65740 96806 65750 96858
rect 65750 96806 65796 96858
rect 65820 96806 65866 96858
rect 65866 96806 65876 96858
rect 65900 96806 65930 96858
rect 65930 96806 65956 96858
rect 65660 96804 65716 96806
rect 65740 96804 65796 96806
rect 65820 96804 65876 96806
rect 65900 96804 65956 96806
rect 65660 95770 65716 95772
rect 65740 95770 65796 95772
rect 65820 95770 65876 95772
rect 65900 95770 65956 95772
rect 65660 95718 65686 95770
rect 65686 95718 65716 95770
rect 65740 95718 65750 95770
rect 65750 95718 65796 95770
rect 65820 95718 65866 95770
rect 65866 95718 65876 95770
rect 65900 95718 65930 95770
rect 65930 95718 65956 95770
rect 65660 95716 65716 95718
rect 65740 95716 65796 95718
rect 65820 95716 65876 95718
rect 65900 95716 65956 95718
rect 65660 94682 65716 94684
rect 65740 94682 65796 94684
rect 65820 94682 65876 94684
rect 65900 94682 65956 94684
rect 65660 94630 65686 94682
rect 65686 94630 65716 94682
rect 65740 94630 65750 94682
rect 65750 94630 65796 94682
rect 65820 94630 65866 94682
rect 65866 94630 65876 94682
rect 65900 94630 65930 94682
rect 65930 94630 65956 94682
rect 65660 94628 65716 94630
rect 65740 94628 65796 94630
rect 65820 94628 65876 94630
rect 65900 94628 65956 94630
rect 65660 93594 65716 93596
rect 65740 93594 65796 93596
rect 65820 93594 65876 93596
rect 65900 93594 65956 93596
rect 65660 93542 65686 93594
rect 65686 93542 65716 93594
rect 65740 93542 65750 93594
rect 65750 93542 65796 93594
rect 65820 93542 65866 93594
rect 65866 93542 65876 93594
rect 65900 93542 65930 93594
rect 65930 93542 65956 93594
rect 65660 93540 65716 93542
rect 65740 93540 65796 93542
rect 65820 93540 65876 93542
rect 65900 93540 65956 93542
rect 65660 92506 65716 92508
rect 65740 92506 65796 92508
rect 65820 92506 65876 92508
rect 65900 92506 65956 92508
rect 65660 92454 65686 92506
rect 65686 92454 65716 92506
rect 65740 92454 65750 92506
rect 65750 92454 65796 92506
rect 65820 92454 65866 92506
rect 65866 92454 65876 92506
rect 65900 92454 65930 92506
rect 65930 92454 65956 92506
rect 65660 92452 65716 92454
rect 65740 92452 65796 92454
rect 65820 92452 65876 92454
rect 65900 92452 65956 92454
rect 65660 91418 65716 91420
rect 65740 91418 65796 91420
rect 65820 91418 65876 91420
rect 65900 91418 65956 91420
rect 65660 91366 65686 91418
rect 65686 91366 65716 91418
rect 65740 91366 65750 91418
rect 65750 91366 65796 91418
rect 65820 91366 65866 91418
rect 65866 91366 65876 91418
rect 65900 91366 65930 91418
rect 65930 91366 65956 91418
rect 65660 91364 65716 91366
rect 65740 91364 65796 91366
rect 65820 91364 65876 91366
rect 65900 91364 65956 91366
rect 65660 90330 65716 90332
rect 65740 90330 65796 90332
rect 65820 90330 65876 90332
rect 65900 90330 65956 90332
rect 65660 90278 65686 90330
rect 65686 90278 65716 90330
rect 65740 90278 65750 90330
rect 65750 90278 65796 90330
rect 65820 90278 65866 90330
rect 65866 90278 65876 90330
rect 65900 90278 65930 90330
rect 65930 90278 65956 90330
rect 65660 90276 65716 90278
rect 65740 90276 65796 90278
rect 65820 90276 65876 90278
rect 65900 90276 65956 90278
rect 65660 89242 65716 89244
rect 65740 89242 65796 89244
rect 65820 89242 65876 89244
rect 65900 89242 65956 89244
rect 65660 89190 65686 89242
rect 65686 89190 65716 89242
rect 65740 89190 65750 89242
rect 65750 89190 65796 89242
rect 65820 89190 65866 89242
rect 65866 89190 65876 89242
rect 65900 89190 65930 89242
rect 65930 89190 65956 89242
rect 65660 89188 65716 89190
rect 65740 89188 65796 89190
rect 65820 89188 65876 89190
rect 65900 89188 65956 89190
rect 65660 88154 65716 88156
rect 65740 88154 65796 88156
rect 65820 88154 65876 88156
rect 65900 88154 65956 88156
rect 65660 88102 65686 88154
rect 65686 88102 65716 88154
rect 65740 88102 65750 88154
rect 65750 88102 65796 88154
rect 65820 88102 65866 88154
rect 65866 88102 65876 88154
rect 65900 88102 65930 88154
rect 65930 88102 65956 88154
rect 65660 88100 65716 88102
rect 65740 88100 65796 88102
rect 65820 88100 65876 88102
rect 65900 88100 65956 88102
rect 65660 87066 65716 87068
rect 65740 87066 65796 87068
rect 65820 87066 65876 87068
rect 65900 87066 65956 87068
rect 65660 87014 65686 87066
rect 65686 87014 65716 87066
rect 65740 87014 65750 87066
rect 65750 87014 65796 87066
rect 65820 87014 65866 87066
rect 65866 87014 65876 87066
rect 65900 87014 65930 87066
rect 65930 87014 65956 87066
rect 65660 87012 65716 87014
rect 65740 87012 65796 87014
rect 65820 87012 65876 87014
rect 65900 87012 65956 87014
rect 65660 85978 65716 85980
rect 65740 85978 65796 85980
rect 65820 85978 65876 85980
rect 65900 85978 65956 85980
rect 65660 85926 65686 85978
rect 65686 85926 65716 85978
rect 65740 85926 65750 85978
rect 65750 85926 65796 85978
rect 65820 85926 65866 85978
rect 65866 85926 65876 85978
rect 65900 85926 65930 85978
rect 65930 85926 65956 85978
rect 65660 85924 65716 85926
rect 65740 85924 65796 85926
rect 65820 85924 65876 85926
rect 65900 85924 65956 85926
rect 65660 84890 65716 84892
rect 65740 84890 65796 84892
rect 65820 84890 65876 84892
rect 65900 84890 65956 84892
rect 65660 84838 65686 84890
rect 65686 84838 65716 84890
rect 65740 84838 65750 84890
rect 65750 84838 65796 84890
rect 65820 84838 65866 84890
rect 65866 84838 65876 84890
rect 65900 84838 65930 84890
rect 65930 84838 65956 84890
rect 65660 84836 65716 84838
rect 65740 84836 65796 84838
rect 65820 84836 65876 84838
rect 65900 84836 65956 84838
rect 65660 83802 65716 83804
rect 65740 83802 65796 83804
rect 65820 83802 65876 83804
rect 65900 83802 65956 83804
rect 65660 83750 65686 83802
rect 65686 83750 65716 83802
rect 65740 83750 65750 83802
rect 65750 83750 65796 83802
rect 65820 83750 65866 83802
rect 65866 83750 65876 83802
rect 65900 83750 65930 83802
rect 65930 83750 65956 83802
rect 65660 83748 65716 83750
rect 65740 83748 65796 83750
rect 65820 83748 65876 83750
rect 65900 83748 65956 83750
rect 65660 82714 65716 82716
rect 65740 82714 65796 82716
rect 65820 82714 65876 82716
rect 65900 82714 65956 82716
rect 65660 82662 65686 82714
rect 65686 82662 65716 82714
rect 65740 82662 65750 82714
rect 65750 82662 65796 82714
rect 65820 82662 65866 82714
rect 65866 82662 65876 82714
rect 65900 82662 65930 82714
rect 65930 82662 65956 82714
rect 65660 82660 65716 82662
rect 65740 82660 65796 82662
rect 65820 82660 65876 82662
rect 65900 82660 65956 82662
rect 65660 81626 65716 81628
rect 65740 81626 65796 81628
rect 65820 81626 65876 81628
rect 65900 81626 65956 81628
rect 65660 81574 65686 81626
rect 65686 81574 65716 81626
rect 65740 81574 65750 81626
rect 65750 81574 65796 81626
rect 65820 81574 65866 81626
rect 65866 81574 65876 81626
rect 65900 81574 65930 81626
rect 65930 81574 65956 81626
rect 65660 81572 65716 81574
rect 65740 81572 65796 81574
rect 65820 81572 65876 81574
rect 65900 81572 65956 81574
rect 65660 80538 65716 80540
rect 65740 80538 65796 80540
rect 65820 80538 65876 80540
rect 65900 80538 65956 80540
rect 65660 80486 65686 80538
rect 65686 80486 65716 80538
rect 65740 80486 65750 80538
rect 65750 80486 65796 80538
rect 65820 80486 65866 80538
rect 65866 80486 65876 80538
rect 65900 80486 65930 80538
rect 65930 80486 65956 80538
rect 65660 80484 65716 80486
rect 65740 80484 65796 80486
rect 65820 80484 65876 80486
rect 65900 80484 65956 80486
rect 65660 79450 65716 79452
rect 65740 79450 65796 79452
rect 65820 79450 65876 79452
rect 65900 79450 65956 79452
rect 65660 79398 65686 79450
rect 65686 79398 65716 79450
rect 65740 79398 65750 79450
rect 65750 79398 65796 79450
rect 65820 79398 65866 79450
rect 65866 79398 65876 79450
rect 65900 79398 65930 79450
rect 65930 79398 65956 79450
rect 65660 79396 65716 79398
rect 65740 79396 65796 79398
rect 65820 79396 65876 79398
rect 65900 79396 65956 79398
rect 65660 78362 65716 78364
rect 65740 78362 65796 78364
rect 65820 78362 65876 78364
rect 65900 78362 65956 78364
rect 65660 78310 65686 78362
rect 65686 78310 65716 78362
rect 65740 78310 65750 78362
rect 65750 78310 65796 78362
rect 65820 78310 65866 78362
rect 65866 78310 65876 78362
rect 65900 78310 65930 78362
rect 65930 78310 65956 78362
rect 65660 78308 65716 78310
rect 65740 78308 65796 78310
rect 65820 78308 65876 78310
rect 65900 78308 65956 78310
rect 65660 77274 65716 77276
rect 65740 77274 65796 77276
rect 65820 77274 65876 77276
rect 65900 77274 65956 77276
rect 65660 77222 65686 77274
rect 65686 77222 65716 77274
rect 65740 77222 65750 77274
rect 65750 77222 65796 77274
rect 65820 77222 65866 77274
rect 65866 77222 65876 77274
rect 65900 77222 65930 77274
rect 65930 77222 65956 77274
rect 65660 77220 65716 77222
rect 65740 77220 65796 77222
rect 65820 77220 65876 77222
rect 65900 77220 65956 77222
rect 65660 76186 65716 76188
rect 65740 76186 65796 76188
rect 65820 76186 65876 76188
rect 65900 76186 65956 76188
rect 65660 76134 65686 76186
rect 65686 76134 65716 76186
rect 65740 76134 65750 76186
rect 65750 76134 65796 76186
rect 65820 76134 65866 76186
rect 65866 76134 65876 76186
rect 65900 76134 65930 76186
rect 65930 76134 65956 76186
rect 65660 76132 65716 76134
rect 65740 76132 65796 76134
rect 65820 76132 65876 76134
rect 65900 76132 65956 76134
rect 65660 75098 65716 75100
rect 65740 75098 65796 75100
rect 65820 75098 65876 75100
rect 65900 75098 65956 75100
rect 65660 75046 65686 75098
rect 65686 75046 65716 75098
rect 65740 75046 65750 75098
rect 65750 75046 65796 75098
rect 65820 75046 65866 75098
rect 65866 75046 65876 75098
rect 65900 75046 65930 75098
rect 65930 75046 65956 75098
rect 65660 75044 65716 75046
rect 65740 75044 65796 75046
rect 65820 75044 65876 75046
rect 65900 75044 65956 75046
rect 65660 74010 65716 74012
rect 65740 74010 65796 74012
rect 65820 74010 65876 74012
rect 65900 74010 65956 74012
rect 65660 73958 65686 74010
rect 65686 73958 65716 74010
rect 65740 73958 65750 74010
rect 65750 73958 65796 74010
rect 65820 73958 65866 74010
rect 65866 73958 65876 74010
rect 65900 73958 65930 74010
rect 65930 73958 65956 74010
rect 65660 73956 65716 73958
rect 65740 73956 65796 73958
rect 65820 73956 65876 73958
rect 65900 73956 65956 73958
rect 65660 72922 65716 72924
rect 65740 72922 65796 72924
rect 65820 72922 65876 72924
rect 65900 72922 65956 72924
rect 65660 72870 65686 72922
rect 65686 72870 65716 72922
rect 65740 72870 65750 72922
rect 65750 72870 65796 72922
rect 65820 72870 65866 72922
rect 65866 72870 65876 72922
rect 65900 72870 65930 72922
rect 65930 72870 65956 72922
rect 65660 72868 65716 72870
rect 65740 72868 65796 72870
rect 65820 72868 65876 72870
rect 65900 72868 65956 72870
rect 65660 71834 65716 71836
rect 65740 71834 65796 71836
rect 65820 71834 65876 71836
rect 65900 71834 65956 71836
rect 65660 71782 65686 71834
rect 65686 71782 65716 71834
rect 65740 71782 65750 71834
rect 65750 71782 65796 71834
rect 65820 71782 65866 71834
rect 65866 71782 65876 71834
rect 65900 71782 65930 71834
rect 65930 71782 65956 71834
rect 65660 71780 65716 71782
rect 65740 71780 65796 71782
rect 65820 71780 65876 71782
rect 65900 71780 65956 71782
rect 65660 70746 65716 70748
rect 65740 70746 65796 70748
rect 65820 70746 65876 70748
rect 65900 70746 65956 70748
rect 65660 70694 65686 70746
rect 65686 70694 65716 70746
rect 65740 70694 65750 70746
rect 65750 70694 65796 70746
rect 65820 70694 65866 70746
rect 65866 70694 65876 70746
rect 65900 70694 65930 70746
rect 65930 70694 65956 70746
rect 65660 70692 65716 70694
rect 65740 70692 65796 70694
rect 65820 70692 65876 70694
rect 65900 70692 65956 70694
rect 65660 69658 65716 69660
rect 65740 69658 65796 69660
rect 65820 69658 65876 69660
rect 65900 69658 65956 69660
rect 65660 69606 65686 69658
rect 65686 69606 65716 69658
rect 65740 69606 65750 69658
rect 65750 69606 65796 69658
rect 65820 69606 65866 69658
rect 65866 69606 65876 69658
rect 65900 69606 65930 69658
rect 65930 69606 65956 69658
rect 65660 69604 65716 69606
rect 65740 69604 65796 69606
rect 65820 69604 65876 69606
rect 65900 69604 65956 69606
rect 65660 68570 65716 68572
rect 65740 68570 65796 68572
rect 65820 68570 65876 68572
rect 65900 68570 65956 68572
rect 65660 68518 65686 68570
rect 65686 68518 65716 68570
rect 65740 68518 65750 68570
rect 65750 68518 65796 68570
rect 65820 68518 65866 68570
rect 65866 68518 65876 68570
rect 65900 68518 65930 68570
rect 65930 68518 65956 68570
rect 65660 68516 65716 68518
rect 65740 68516 65796 68518
rect 65820 68516 65876 68518
rect 65900 68516 65956 68518
rect 65660 67482 65716 67484
rect 65740 67482 65796 67484
rect 65820 67482 65876 67484
rect 65900 67482 65956 67484
rect 65660 67430 65686 67482
rect 65686 67430 65716 67482
rect 65740 67430 65750 67482
rect 65750 67430 65796 67482
rect 65820 67430 65866 67482
rect 65866 67430 65876 67482
rect 65900 67430 65930 67482
rect 65930 67430 65956 67482
rect 65660 67428 65716 67430
rect 65740 67428 65796 67430
rect 65820 67428 65876 67430
rect 65900 67428 65956 67430
rect 65660 66394 65716 66396
rect 65740 66394 65796 66396
rect 65820 66394 65876 66396
rect 65900 66394 65956 66396
rect 65660 66342 65686 66394
rect 65686 66342 65716 66394
rect 65740 66342 65750 66394
rect 65750 66342 65796 66394
rect 65820 66342 65866 66394
rect 65866 66342 65876 66394
rect 65900 66342 65930 66394
rect 65930 66342 65956 66394
rect 65660 66340 65716 66342
rect 65740 66340 65796 66342
rect 65820 66340 65876 66342
rect 65900 66340 65956 66342
rect 65660 65306 65716 65308
rect 65740 65306 65796 65308
rect 65820 65306 65876 65308
rect 65900 65306 65956 65308
rect 65660 65254 65686 65306
rect 65686 65254 65716 65306
rect 65740 65254 65750 65306
rect 65750 65254 65796 65306
rect 65820 65254 65866 65306
rect 65866 65254 65876 65306
rect 65900 65254 65930 65306
rect 65930 65254 65956 65306
rect 65660 65252 65716 65254
rect 65740 65252 65796 65254
rect 65820 65252 65876 65254
rect 65900 65252 65956 65254
rect 65660 64218 65716 64220
rect 65740 64218 65796 64220
rect 65820 64218 65876 64220
rect 65900 64218 65956 64220
rect 65660 64166 65686 64218
rect 65686 64166 65716 64218
rect 65740 64166 65750 64218
rect 65750 64166 65796 64218
rect 65820 64166 65866 64218
rect 65866 64166 65876 64218
rect 65900 64166 65930 64218
rect 65930 64166 65956 64218
rect 65660 64164 65716 64166
rect 65740 64164 65796 64166
rect 65820 64164 65876 64166
rect 65900 64164 65956 64166
rect 65660 63130 65716 63132
rect 65740 63130 65796 63132
rect 65820 63130 65876 63132
rect 65900 63130 65956 63132
rect 65660 63078 65686 63130
rect 65686 63078 65716 63130
rect 65740 63078 65750 63130
rect 65750 63078 65796 63130
rect 65820 63078 65866 63130
rect 65866 63078 65876 63130
rect 65900 63078 65930 63130
rect 65930 63078 65956 63130
rect 65660 63076 65716 63078
rect 65740 63076 65796 63078
rect 65820 63076 65876 63078
rect 65900 63076 65956 63078
rect 65660 62042 65716 62044
rect 65740 62042 65796 62044
rect 65820 62042 65876 62044
rect 65900 62042 65956 62044
rect 65660 61990 65686 62042
rect 65686 61990 65716 62042
rect 65740 61990 65750 62042
rect 65750 61990 65796 62042
rect 65820 61990 65866 62042
rect 65866 61990 65876 62042
rect 65900 61990 65930 62042
rect 65930 61990 65956 62042
rect 65660 61988 65716 61990
rect 65740 61988 65796 61990
rect 65820 61988 65876 61990
rect 65900 61988 65956 61990
rect 65660 60954 65716 60956
rect 65740 60954 65796 60956
rect 65820 60954 65876 60956
rect 65900 60954 65956 60956
rect 65660 60902 65686 60954
rect 65686 60902 65716 60954
rect 65740 60902 65750 60954
rect 65750 60902 65796 60954
rect 65820 60902 65866 60954
rect 65866 60902 65876 60954
rect 65900 60902 65930 60954
rect 65930 60902 65956 60954
rect 65660 60900 65716 60902
rect 65740 60900 65796 60902
rect 65820 60900 65876 60902
rect 65900 60900 65956 60902
rect 65660 59866 65716 59868
rect 65740 59866 65796 59868
rect 65820 59866 65876 59868
rect 65900 59866 65956 59868
rect 65660 59814 65686 59866
rect 65686 59814 65716 59866
rect 65740 59814 65750 59866
rect 65750 59814 65796 59866
rect 65820 59814 65866 59866
rect 65866 59814 65876 59866
rect 65900 59814 65930 59866
rect 65930 59814 65956 59866
rect 65660 59812 65716 59814
rect 65740 59812 65796 59814
rect 65820 59812 65876 59814
rect 65900 59812 65956 59814
rect 65660 58778 65716 58780
rect 65740 58778 65796 58780
rect 65820 58778 65876 58780
rect 65900 58778 65956 58780
rect 65660 58726 65686 58778
rect 65686 58726 65716 58778
rect 65740 58726 65750 58778
rect 65750 58726 65796 58778
rect 65820 58726 65866 58778
rect 65866 58726 65876 58778
rect 65900 58726 65930 58778
rect 65930 58726 65956 58778
rect 65660 58724 65716 58726
rect 65740 58724 65796 58726
rect 65820 58724 65876 58726
rect 65900 58724 65956 58726
rect 65660 57690 65716 57692
rect 65740 57690 65796 57692
rect 65820 57690 65876 57692
rect 65900 57690 65956 57692
rect 65660 57638 65686 57690
rect 65686 57638 65716 57690
rect 65740 57638 65750 57690
rect 65750 57638 65796 57690
rect 65820 57638 65866 57690
rect 65866 57638 65876 57690
rect 65900 57638 65930 57690
rect 65930 57638 65956 57690
rect 65660 57636 65716 57638
rect 65740 57636 65796 57638
rect 65820 57636 65876 57638
rect 65900 57636 65956 57638
rect 65660 56602 65716 56604
rect 65740 56602 65796 56604
rect 65820 56602 65876 56604
rect 65900 56602 65956 56604
rect 65660 56550 65686 56602
rect 65686 56550 65716 56602
rect 65740 56550 65750 56602
rect 65750 56550 65796 56602
rect 65820 56550 65866 56602
rect 65866 56550 65876 56602
rect 65900 56550 65930 56602
rect 65930 56550 65956 56602
rect 65660 56548 65716 56550
rect 65740 56548 65796 56550
rect 65820 56548 65876 56550
rect 65900 56548 65956 56550
rect 65660 55514 65716 55516
rect 65740 55514 65796 55516
rect 65820 55514 65876 55516
rect 65900 55514 65956 55516
rect 65660 55462 65686 55514
rect 65686 55462 65716 55514
rect 65740 55462 65750 55514
rect 65750 55462 65796 55514
rect 65820 55462 65866 55514
rect 65866 55462 65876 55514
rect 65900 55462 65930 55514
rect 65930 55462 65956 55514
rect 65660 55460 65716 55462
rect 65740 55460 65796 55462
rect 65820 55460 65876 55462
rect 65900 55460 65956 55462
rect 65660 54426 65716 54428
rect 65740 54426 65796 54428
rect 65820 54426 65876 54428
rect 65900 54426 65956 54428
rect 65660 54374 65686 54426
rect 65686 54374 65716 54426
rect 65740 54374 65750 54426
rect 65750 54374 65796 54426
rect 65820 54374 65866 54426
rect 65866 54374 65876 54426
rect 65900 54374 65930 54426
rect 65930 54374 65956 54426
rect 65660 54372 65716 54374
rect 65740 54372 65796 54374
rect 65820 54372 65876 54374
rect 65900 54372 65956 54374
rect 65660 53338 65716 53340
rect 65740 53338 65796 53340
rect 65820 53338 65876 53340
rect 65900 53338 65956 53340
rect 65660 53286 65686 53338
rect 65686 53286 65716 53338
rect 65740 53286 65750 53338
rect 65750 53286 65796 53338
rect 65820 53286 65866 53338
rect 65866 53286 65876 53338
rect 65900 53286 65930 53338
rect 65930 53286 65956 53338
rect 65660 53284 65716 53286
rect 65740 53284 65796 53286
rect 65820 53284 65876 53286
rect 65900 53284 65956 53286
rect 65660 52250 65716 52252
rect 65740 52250 65796 52252
rect 65820 52250 65876 52252
rect 65900 52250 65956 52252
rect 65660 52198 65686 52250
rect 65686 52198 65716 52250
rect 65740 52198 65750 52250
rect 65750 52198 65796 52250
rect 65820 52198 65866 52250
rect 65866 52198 65876 52250
rect 65900 52198 65930 52250
rect 65930 52198 65956 52250
rect 65660 52196 65716 52198
rect 65740 52196 65796 52198
rect 65820 52196 65876 52198
rect 65900 52196 65956 52198
rect 65660 51162 65716 51164
rect 65740 51162 65796 51164
rect 65820 51162 65876 51164
rect 65900 51162 65956 51164
rect 65660 51110 65686 51162
rect 65686 51110 65716 51162
rect 65740 51110 65750 51162
rect 65750 51110 65796 51162
rect 65820 51110 65866 51162
rect 65866 51110 65876 51162
rect 65900 51110 65930 51162
rect 65930 51110 65956 51162
rect 65660 51108 65716 51110
rect 65740 51108 65796 51110
rect 65820 51108 65876 51110
rect 65900 51108 65956 51110
rect 65660 50074 65716 50076
rect 65740 50074 65796 50076
rect 65820 50074 65876 50076
rect 65900 50074 65956 50076
rect 65660 50022 65686 50074
rect 65686 50022 65716 50074
rect 65740 50022 65750 50074
rect 65750 50022 65796 50074
rect 65820 50022 65866 50074
rect 65866 50022 65876 50074
rect 65900 50022 65930 50074
rect 65930 50022 65956 50074
rect 65660 50020 65716 50022
rect 65740 50020 65796 50022
rect 65820 50020 65876 50022
rect 65900 50020 65956 50022
rect 65660 48986 65716 48988
rect 65740 48986 65796 48988
rect 65820 48986 65876 48988
rect 65900 48986 65956 48988
rect 65660 48934 65686 48986
rect 65686 48934 65716 48986
rect 65740 48934 65750 48986
rect 65750 48934 65796 48986
rect 65820 48934 65866 48986
rect 65866 48934 65876 48986
rect 65900 48934 65930 48986
rect 65930 48934 65956 48986
rect 65660 48932 65716 48934
rect 65740 48932 65796 48934
rect 65820 48932 65876 48934
rect 65900 48932 65956 48934
rect 65660 47898 65716 47900
rect 65740 47898 65796 47900
rect 65820 47898 65876 47900
rect 65900 47898 65956 47900
rect 65660 47846 65686 47898
rect 65686 47846 65716 47898
rect 65740 47846 65750 47898
rect 65750 47846 65796 47898
rect 65820 47846 65866 47898
rect 65866 47846 65876 47898
rect 65900 47846 65930 47898
rect 65930 47846 65956 47898
rect 65660 47844 65716 47846
rect 65740 47844 65796 47846
rect 65820 47844 65876 47846
rect 65900 47844 65956 47846
rect 65660 46810 65716 46812
rect 65740 46810 65796 46812
rect 65820 46810 65876 46812
rect 65900 46810 65956 46812
rect 65660 46758 65686 46810
rect 65686 46758 65716 46810
rect 65740 46758 65750 46810
rect 65750 46758 65796 46810
rect 65820 46758 65866 46810
rect 65866 46758 65876 46810
rect 65900 46758 65930 46810
rect 65930 46758 65956 46810
rect 65660 46756 65716 46758
rect 65740 46756 65796 46758
rect 65820 46756 65876 46758
rect 65900 46756 65956 46758
rect 65660 45722 65716 45724
rect 65740 45722 65796 45724
rect 65820 45722 65876 45724
rect 65900 45722 65956 45724
rect 65660 45670 65686 45722
rect 65686 45670 65716 45722
rect 65740 45670 65750 45722
rect 65750 45670 65796 45722
rect 65820 45670 65866 45722
rect 65866 45670 65876 45722
rect 65900 45670 65930 45722
rect 65930 45670 65956 45722
rect 65660 45668 65716 45670
rect 65740 45668 65796 45670
rect 65820 45668 65876 45670
rect 65900 45668 65956 45670
rect 65660 44634 65716 44636
rect 65740 44634 65796 44636
rect 65820 44634 65876 44636
rect 65900 44634 65956 44636
rect 65660 44582 65686 44634
rect 65686 44582 65716 44634
rect 65740 44582 65750 44634
rect 65750 44582 65796 44634
rect 65820 44582 65866 44634
rect 65866 44582 65876 44634
rect 65900 44582 65930 44634
rect 65930 44582 65956 44634
rect 65660 44580 65716 44582
rect 65740 44580 65796 44582
rect 65820 44580 65876 44582
rect 65900 44580 65956 44582
rect 65660 43546 65716 43548
rect 65740 43546 65796 43548
rect 65820 43546 65876 43548
rect 65900 43546 65956 43548
rect 65660 43494 65686 43546
rect 65686 43494 65716 43546
rect 65740 43494 65750 43546
rect 65750 43494 65796 43546
rect 65820 43494 65866 43546
rect 65866 43494 65876 43546
rect 65900 43494 65930 43546
rect 65930 43494 65956 43546
rect 65660 43492 65716 43494
rect 65740 43492 65796 43494
rect 65820 43492 65876 43494
rect 65900 43492 65956 43494
rect 65660 42458 65716 42460
rect 65740 42458 65796 42460
rect 65820 42458 65876 42460
rect 65900 42458 65956 42460
rect 65660 42406 65686 42458
rect 65686 42406 65716 42458
rect 65740 42406 65750 42458
rect 65750 42406 65796 42458
rect 65820 42406 65866 42458
rect 65866 42406 65876 42458
rect 65900 42406 65930 42458
rect 65930 42406 65956 42458
rect 65660 42404 65716 42406
rect 65740 42404 65796 42406
rect 65820 42404 65876 42406
rect 65900 42404 65956 42406
rect 65660 41370 65716 41372
rect 65740 41370 65796 41372
rect 65820 41370 65876 41372
rect 65900 41370 65956 41372
rect 65660 41318 65686 41370
rect 65686 41318 65716 41370
rect 65740 41318 65750 41370
rect 65750 41318 65796 41370
rect 65820 41318 65866 41370
rect 65866 41318 65876 41370
rect 65900 41318 65930 41370
rect 65930 41318 65956 41370
rect 65660 41316 65716 41318
rect 65740 41316 65796 41318
rect 65820 41316 65876 41318
rect 65900 41316 65956 41318
rect 65660 40282 65716 40284
rect 65740 40282 65796 40284
rect 65820 40282 65876 40284
rect 65900 40282 65956 40284
rect 65660 40230 65686 40282
rect 65686 40230 65716 40282
rect 65740 40230 65750 40282
rect 65750 40230 65796 40282
rect 65820 40230 65866 40282
rect 65866 40230 65876 40282
rect 65900 40230 65930 40282
rect 65930 40230 65956 40282
rect 65660 40228 65716 40230
rect 65740 40228 65796 40230
rect 65820 40228 65876 40230
rect 65900 40228 65956 40230
rect 65660 39194 65716 39196
rect 65740 39194 65796 39196
rect 65820 39194 65876 39196
rect 65900 39194 65956 39196
rect 65660 39142 65686 39194
rect 65686 39142 65716 39194
rect 65740 39142 65750 39194
rect 65750 39142 65796 39194
rect 65820 39142 65866 39194
rect 65866 39142 65876 39194
rect 65900 39142 65930 39194
rect 65930 39142 65956 39194
rect 65660 39140 65716 39142
rect 65740 39140 65796 39142
rect 65820 39140 65876 39142
rect 65900 39140 65956 39142
rect 65660 38106 65716 38108
rect 65740 38106 65796 38108
rect 65820 38106 65876 38108
rect 65900 38106 65956 38108
rect 65660 38054 65686 38106
rect 65686 38054 65716 38106
rect 65740 38054 65750 38106
rect 65750 38054 65796 38106
rect 65820 38054 65866 38106
rect 65866 38054 65876 38106
rect 65900 38054 65930 38106
rect 65930 38054 65956 38106
rect 65660 38052 65716 38054
rect 65740 38052 65796 38054
rect 65820 38052 65876 38054
rect 65900 38052 65956 38054
rect 65660 37018 65716 37020
rect 65740 37018 65796 37020
rect 65820 37018 65876 37020
rect 65900 37018 65956 37020
rect 65660 36966 65686 37018
rect 65686 36966 65716 37018
rect 65740 36966 65750 37018
rect 65750 36966 65796 37018
rect 65820 36966 65866 37018
rect 65866 36966 65876 37018
rect 65900 36966 65930 37018
rect 65930 36966 65956 37018
rect 65660 36964 65716 36966
rect 65740 36964 65796 36966
rect 65820 36964 65876 36966
rect 65900 36964 65956 36966
rect 65660 35930 65716 35932
rect 65740 35930 65796 35932
rect 65820 35930 65876 35932
rect 65900 35930 65956 35932
rect 65660 35878 65686 35930
rect 65686 35878 65716 35930
rect 65740 35878 65750 35930
rect 65750 35878 65796 35930
rect 65820 35878 65866 35930
rect 65866 35878 65876 35930
rect 65900 35878 65930 35930
rect 65930 35878 65956 35930
rect 65660 35876 65716 35878
rect 65740 35876 65796 35878
rect 65820 35876 65876 35878
rect 65900 35876 65956 35878
rect 65660 34842 65716 34844
rect 65740 34842 65796 34844
rect 65820 34842 65876 34844
rect 65900 34842 65956 34844
rect 65660 34790 65686 34842
rect 65686 34790 65716 34842
rect 65740 34790 65750 34842
rect 65750 34790 65796 34842
rect 65820 34790 65866 34842
rect 65866 34790 65876 34842
rect 65900 34790 65930 34842
rect 65930 34790 65956 34842
rect 65660 34788 65716 34790
rect 65740 34788 65796 34790
rect 65820 34788 65876 34790
rect 65900 34788 65956 34790
rect 65660 33754 65716 33756
rect 65740 33754 65796 33756
rect 65820 33754 65876 33756
rect 65900 33754 65956 33756
rect 65660 33702 65686 33754
rect 65686 33702 65716 33754
rect 65740 33702 65750 33754
rect 65750 33702 65796 33754
rect 65820 33702 65866 33754
rect 65866 33702 65876 33754
rect 65900 33702 65930 33754
rect 65930 33702 65956 33754
rect 65660 33700 65716 33702
rect 65740 33700 65796 33702
rect 65820 33700 65876 33702
rect 65900 33700 65956 33702
rect 65660 32666 65716 32668
rect 65740 32666 65796 32668
rect 65820 32666 65876 32668
rect 65900 32666 65956 32668
rect 65660 32614 65686 32666
rect 65686 32614 65716 32666
rect 65740 32614 65750 32666
rect 65750 32614 65796 32666
rect 65820 32614 65866 32666
rect 65866 32614 65876 32666
rect 65900 32614 65930 32666
rect 65930 32614 65956 32666
rect 65660 32612 65716 32614
rect 65740 32612 65796 32614
rect 65820 32612 65876 32614
rect 65900 32612 65956 32614
rect 65660 31578 65716 31580
rect 65740 31578 65796 31580
rect 65820 31578 65876 31580
rect 65900 31578 65956 31580
rect 65660 31526 65686 31578
rect 65686 31526 65716 31578
rect 65740 31526 65750 31578
rect 65750 31526 65796 31578
rect 65820 31526 65866 31578
rect 65866 31526 65876 31578
rect 65900 31526 65930 31578
rect 65930 31526 65956 31578
rect 65660 31524 65716 31526
rect 65740 31524 65796 31526
rect 65820 31524 65876 31526
rect 65900 31524 65956 31526
rect 65660 30490 65716 30492
rect 65740 30490 65796 30492
rect 65820 30490 65876 30492
rect 65900 30490 65956 30492
rect 65660 30438 65686 30490
rect 65686 30438 65716 30490
rect 65740 30438 65750 30490
rect 65750 30438 65796 30490
rect 65820 30438 65866 30490
rect 65866 30438 65876 30490
rect 65900 30438 65930 30490
rect 65930 30438 65956 30490
rect 65660 30436 65716 30438
rect 65740 30436 65796 30438
rect 65820 30436 65876 30438
rect 65900 30436 65956 30438
rect 65660 29402 65716 29404
rect 65740 29402 65796 29404
rect 65820 29402 65876 29404
rect 65900 29402 65956 29404
rect 65660 29350 65686 29402
rect 65686 29350 65716 29402
rect 65740 29350 65750 29402
rect 65750 29350 65796 29402
rect 65820 29350 65866 29402
rect 65866 29350 65876 29402
rect 65900 29350 65930 29402
rect 65930 29350 65956 29402
rect 65660 29348 65716 29350
rect 65740 29348 65796 29350
rect 65820 29348 65876 29350
rect 65900 29348 65956 29350
rect 65660 28314 65716 28316
rect 65740 28314 65796 28316
rect 65820 28314 65876 28316
rect 65900 28314 65956 28316
rect 65660 28262 65686 28314
rect 65686 28262 65716 28314
rect 65740 28262 65750 28314
rect 65750 28262 65796 28314
rect 65820 28262 65866 28314
rect 65866 28262 65876 28314
rect 65900 28262 65930 28314
rect 65930 28262 65956 28314
rect 65660 28260 65716 28262
rect 65740 28260 65796 28262
rect 65820 28260 65876 28262
rect 65900 28260 65956 28262
rect 65660 27226 65716 27228
rect 65740 27226 65796 27228
rect 65820 27226 65876 27228
rect 65900 27226 65956 27228
rect 65660 27174 65686 27226
rect 65686 27174 65716 27226
rect 65740 27174 65750 27226
rect 65750 27174 65796 27226
rect 65820 27174 65866 27226
rect 65866 27174 65876 27226
rect 65900 27174 65930 27226
rect 65930 27174 65956 27226
rect 65660 27172 65716 27174
rect 65740 27172 65796 27174
rect 65820 27172 65876 27174
rect 65900 27172 65956 27174
rect 65660 26138 65716 26140
rect 65740 26138 65796 26140
rect 65820 26138 65876 26140
rect 65900 26138 65956 26140
rect 65660 26086 65686 26138
rect 65686 26086 65716 26138
rect 65740 26086 65750 26138
rect 65750 26086 65796 26138
rect 65820 26086 65866 26138
rect 65866 26086 65876 26138
rect 65900 26086 65930 26138
rect 65930 26086 65956 26138
rect 65660 26084 65716 26086
rect 65740 26084 65796 26086
rect 65820 26084 65876 26086
rect 65900 26084 65956 26086
rect 65660 25050 65716 25052
rect 65740 25050 65796 25052
rect 65820 25050 65876 25052
rect 65900 25050 65956 25052
rect 65660 24998 65686 25050
rect 65686 24998 65716 25050
rect 65740 24998 65750 25050
rect 65750 24998 65796 25050
rect 65820 24998 65866 25050
rect 65866 24998 65876 25050
rect 65900 24998 65930 25050
rect 65930 24998 65956 25050
rect 65660 24996 65716 24998
rect 65740 24996 65796 24998
rect 65820 24996 65876 24998
rect 65900 24996 65956 24998
rect 65660 23962 65716 23964
rect 65740 23962 65796 23964
rect 65820 23962 65876 23964
rect 65900 23962 65956 23964
rect 65660 23910 65686 23962
rect 65686 23910 65716 23962
rect 65740 23910 65750 23962
rect 65750 23910 65796 23962
rect 65820 23910 65866 23962
rect 65866 23910 65876 23962
rect 65900 23910 65930 23962
rect 65930 23910 65956 23962
rect 65660 23908 65716 23910
rect 65740 23908 65796 23910
rect 65820 23908 65876 23910
rect 65900 23908 65956 23910
rect 65660 22874 65716 22876
rect 65740 22874 65796 22876
rect 65820 22874 65876 22876
rect 65900 22874 65956 22876
rect 65660 22822 65686 22874
rect 65686 22822 65716 22874
rect 65740 22822 65750 22874
rect 65750 22822 65796 22874
rect 65820 22822 65866 22874
rect 65866 22822 65876 22874
rect 65900 22822 65930 22874
rect 65930 22822 65956 22874
rect 65660 22820 65716 22822
rect 65740 22820 65796 22822
rect 65820 22820 65876 22822
rect 65900 22820 65956 22822
rect 65660 21786 65716 21788
rect 65740 21786 65796 21788
rect 65820 21786 65876 21788
rect 65900 21786 65956 21788
rect 65660 21734 65686 21786
rect 65686 21734 65716 21786
rect 65740 21734 65750 21786
rect 65750 21734 65796 21786
rect 65820 21734 65866 21786
rect 65866 21734 65876 21786
rect 65900 21734 65930 21786
rect 65930 21734 65956 21786
rect 65660 21732 65716 21734
rect 65740 21732 65796 21734
rect 65820 21732 65876 21734
rect 65900 21732 65956 21734
rect 65660 20698 65716 20700
rect 65740 20698 65796 20700
rect 65820 20698 65876 20700
rect 65900 20698 65956 20700
rect 65660 20646 65686 20698
rect 65686 20646 65716 20698
rect 65740 20646 65750 20698
rect 65750 20646 65796 20698
rect 65820 20646 65866 20698
rect 65866 20646 65876 20698
rect 65900 20646 65930 20698
rect 65930 20646 65956 20698
rect 65660 20644 65716 20646
rect 65740 20644 65796 20646
rect 65820 20644 65876 20646
rect 65900 20644 65956 20646
rect 65660 19610 65716 19612
rect 65740 19610 65796 19612
rect 65820 19610 65876 19612
rect 65900 19610 65956 19612
rect 65660 19558 65686 19610
rect 65686 19558 65716 19610
rect 65740 19558 65750 19610
rect 65750 19558 65796 19610
rect 65820 19558 65866 19610
rect 65866 19558 65876 19610
rect 65900 19558 65930 19610
rect 65930 19558 65956 19610
rect 65660 19556 65716 19558
rect 65740 19556 65796 19558
rect 65820 19556 65876 19558
rect 65900 19556 65956 19558
rect 65660 18522 65716 18524
rect 65740 18522 65796 18524
rect 65820 18522 65876 18524
rect 65900 18522 65956 18524
rect 65660 18470 65686 18522
rect 65686 18470 65716 18522
rect 65740 18470 65750 18522
rect 65750 18470 65796 18522
rect 65820 18470 65866 18522
rect 65866 18470 65876 18522
rect 65900 18470 65930 18522
rect 65930 18470 65956 18522
rect 65660 18468 65716 18470
rect 65740 18468 65796 18470
rect 65820 18468 65876 18470
rect 65900 18468 65956 18470
rect 65660 17434 65716 17436
rect 65740 17434 65796 17436
rect 65820 17434 65876 17436
rect 65900 17434 65956 17436
rect 65660 17382 65686 17434
rect 65686 17382 65716 17434
rect 65740 17382 65750 17434
rect 65750 17382 65796 17434
rect 65820 17382 65866 17434
rect 65866 17382 65876 17434
rect 65900 17382 65930 17434
rect 65930 17382 65956 17434
rect 65660 17380 65716 17382
rect 65740 17380 65796 17382
rect 65820 17380 65876 17382
rect 65900 17380 65956 17382
rect 61198 7148 61200 7168
rect 61200 7148 61252 7168
rect 61252 7148 61254 7168
rect 61198 7112 61254 7148
rect 61566 7268 61622 7304
rect 61566 7248 61568 7268
rect 61568 7248 61620 7268
rect 61620 7248 61622 7268
rect 60646 6316 60702 6352
rect 60646 6296 60648 6316
rect 60648 6296 60700 6316
rect 60700 6296 60702 6316
rect 61566 6568 61622 6624
rect 61014 5480 61070 5536
rect 62302 7404 62358 7440
rect 62302 7384 62331 7404
rect 62331 7384 62358 7404
rect 62026 6996 62082 7032
rect 62026 6976 62028 6996
rect 62028 6976 62080 6996
rect 62080 6976 62082 6996
rect 62578 7812 62634 7848
rect 62578 7792 62580 7812
rect 62580 7792 62632 7812
rect 62632 7792 62634 7812
rect 62394 6704 62450 6760
rect 63130 6452 63186 6488
rect 63130 6432 63132 6452
rect 63132 6432 63184 6452
rect 63184 6432 63186 6452
rect 63130 5908 63186 5944
rect 63130 5888 63132 5908
rect 63132 5888 63184 5908
rect 63184 5888 63186 5908
rect 63314 7404 63370 7440
rect 63314 7384 63316 7404
rect 63316 7384 63368 7404
rect 63368 7384 63370 7404
rect 63314 6724 63370 6760
rect 63314 6704 63316 6724
rect 63316 6704 63368 6724
rect 63368 6704 63370 6724
rect 63406 5616 63462 5672
rect 63866 7248 63922 7304
rect 64234 7812 64290 7848
rect 64234 7792 64236 7812
rect 64236 7792 64288 7812
rect 64288 7792 64290 7812
rect 64418 6840 64474 6896
rect 65660 16346 65716 16348
rect 65740 16346 65796 16348
rect 65820 16346 65876 16348
rect 65900 16346 65956 16348
rect 65660 16294 65686 16346
rect 65686 16294 65716 16346
rect 65740 16294 65750 16346
rect 65750 16294 65796 16346
rect 65820 16294 65866 16346
rect 65866 16294 65876 16346
rect 65900 16294 65930 16346
rect 65930 16294 65956 16346
rect 65660 16292 65716 16294
rect 65740 16292 65796 16294
rect 65820 16292 65876 16294
rect 65900 16292 65956 16294
rect 65660 15258 65716 15260
rect 65740 15258 65796 15260
rect 65820 15258 65876 15260
rect 65900 15258 65956 15260
rect 65660 15206 65686 15258
rect 65686 15206 65716 15258
rect 65740 15206 65750 15258
rect 65750 15206 65796 15258
rect 65820 15206 65866 15258
rect 65866 15206 65876 15258
rect 65900 15206 65930 15258
rect 65930 15206 65956 15258
rect 65660 15204 65716 15206
rect 65740 15204 65796 15206
rect 65820 15204 65876 15206
rect 65900 15204 65956 15206
rect 65660 14170 65716 14172
rect 65740 14170 65796 14172
rect 65820 14170 65876 14172
rect 65900 14170 65956 14172
rect 65660 14118 65686 14170
rect 65686 14118 65716 14170
rect 65740 14118 65750 14170
rect 65750 14118 65796 14170
rect 65820 14118 65866 14170
rect 65866 14118 65876 14170
rect 65900 14118 65930 14170
rect 65930 14118 65956 14170
rect 65660 14116 65716 14118
rect 65740 14116 65796 14118
rect 65820 14116 65876 14118
rect 65900 14116 65956 14118
rect 65660 13082 65716 13084
rect 65740 13082 65796 13084
rect 65820 13082 65876 13084
rect 65900 13082 65956 13084
rect 65660 13030 65686 13082
rect 65686 13030 65716 13082
rect 65740 13030 65750 13082
rect 65750 13030 65796 13082
rect 65820 13030 65866 13082
rect 65866 13030 65876 13082
rect 65900 13030 65930 13082
rect 65930 13030 65956 13082
rect 65660 13028 65716 13030
rect 65740 13028 65796 13030
rect 65820 13028 65876 13030
rect 65900 13028 65956 13030
rect 64786 6840 64842 6896
rect 65154 7112 65210 7168
rect 64602 6296 64658 6352
rect 64418 6024 64474 6080
rect 64234 5772 64290 5808
rect 64234 5752 64236 5772
rect 64236 5752 64288 5772
rect 64288 5752 64290 5772
rect 64602 5636 64658 5672
rect 64602 5616 64604 5636
rect 64604 5616 64656 5636
rect 64656 5616 64658 5636
rect 65660 11994 65716 11996
rect 65740 11994 65796 11996
rect 65820 11994 65876 11996
rect 65900 11994 65956 11996
rect 65660 11942 65686 11994
rect 65686 11942 65716 11994
rect 65740 11942 65750 11994
rect 65750 11942 65796 11994
rect 65820 11942 65866 11994
rect 65866 11942 65876 11994
rect 65900 11942 65930 11994
rect 65930 11942 65956 11994
rect 65660 11940 65716 11942
rect 65740 11940 65796 11942
rect 65820 11940 65876 11942
rect 65900 11940 65956 11942
rect 65660 10906 65716 10908
rect 65740 10906 65796 10908
rect 65820 10906 65876 10908
rect 65900 10906 65956 10908
rect 65660 10854 65686 10906
rect 65686 10854 65716 10906
rect 65740 10854 65750 10906
rect 65750 10854 65796 10906
rect 65820 10854 65866 10906
rect 65866 10854 65876 10906
rect 65900 10854 65930 10906
rect 65930 10854 65956 10906
rect 65660 10852 65716 10854
rect 65740 10852 65796 10854
rect 65820 10852 65876 10854
rect 65900 10852 65956 10854
rect 65660 9818 65716 9820
rect 65740 9818 65796 9820
rect 65820 9818 65876 9820
rect 65900 9818 65956 9820
rect 65660 9766 65686 9818
rect 65686 9766 65716 9818
rect 65740 9766 65750 9818
rect 65750 9766 65796 9818
rect 65820 9766 65866 9818
rect 65866 9766 65876 9818
rect 65900 9766 65930 9818
rect 65930 9766 65956 9818
rect 65660 9764 65716 9766
rect 65740 9764 65796 9766
rect 65820 9764 65876 9766
rect 65900 9764 65956 9766
rect 65660 8730 65716 8732
rect 65740 8730 65796 8732
rect 65820 8730 65876 8732
rect 65900 8730 65956 8732
rect 65660 8678 65686 8730
rect 65686 8678 65716 8730
rect 65740 8678 65750 8730
rect 65750 8678 65796 8730
rect 65820 8678 65866 8730
rect 65866 8678 65876 8730
rect 65900 8678 65930 8730
rect 65930 8678 65956 8730
rect 65660 8676 65716 8678
rect 65740 8676 65796 8678
rect 65820 8676 65876 8678
rect 65900 8676 65956 8678
rect 65338 7112 65394 7168
rect 65246 5908 65302 5944
rect 65246 5888 65248 5908
rect 65248 5888 65300 5908
rect 65300 5888 65302 5908
rect 65246 5752 65302 5808
rect 65660 7642 65716 7644
rect 65740 7642 65796 7644
rect 65820 7642 65876 7644
rect 65900 7642 65956 7644
rect 65660 7590 65686 7642
rect 65686 7590 65716 7642
rect 65740 7590 65750 7642
rect 65750 7590 65796 7642
rect 65820 7590 65866 7642
rect 65866 7590 65876 7642
rect 65900 7590 65930 7642
rect 65930 7590 65956 7642
rect 65660 7588 65716 7590
rect 65740 7588 65796 7590
rect 65820 7588 65876 7590
rect 65900 7588 65956 7590
rect 65430 6740 65432 6760
rect 65432 6740 65484 6760
rect 65484 6740 65486 6760
rect 65430 6704 65486 6740
rect 65522 6604 65524 6624
rect 65524 6604 65576 6624
rect 65576 6604 65578 6624
rect 65522 6568 65578 6604
rect 65660 6554 65716 6556
rect 65740 6554 65796 6556
rect 65820 6554 65876 6556
rect 65900 6554 65956 6556
rect 65660 6502 65686 6554
rect 65686 6502 65716 6554
rect 65740 6502 65750 6554
rect 65750 6502 65796 6554
rect 65820 6502 65866 6554
rect 65866 6502 65876 6554
rect 65900 6502 65930 6554
rect 65930 6502 65956 6554
rect 65660 6500 65716 6502
rect 65740 6500 65796 6502
rect 65820 6500 65876 6502
rect 65900 6500 65956 6502
rect 65982 6024 66038 6080
rect 65798 5616 65854 5672
rect 65522 5480 65578 5536
rect 65660 5466 65716 5468
rect 65740 5466 65796 5468
rect 65820 5466 65876 5468
rect 65900 5466 65956 5468
rect 65660 5414 65686 5466
rect 65686 5414 65716 5466
rect 65740 5414 65750 5466
rect 65750 5414 65796 5466
rect 65820 5414 65866 5466
rect 65866 5414 65876 5466
rect 65900 5414 65930 5466
rect 65930 5414 65956 5466
rect 65660 5412 65716 5414
rect 65740 5412 65796 5414
rect 65820 5412 65876 5414
rect 65900 5412 65956 5414
rect 65660 4378 65716 4380
rect 65740 4378 65796 4380
rect 65820 4378 65876 4380
rect 65900 4378 65956 4380
rect 65660 4326 65686 4378
rect 65686 4326 65716 4378
rect 65740 4326 65750 4378
rect 65750 4326 65796 4378
rect 65820 4326 65866 4378
rect 65866 4326 65876 4378
rect 65900 4326 65930 4378
rect 65930 4326 65956 4378
rect 65660 4324 65716 4326
rect 65740 4324 65796 4326
rect 65820 4324 65876 4326
rect 65900 4324 65956 4326
rect 65660 3290 65716 3292
rect 65740 3290 65796 3292
rect 65820 3290 65876 3292
rect 65900 3290 65956 3292
rect 65660 3238 65686 3290
rect 65686 3238 65716 3290
rect 65740 3238 65750 3290
rect 65750 3238 65796 3290
rect 65820 3238 65866 3290
rect 65866 3238 65876 3290
rect 65900 3238 65930 3290
rect 65930 3238 65956 3290
rect 65660 3236 65716 3238
rect 65740 3236 65796 3238
rect 65820 3236 65876 3238
rect 65900 3236 65956 3238
rect 65660 2202 65716 2204
rect 65740 2202 65796 2204
rect 65820 2202 65876 2204
rect 65900 2202 65956 2204
rect 65660 2150 65686 2202
rect 65686 2150 65716 2202
rect 65740 2150 65750 2202
rect 65750 2150 65796 2202
rect 65820 2150 65866 2202
rect 65866 2150 65876 2202
rect 65900 2150 65930 2202
rect 65930 2150 65956 2202
rect 65660 2148 65716 2150
rect 65740 2148 65796 2150
rect 65820 2148 65876 2150
rect 65900 2148 65956 2150
rect 66258 6976 66314 7032
rect 66902 6296 66958 6352
rect 68282 3712 68338 3768
rect 68558 3304 68614 3360
rect 68650 2916 68706 2952
rect 68650 2896 68652 2916
rect 68652 2896 68704 2916
rect 68704 2896 68706 2916
rect 81020 116986 81076 116988
rect 81100 116986 81156 116988
rect 81180 116986 81236 116988
rect 81260 116986 81316 116988
rect 81020 116934 81046 116986
rect 81046 116934 81076 116986
rect 81100 116934 81110 116986
rect 81110 116934 81156 116986
rect 81180 116934 81226 116986
rect 81226 116934 81236 116986
rect 81260 116934 81290 116986
rect 81290 116934 81316 116986
rect 81020 116932 81076 116934
rect 81100 116932 81156 116934
rect 81180 116932 81236 116934
rect 81260 116932 81316 116934
rect 96380 116442 96436 116444
rect 96460 116442 96516 116444
rect 96540 116442 96596 116444
rect 96620 116442 96676 116444
rect 96380 116390 96406 116442
rect 96406 116390 96436 116442
rect 96460 116390 96470 116442
rect 96470 116390 96516 116442
rect 96540 116390 96586 116442
rect 96586 116390 96596 116442
rect 96620 116390 96650 116442
rect 96650 116390 96676 116442
rect 96380 116388 96436 116390
rect 96460 116388 96516 116390
rect 96540 116388 96596 116390
rect 96620 116388 96676 116390
rect 111740 116986 111796 116988
rect 111820 116986 111876 116988
rect 111900 116986 111956 116988
rect 111980 116986 112036 116988
rect 111740 116934 111766 116986
rect 111766 116934 111796 116986
rect 111820 116934 111830 116986
rect 111830 116934 111876 116986
rect 111900 116934 111946 116986
rect 111946 116934 111956 116986
rect 111980 116934 112010 116986
rect 112010 116934 112036 116986
rect 111740 116932 111796 116934
rect 111820 116932 111876 116934
rect 111900 116932 111956 116934
rect 111980 116932 112036 116934
rect 81020 115898 81076 115900
rect 81100 115898 81156 115900
rect 81180 115898 81236 115900
rect 81260 115898 81316 115900
rect 81020 115846 81046 115898
rect 81046 115846 81076 115898
rect 81100 115846 81110 115898
rect 81110 115846 81156 115898
rect 81180 115846 81226 115898
rect 81226 115846 81236 115898
rect 81260 115846 81290 115898
rect 81290 115846 81316 115898
rect 81020 115844 81076 115846
rect 81100 115844 81156 115846
rect 81180 115844 81236 115846
rect 81260 115844 81316 115846
rect 111740 115898 111796 115900
rect 111820 115898 111876 115900
rect 111900 115898 111956 115900
rect 111980 115898 112036 115900
rect 111740 115846 111766 115898
rect 111766 115846 111796 115898
rect 111820 115846 111830 115898
rect 111830 115846 111876 115898
rect 111900 115846 111946 115898
rect 111946 115846 111956 115898
rect 111980 115846 112010 115898
rect 112010 115846 112036 115898
rect 111740 115844 111796 115846
rect 111820 115844 111876 115846
rect 111900 115844 111956 115846
rect 111980 115844 112036 115846
rect 96380 115354 96436 115356
rect 96460 115354 96516 115356
rect 96540 115354 96596 115356
rect 96620 115354 96676 115356
rect 96380 115302 96406 115354
rect 96406 115302 96436 115354
rect 96460 115302 96470 115354
rect 96470 115302 96516 115354
rect 96540 115302 96586 115354
rect 96586 115302 96596 115354
rect 96620 115302 96650 115354
rect 96650 115302 96676 115354
rect 96380 115300 96436 115302
rect 96460 115300 96516 115302
rect 96540 115300 96596 115302
rect 96620 115300 96676 115302
rect 81020 114810 81076 114812
rect 81100 114810 81156 114812
rect 81180 114810 81236 114812
rect 81260 114810 81316 114812
rect 81020 114758 81046 114810
rect 81046 114758 81076 114810
rect 81100 114758 81110 114810
rect 81110 114758 81156 114810
rect 81180 114758 81226 114810
rect 81226 114758 81236 114810
rect 81260 114758 81290 114810
rect 81290 114758 81316 114810
rect 81020 114756 81076 114758
rect 81100 114756 81156 114758
rect 81180 114756 81236 114758
rect 81260 114756 81316 114758
rect 111740 114810 111796 114812
rect 111820 114810 111876 114812
rect 111900 114810 111956 114812
rect 111980 114810 112036 114812
rect 111740 114758 111766 114810
rect 111766 114758 111796 114810
rect 111820 114758 111830 114810
rect 111830 114758 111876 114810
rect 111900 114758 111946 114810
rect 111946 114758 111956 114810
rect 111980 114758 112010 114810
rect 112010 114758 112036 114810
rect 111740 114756 111796 114758
rect 111820 114756 111876 114758
rect 111900 114756 111956 114758
rect 111980 114756 112036 114758
rect 96380 114266 96436 114268
rect 96460 114266 96516 114268
rect 96540 114266 96596 114268
rect 96620 114266 96676 114268
rect 96380 114214 96406 114266
rect 96406 114214 96436 114266
rect 96460 114214 96470 114266
rect 96470 114214 96516 114266
rect 96540 114214 96586 114266
rect 96586 114214 96596 114266
rect 96620 114214 96650 114266
rect 96650 114214 96676 114266
rect 96380 114212 96436 114214
rect 96460 114212 96516 114214
rect 96540 114212 96596 114214
rect 96620 114212 96676 114214
rect 81020 113722 81076 113724
rect 81100 113722 81156 113724
rect 81180 113722 81236 113724
rect 81260 113722 81316 113724
rect 81020 113670 81046 113722
rect 81046 113670 81076 113722
rect 81100 113670 81110 113722
rect 81110 113670 81156 113722
rect 81180 113670 81226 113722
rect 81226 113670 81236 113722
rect 81260 113670 81290 113722
rect 81290 113670 81316 113722
rect 81020 113668 81076 113670
rect 81100 113668 81156 113670
rect 81180 113668 81236 113670
rect 81260 113668 81316 113670
rect 111740 113722 111796 113724
rect 111820 113722 111876 113724
rect 111900 113722 111956 113724
rect 111980 113722 112036 113724
rect 111740 113670 111766 113722
rect 111766 113670 111796 113722
rect 111820 113670 111830 113722
rect 111830 113670 111876 113722
rect 111900 113670 111946 113722
rect 111946 113670 111956 113722
rect 111980 113670 112010 113722
rect 112010 113670 112036 113722
rect 111740 113668 111796 113670
rect 111820 113668 111876 113670
rect 111900 113668 111956 113670
rect 111980 113668 112036 113670
rect 96380 113178 96436 113180
rect 96460 113178 96516 113180
rect 96540 113178 96596 113180
rect 96620 113178 96676 113180
rect 96380 113126 96406 113178
rect 96406 113126 96436 113178
rect 96460 113126 96470 113178
rect 96470 113126 96516 113178
rect 96540 113126 96586 113178
rect 96586 113126 96596 113178
rect 96620 113126 96650 113178
rect 96650 113126 96676 113178
rect 96380 113124 96436 113126
rect 96460 113124 96516 113126
rect 96540 113124 96596 113126
rect 96620 113124 96676 113126
rect 81020 112634 81076 112636
rect 81100 112634 81156 112636
rect 81180 112634 81236 112636
rect 81260 112634 81316 112636
rect 81020 112582 81046 112634
rect 81046 112582 81076 112634
rect 81100 112582 81110 112634
rect 81110 112582 81156 112634
rect 81180 112582 81226 112634
rect 81226 112582 81236 112634
rect 81260 112582 81290 112634
rect 81290 112582 81316 112634
rect 81020 112580 81076 112582
rect 81100 112580 81156 112582
rect 81180 112580 81236 112582
rect 81260 112580 81316 112582
rect 111740 112634 111796 112636
rect 111820 112634 111876 112636
rect 111900 112634 111956 112636
rect 111980 112634 112036 112636
rect 111740 112582 111766 112634
rect 111766 112582 111796 112634
rect 111820 112582 111830 112634
rect 111830 112582 111876 112634
rect 111900 112582 111946 112634
rect 111946 112582 111956 112634
rect 111980 112582 112010 112634
rect 112010 112582 112036 112634
rect 111740 112580 111796 112582
rect 111820 112580 111876 112582
rect 111900 112580 111956 112582
rect 111980 112580 112036 112582
rect 96380 112090 96436 112092
rect 96460 112090 96516 112092
rect 96540 112090 96596 112092
rect 96620 112090 96676 112092
rect 96380 112038 96406 112090
rect 96406 112038 96436 112090
rect 96460 112038 96470 112090
rect 96470 112038 96516 112090
rect 96540 112038 96586 112090
rect 96586 112038 96596 112090
rect 96620 112038 96650 112090
rect 96650 112038 96676 112090
rect 96380 112036 96436 112038
rect 96460 112036 96516 112038
rect 96540 112036 96596 112038
rect 96620 112036 96676 112038
rect 81020 111546 81076 111548
rect 81100 111546 81156 111548
rect 81180 111546 81236 111548
rect 81260 111546 81316 111548
rect 81020 111494 81046 111546
rect 81046 111494 81076 111546
rect 81100 111494 81110 111546
rect 81110 111494 81156 111546
rect 81180 111494 81226 111546
rect 81226 111494 81236 111546
rect 81260 111494 81290 111546
rect 81290 111494 81316 111546
rect 81020 111492 81076 111494
rect 81100 111492 81156 111494
rect 81180 111492 81236 111494
rect 81260 111492 81316 111494
rect 111740 111546 111796 111548
rect 111820 111546 111876 111548
rect 111900 111546 111956 111548
rect 111980 111546 112036 111548
rect 111740 111494 111766 111546
rect 111766 111494 111796 111546
rect 111820 111494 111830 111546
rect 111830 111494 111876 111546
rect 111900 111494 111946 111546
rect 111946 111494 111956 111546
rect 111980 111494 112010 111546
rect 112010 111494 112036 111546
rect 111740 111492 111796 111494
rect 111820 111492 111876 111494
rect 111900 111492 111956 111494
rect 111980 111492 112036 111494
rect 96380 111002 96436 111004
rect 96460 111002 96516 111004
rect 96540 111002 96596 111004
rect 96620 111002 96676 111004
rect 96380 110950 96406 111002
rect 96406 110950 96436 111002
rect 96460 110950 96470 111002
rect 96470 110950 96516 111002
rect 96540 110950 96586 111002
rect 96586 110950 96596 111002
rect 96620 110950 96650 111002
rect 96650 110950 96676 111002
rect 96380 110948 96436 110950
rect 96460 110948 96516 110950
rect 96540 110948 96596 110950
rect 96620 110948 96676 110950
rect 81020 110458 81076 110460
rect 81100 110458 81156 110460
rect 81180 110458 81236 110460
rect 81260 110458 81316 110460
rect 81020 110406 81046 110458
rect 81046 110406 81076 110458
rect 81100 110406 81110 110458
rect 81110 110406 81156 110458
rect 81180 110406 81226 110458
rect 81226 110406 81236 110458
rect 81260 110406 81290 110458
rect 81290 110406 81316 110458
rect 81020 110404 81076 110406
rect 81100 110404 81156 110406
rect 81180 110404 81236 110406
rect 81260 110404 81316 110406
rect 111740 110458 111796 110460
rect 111820 110458 111876 110460
rect 111900 110458 111956 110460
rect 111980 110458 112036 110460
rect 111740 110406 111766 110458
rect 111766 110406 111796 110458
rect 111820 110406 111830 110458
rect 111830 110406 111876 110458
rect 111900 110406 111946 110458
rect 111946 110406 111956 110458
rect 111980 110406 112010 110458
rect 112010 110406 112036 110458
rect 111740 110404 111796 110406
rect 111820 110404 111876 110406
rect 111900 110404 111956 110406
rect 111980 110404 112036 110406
rect 96380 109914 96436 109916
rect 96460 109914 96516 109916
rect 96540 109914 96596 109916
rect 96620 109914 96676 109916
rect 96380 109862 96406 109914
rect 96406 109862 96436 109914
rect 96460 109862 96470 109914
rect 96470 109862 96516 109914
rect 96540 109862 96586 109914
rect 96586 109862 96596 109914
rect 96620 109862 96650 109914
rect 96650 109862 96676 109914
rect 96380 109860 96436 109862
rect 96460 109860 96516 109862
rect 96540 109860 96596 109862
rect 96620 109860 96676 109862
rect 81020 109370 81076 109372
rect 81100 109370 81156 109372
rect 81180 109370 81236 109372
rect 81260 109370 81316 109372
rect 81020 109318 81046 109370
rect 81046 109318 81076 109370
rect 81100 109318 81110 109370
rect 81110 109318 81156 109370
rect 81180 109318 81226 109370
rect 81226 109318 81236 109370
rect 81260 109318 81290 109370
rect 81290 109318 81316 109370
rect 81020 109316 81076 109318
rect 81100 109316 81156 109318
rect 81180 109316 81236 109318
rect 81260 109316 81316 109318
rect 111740 109370 111796 109372
rect 111820 109370 111876 109372
rect 111900 109370 111956 109372
rect 111980 109370 112036 109372
rect 111740 109318 111766 109370
rect 111766 109318 111796 109370
rect 111820 109318 111830 109370
rect 111830 109318 111876 109370
rect 111900 109318 111946 109370
rect 111946 109318 111956 109370
rect 111980 109318 112010 109370
rect 112010 109318 112036 109370
rect 111740 109316 111796 109318
rect 111820 109316 111876 109318
rect 111900 109316 111956 109318
rect 111980 109316 112036 109318
rect 96380 108826 96436 108828
rect 96460 108826 96516 108828
rect 96540 108826 96596 108828
rect 96620 108826 96676 108828
rect 96380 108774 96406 108826
rect 96406 108774 96436 108826
rect 96460 108774 96470 108826
rect 96470 108774 96516 108826
rect 96540 108774 96586 108826
rect 96586 108774 96596 108826
rect 96620 108774 96650 108826
rect 96650 108774 96676 108826
rect 96380 108772 96436 108774
rect 96460 108772 96516 108774
rect 96540 108772 96596 108774
rect 96620 108772 96676 108774
rect 81020 108282 81076 108284
rect 81100 108282 81156 108284
rect 81180 108282 81236 108284
rect 81260 108282 81316 108284
rect 81020 108230 81046 108282
rect 81046 108230 81076 108282
rect 81100 108230 81110 108282
rect 81110 108230 81156 108282
rect 81180 108230 81226 108282
rect 81226 108230 81236 108282
rect 81260 108230 81290 108282
rect 81290 108230 81316 108282
rect 81020 108228 81076 108230
rect 81100 108228 81156 108230
rect 81180 108228 81236 108230
rect 81260 108228 81316 108230
rect 111740 108282 111796 108284
rect 111820 108282 111876 108284
rect 111900 108282 111956 108284
rect 111980 108282 112036 108284
rect 111740 108230 111766 108282
rect 111766 108230 111796 108282
rect 111820 108230 111830 108282
rect 111830 108230 111876 108282
rect 111900 108230 111946 108282
rect 111946 108230 111956 108282
rect 111980 108230 112010 108282
rect 112010 108230 112036 108282
rect 111740 108228 111796 108230
rect 111820 108228 111876 108230
rect 111900 108228 111956 108230
rect 111980 108228 112036 108230
rect 96380 107738 96436 107740
rect 96460 107738 96516 107740
rect 96540 107738 96596 107740
rect 96620 107738 96676 107740
rect 96380 107686 96406 107738
rect 96406 107686 96436 107738
rect 96460 107686 96470 107738
rect 96470 107686 96516 107738
rect 96540 107686 96586 107738
rect 96586 107686 96596 107738
rect 96620 107686 96650 107738
rect 96650 107686 96676 107738
rect 96380 107684 96436 107686
rect 96460 107684 96516 107686
rect 96540 107684 96596 107686
rect 96620 107684 96676 107686
rect 81020 107194 81076 107196
rect 81100 107194 81156 107196
rect 81180 107194 81236 107196
rect 81260 107194 81316 107196
rect 81020 107142 81046 107194
rect 81046 107142 81076 107194
rect 81100 107142 81110 107194
rect 81110 107142 81156 107194
rect 81180 107142 81226 107194
rect 81226 107142 81236 107194
rect 81260 107142 81290 107194
rect 81290 107142 81316 107194
rect 81020 107140 81076 107142
rect 81100 107140 81156 107142
rect 81180 107140 81236 107142
rect 81260 107140 81316 107142
rect 111740 107194 111796 107196
rect 111820 107194 111876 107196
rect 111900 107194 111956 107196
rect 111980 107194 112036 107196
rect 111740 107142 111766 107194
rect 111766 107142 111796 107194
rect 111820 107142 111830 107194
rect 111830 107142 111876 107194
rect 111900 107142 111946 107194
rect 111946 107142 111956 107194
rect 111980 107142 112010 107194
rect 112010 107142 112036 107194
rect 111740 107140 111796 107142
rect 111820 107140 111876 107142
rect 111900 107140 111956 107142
rect 111980 107140 112036 107142
rect 96380 106650 96436 106652
rect 96460 106650 96516 106652
rect 96540 106650 96596 106652
rect 96620 106650 96676 106652
rect 96380 106598 96406 106650
rect 96406 106598 96436 106650
rect 96460 106598 96470 106650
rect 96470 106598 96516 106650
rect 96540 106598 96586 106650
rect 96586 106598 96596 106650
rect 96620 106598 96650 106650
rect 96650 106598 96676 106650
rect 96380 106596 96436 106598
rect 96460 106596 96516 106598
rect 96540 106596 96596 106598
rect 96620 106596 96676 106598
rect 81020 106106 81076 106108
rect 81100 106106 81156 106108
rect 81180 106106 81236 106108
rect 81260 106106 81316 106108
rect 81020 106054 81046 106106
rect 81046 106054 81076 106106
rect 81100 106054 81110 106106
rect 81110 106054 81156 106106
rect 81180 106054 81226 106106
rect 81226 106054 81236 106106
rect 81260 106054 81290 106106
rect 81290 106054 81316 106106
rect 81020 106052 81076 106054
rect 81100 106052 81156 106054
rect 81180 106052 81236 106054
rect 81260 106052 81316 106054
rect 111740 106106 111796 106108
rect 111820 106106 111876 106108
rect 111900 106106 111956 106108
rect 111980 106106 112036 106108
rect 111740 106054 111766 106106
rect 111766 106054 111796 106106
rect 111820 106054 111830 106106
rect 111830 106054 111876 106106
rect 111900 106054 111946 106106
rect 111946 106054 111956 106106
rect 111980 106054 112010 106106
rect 112010 106054 112036 106106
rect 111740 106052 111796 106054
rect 111820 106052 111876 106054
rect 111900 106052 111956 106054
rect 111980 106052 112036 106054
rect 96380 105562 96436 105564
rect 96460 105562 96516 105564
rect 96540 105562 96596 105564
rect 96620 105562 96676 105564
rect 96380 105510 96406 105562
rect 96406 105510 96436 105562
rect 96460 105510 96470 105562
rect 96470 105510 96516 105562
rect 96540 105510 96586 105562
rect 96586 105510 96596 105562
rect 96620 105510 96650 105562
rect 96650 105510 96676 105562
rect 96380 105508 96436 105510
rect 96460 105508 96516 105510
rect 96540 105508 96596 105510
rect 96620 105508 96676 105510
rect 81020 105018 81076 105020
rect 81100 105018 81156 105020
rect 81180 105018 81236 105020
rect 81260 105018 81316 105020
rect 81020 104966 81046 105018
rect 81046 104966 81076 105018
rect 81100 104966 81110 105018
rect 81110 104966 81156 105018
rect 81180 104966 81226 105018
rect 81226 104966 81236 105018
rect 81260 104966 81290 105018
rect 81290 104966 81316 105018
rect 81020 104964 81076 104966
rect 81100 104964 81156 104966
rect 81180 104964 81236 104966
rect 81260 104964 81316 104966
rect 111740 105018 111796 105020
rect 111820 105018 111876 105020
rect 111900 105018 111956 105020
rect 111980 105018 112036 105020
rect 111740 104966 111766 105018
rect 111766 104966 111796 105018
rect 111820 104966 111830 105018
rect 111830 104966 111876 105018
rect 111900 104966 111946 105018
rect 111946 104966 111956 105018
rect 111980 104966 112010 105018
rect 112010 104966 112036 105018
rect 111740 104964 111796 104966
rect 111820 104964 111876 104966
rect 111900 104964 111956 104966
rect 111980 104964 112036 104966
rect 96380 104474 96436 104476
rect 96460 104474 96516 104476
rect 96540 104474 96596 104476
rect 96620 104474 96676 104476
rect 96380 104422 96406 104474
rect 96406 104422 96436 104474
rect 96460 104422 96470 104474
rect 96470 104422 96516 104474
rect 96540 104422 96586 104474
rect 96586 104422 96596 104474
rect 96620 104422 96650 104474
rect 96650 104422 96676 104474
rect 96380 104420 96436 104422
rect 96460 104420 96516 104422
rect 96540 104420 96596 104422
rect 96620 104420 96676 104422
rect 81020 103930 81076 103932
rect 81100 103930 81156 103932
rect 81180 103930 81236 103932
rect 81260 103930 81316 103932
rect 81020 103878 81046 103930
rect 81046 103878 81076 103930
rect 81100 103878 81110 103930
rect 81110 103878 81156 103930
rect 81180 103878 81226 103930
rect 81226 103878 81236 103930
rect 81260 103878 81290 103930
rect 81290 103878 81316 103930
rect 81020 103876 81076 103878
rect 81100 103876 81156 103878
rect 81180 103876 81236 103878
rect 81260 103876 81316 103878
rect 111740 103930 111796 103932
rect 111820 103930 111876 103932
rect 111900 103930 111956 103932
rect 111980 103930 112036 103932
rect 111740 103878 111766 103930
rect 111766 103878 111796 103930
rect 111820 103878 111830 103930
rect 111830 103878 111876 103930
rect 111900 103878 111946 103930
rect 111946 103878 111956 103930
rect 111980 103878 112010 103930
rect 112010 103878 112036 103930
rect 111740 103876 111796 103878
rect 111820 103876 111876 103878
rect 111900 103876 111956 103878
rect 111980 103876 112036 103878
rect 96380 103386 96436 103388
rect 96460 103386 96516 103388
rect 96540 103386 96596 103388
rect 96620 103386 96676 103388
rect 96380 103334 96406 103386
rect 96406 103334 96436 103386
rect 96460 103334 96470 103386
rect 96470 103334 96516 103386
rect 96540 103334 96586 103386
rect 96586 103334 96596 103386
rect 96620 103334 96650 103386
rect 96650 103334 96676 103386
rect 96380 103332 96436 103334
rect 96460 103332 96516 103334
rect 96540 103332 96596 103334
rect 96620 103332 96676 103334
rect 81020 102842 81076 102844
rect 81100 102842 81156 102844
rect 81180 102842 81236 102844
rect 81260 102842 81316 102844
rect 81020 102790 81046 102842
rect 81046 102790 81076 102842
rect 81100 102790 81110 102842
rect 81110 102790 81156 102842
rect 81180 102790 81226 102842
rect 81226 102790 81236 102842
rect 81260 102790 81290 102842
rect 81290 102790 81316 102842
rect 81020 102788 81076 102790
rect 81100 102788 81156 102790
rect 81180 102788 81236 102790
rect 81260 102788 81316 102790
rect 111740 102842 111796 102844
rect 111820 102842 111876 102844
rect 111900 102842 111956 102844
rect 111980 102842 112036 102844
rect 111740 102790 111766 102842
rect 111766 102790 111796 102842
rect 111820 102790 111830 102842
rect 111830 102790 111876 102842
rect 111900 102790 111946 102842
rect 111946 102790 111956 102842
rect 111980 102790 112010 102842
rect 112010 102790 112036 102842
rect 111740 102788 111796 102790
rect 111820 102788 111876 102790
rect 111900 102788 111956 102790
rect 111980 102788 112036 102790
rect 96380 102298 96436 102300
rect 96460 102298 96516 102300
rect 96540 102298 96596 102300
rect 96620 102298 96676 102300
rect 96380 102246 96406 102298
rect 96406 102246 96436 102298
rect 96460 102246 96470 102298
rect 96470 102246 96516 102298
rect 96540 102246 96586 102298
rect 96586 102246 96596 102298
rect 96620 102246 96650 102298
rect 96650 102246 96676 102298
rect 96380 102244 96436 102246
rect 96460 102244 96516 102246
rect 96540 102244 96596 102246
rect 96620 102244 96676 102246
rect 81020 101754 81076 101756
rect 81100 101754 81156 101756
rect 81180 101754 81236 101756
rect 81260 101754 81316 101756
rect 81020 101702 81046 101754
rect 81046 101702 81076 101754
rect 81100 101702 81110 101754
rect 81110 101702 81156 101754
rect 81180 101702 81226 101754
rect 81226 101702 81236 101754
rect 81260 101702 81290 101754
rect 81290 101702 81316 101754
rect 81020 101700 81076 101702
rect 81100 101700 81156 101702
rect 81180 101700 81236 101702
rect 81260 101700 81316 101702
rect 111740 101754 111796 101756
rect 111820 101754 111876 101756
rect 111900 101754 111956 101756
rect 111980 101754 112036 101756
rect 111740 101702 111766 101754
rect 111766 101702 111796 101754
rect 111820 101702 111830 101754
rect 111830 101702 111876 101754
rect 111900 101702 111946 101754
rect 111946 101702 111956 101754
rect 111980 101702 112010 101754
rect 112010 101702 112036 101754
rect 111740 101700 111796 101702
rect 111820 101700 111876 101702
rect 111900 101700 111956 101702
rect 111980 101700 112036 101702
rect 96380 101210 96436 101212
rect 96460 101210 96516 101212
rect 96540 101210 96596 101212
rect 96620 101210 96676 101212
rect 96380 101158 96406 101210
rect 96406 101158 96436 101210
rect 96460 101158 96470 101210
rect 96470 101158 96516 101210
rect 96540 101158 96586 101210
rect 96586 101158 96596 101210
rect 96620 101158 96650 101210
rect 96650 101158 96676 101210
rect 96380 101156 96436 101158
rect 96460 101156 96516 101158
rect 96540 101156 96596 101158
rect 96620 101156 96676 101158
rect 81020 100666 81076 100668
rect 81100 100666 81156 100668
rect 81180 100666 81236 100668
rect 81260 100666 81316 100668
rect 81020 100614 81046 100666
rect 81046 100614 81076 100666
rect 81100 100614 81110 100666
rect 81110 100614 81156 100666
rect 81180 100614 81226 100666
rect 81226 100614 81236 100666
rect 81260 100614 81290 100666
rect 81290 100614 81316 100666
rect 81020 100612 81076 100614
rect 81100 100612 81156 100614
rect 81180 100612 81236 100614
rect 81260 100612 81316 100614
rect 111740 100666 111796 100668
rect 111820 100666 111876 100668
rect 111900 100666 111956 100668
rect 111980 100666 112036 100668
rect 111740 100614 111766 100666
rect 111766 100614 111796 100666
rect 111820 100614 111830 100666
rect 111830 100614 111876 100666
rect 111900 100614 111946 100666
rect 111946 100614 111956 100666
rect 111980 100614 112010 100666
rect 112010 100614 112036 100666
rect 111740 100612 111796 100614
rect 111820 100612 111876 100614
rect 111900 100612 111956 100614
rect 111980 100612 112036 100614
rect 96380 100122 96436 100124
rect 96460 100122 96516 100124
rect 96540 100122 96596 100124
rect 96620 100122 96676 100124
rect 96380 100070 96406 100122
rect 96406 100070 96436 100122
rect 96460 100070 96470 100122
rect 96470 100070 96516 100122
rect 96540 100070 96586 100122
rect 96586 100070 96596 100122
rect 96620 100070 96650 100122
rect 96650 100070 96676 100122
rect 96380 100068 96436 100070
rect 96460 100068 96516 100070
rect 96540 100068 96596 100070
rect 96620 100068 96676 100070
rect 81020 99578 81076 99580
rect 81100 99578 81156 99580
rect 81180 99578 81236 99580
rect 81260 99578 81316 99580
rect 81020 99526 81046 99578
rect 81046 99526 81076 99578
rect 81100 99526 81110 99578
rect 81110 99526 81156 99578
rect 81180 99526 81226 99578
rect 81226 99526 81236 99578
rect 81260 99526 81290 99578
rect 81290 99526 81316 99578
rect 81020 99524 81076 99526
rect 81100 99524 81156 99526
rect 81180 99524 81236 99526
rect 81260 99524 81316 99526
rect 111740 99578 111796 99580
rect 111820 99578 111876 99580
rect 111900 99578 111956 99580
rect 111980 99578 112036 99580
rect 111740 99526 111766 99578
rect 111766 99526 111796 99578
rect 111820 99526 111830 99578
rect 111830 99526 111876 99578
rect 111900 99526 111946 99578
rect 111946 99526 111956 99578
rect 111980 99526 112010 99578
rect 112010 99526 112036 99578
rect 111740 99524 111796 99526
rect 111820 99524 111876 99526
rect 111900 99524 111956 99526
rect 111980 99524 112036 99526
rect 96380 99034 96436 99036
rect 96460 99034 96516 99036
rect 96540 99034 96596 99036
rect 96620 99034 96676 99036
rect 96380 98982 96406 99034
rect 96406 98982 96436 99034
rect 96460 98982 96470 99034
rect 96470 98982 96516 99034
rect 96540 98982 96586 99034
rect 96586 98982 96596 99034
rect 96620 98982 96650 99034
rect 96650 98982 96676 99034
rect 96380 98980 96436 98982
rect 96460 98980 96516 98982
rect 96540 98980 96596 98982
rect 96620 98980 96676 98982
rect 81020 98490 81076 98492
rect 81100 98490 81156 98492
rect 81180 98490 81236 98492
rect 81260 98490 81316 98492
rect 81020 98438 81046 98490
rect 81046 98438 81076 98490
rect 81100 98438 81110 98490
rect 81110 98438 81156 98490
rect 81180 98438 81226 98490
rect 81226 98438 81236 98490
rect 81260 98438 81290 98490
rect 81290 98438 81316 98490
rect 81020 98436 81076 98438
rect 81100 98436 81156 98438
rect 81180 98436 81236 98438
rect 81260 98436 81316 98438
rect 111740 98490 111796 98492
rect 111820 98490 111876 98492
rect 111900 98490 111956 98492
rect 111980 98490 112036 98492
rect 111740 98438 111766 98490
rect 111766 98438 111796 98490
rect 111820 98438 111830 98490
rect 111830 98438 111876 98490
rect 111900 98438 111946 98490
rect 111946 98438 111956 98490
rect 111980 98438 112010 98490
rect 112010 98438 112036 98490
rect 111740 98436 111796 98438
rect 111820 98436 111876 98438
rect 111900 98436 111956 98438
rect 111980 98436 112036 98438
rect 96380 97946 96436 97948
rect 96460 97946 96516 97948
rect 96540 97946 96596 97948
rect 96620 97946 96676 97948
rect 96380 97894 96406 97946
rect 96406 97894 96436 97946
rect 96460 97894 96470 97946
rect 96470 97894 96516 97946
rect 96540 97894 96586 97946
rect 96586 97894 96596 97946
rect 96620 97894 96650 97946
rect 96650 97894 96676 97946
rect 96380 97892 96436 97894
rect 96460 97892 96516 97894
rect 96540 97892 96596 97894
rect 96620 97892 96676 97894
rect 81020 97402 81076 97404
rect 81100 97402 81156 97404
rect 81180 97402 81236 97404
rect 81260 97402 81316 97404
rect 81020 97350 81046 97402
rect 81046 97350 81076 97402
rect 81100 97350 81110 97402
rect 81110 97350 81156 97402
rect 81180 97350 81226 97402
rect 81226 97350 81236 97402
rect 81260 97350 81290 97402
rect 81290 97350 81316 97402
rect 81020 97348 81076 97350
rect 81100 97348 81156 97350
rect 81180 97348 81236 97350
rect 81260 97348 81316 97350
rect 111740 97402 111796 97404
rect 111820 97402 111876 97404
rect 111900 97402 111956 97404
rect 111980 97402 112036 97404
rect 111740 97350 111766 97402
rect 111766 97350 111796 97402
rect 111820 97350 111830 97402
rect 111830 97350 111876 97402
rect 111900 97350 111946 97402
rect 111946 97350 111956 97402
rect 111980 97350 112010 97402
rect 112010 97350 112036 97402
rect 111740 97348 111796 97350
rect 111820 97348 111876 97350
rect 111900 97348 111956 97350
rect 111980 97348 112036 97350
rect 96380 96858 96436 96860
rect 96460 96858 96516 96860
rect 96540 96858 96596 96860
rect 96620 96858 96676 96860
rect 96380 96806 96406 96858
rect 96406 96806 96436 96858
rect 96460 96806 96470 96858
rect 96470 96806 96516 96858
rect 96540 96806 96586 96858
rect 96586 96806 96596 96858
rect 96620 96806 96650 96858
rect 96650 96806 96676 96858
rect 96380 96804 96436 96806
rect 96460 96804 96516 96806
rect 96540 96804 96596 96806
rect 96620 96804 96676 96806
rect 81020 96314 81076 96316
rect 81100 96314 81156 96316
rect 81180 96314 81236 96316
rect 81260 96314 81316 96316
rect 81020 96262 81046 96314
rect 81046 96262 81076 96314
rect 81100 96262 81110 96314
rect 81110 96262 81156 96314
rect 81180 96262 81226 96314
rect 81226 96262 81236 96314
rect 81260 96262 81290 96314
rect 81290 96262 81316 96314
rect 81020 96260 81076 96262
rect 81100 96260 81156 96262
rect 81180 96260 81236 96262
rect 81260 96260 81316 96262
rect 111740 96314 111796 96316
rect 111820 96314 111876 96316
rect 111900 96314 111956 96316
rect 111980 96314 112036 96316
rect 111740 96262 111766 96314
rect 111766 96262 111796 96314
rect 111820 96262 111830 96314
rect 111830 96262 111876 96314
rect 111900 96262 111946 96314
rect 111946 96262 111956 96314
rect 111980 96262 112010 96314
rect 112010 96262 112036 96314
rect 111740 96260 111796 96262
rect 111820 96260 111876 96262
rect 111900 96260 111956 96262
rect 111980 96260 112036 96262
rect 96380 95770 96436 95772
rect 96460 95770 96516 95772
rect 96540 95770 96596 95772
rect 96620 95770 96676 95772
rect 96380 95718 96406 95770
rect 96406 95718 96436 95770
rect 96460 95718 96470 95770
rect 96470 95718 96516 95770
rect 96540 95718 96586 95770
rect 96586 95718 96596 95770
rect 96620 95718 96650 95770
rect 96650 95718 96676 95770
rect 96380 95716 96436 95718
rect 96460 95716 96516 95718
rect 96540 95716 96596 95718
rect 96620 95716 96676 95718
rect 81020 95226 81076 95228
rect 81100 95226 81156 95228
rect 81180 95226 81236 95228
rect 81260 95226 81316 95228
rect 81020 95174 81046 95226
rect 81046 95174 81076 95226
rect 81100 95174 81110 95226
rect 81110 95174 81156 95226
rect 81180 95174 81226 95226
rect 81226 95174 81236 95226
rect 81260 95174 81290 95226
rect 81290 95174 81316 95226
rect 81020 95172 81076 95174
rect 81100 95172 81156 95174
rect 81180 95172 81236 95174
rect 81260 95172 81316 95174
rect 111740 95226 111796 95228
rect 111820 95226 111876 95228
rect 111900 95226 111956 95228
rect 111980 95226 112036 95228
rect 111740 95174 111766 95226
rect 111766 95174 111796 95226
rect 111820 95174 111830 95226
rect 111830 95174 111876 95226
rect 111900 95174 111946 95226
rect 111946 95174 111956 95226
rect 111980 95174 112010 95226
rect 112010 95174 112036 95226
rect 111740 95172 111796 95174
rect 111820 95172 111876 95174
rect 111900 95172 111956 95174
rect 111980 95172 112036 95174
rect 96380 94682 96436 94684
rect 96460 94682 96516 94684
rect 96540 94682 96596 94684
rect 96620 94682 96676 94684
rect 96380 94630 96406 94682
rect 96406 94630 96436 94682
rect 96460 94630 96470 94682
rect 96470 94630 96516 94682
rect 96540 94630 96586 94682
rect 96586 94630 96596 94682
rect 96620 94630 96650 94682
rect 96650 94630 96676 94682
rect 96380 94628 96436 94630
rect 96460 94628 96516 94630
rect 96540 94628 96596 94630
rect 96620 94628 96676 94630
rect 81020 94138 81076 94140
rect 81100 94138 81156 94140
rect 81180 94138 81236 94140
rect 81260 94138 81316 94140
rect 81020 94086 81046 94138
rect 81046 94086 81076 94138
rect 81100 94086 81110 94138
rect 81110 94086 81156 94138
rect 81180 94086 81226 94138
rect 81226 94086 81236 94138
rect 81260 94086 81290 94138
rect 81290 94086 81316 94138
rect 81020 94084 81076 94086
rect 81100 94084 81156 94086
rect 81180 94084 81236 94086
rect 81260 94084 81316 94086
rect 111740 94138 111796 94140
rect 111820 94138 111876 94140
rect 111900 94138 111956 94140
rect 111980 94138 112036 94140
rect 111740 94086 111766 94138
rect 111766 94086 111796 94138
rect 111820 94086 111830 94138
rect 111830 94086 111876 94138
rect 111900 94086 111946 94138
rect 111946 94086 111956 94138
rect 111980 94086 112010 94138
rect 112010 94086 112036 94138
rect 111740 94084 111796 94086
rect 111820 94084 111876 94086
rect 111900 94084 111956 94086
rect 111980 94084 112036 94086
rect 96380 93594 96436 93596
rect 96460 93594 96516 93596
rect 96540 93594 96596 93596
rect 96620 93594 96676 93596
rect 96380 93542 96406 93594
rect 96406 93542 96436 93594
rect 96460 93542 96470 93594
rect 96470 93542 96516 93594
rect 96540 93542 96586 93594
rect 96586 93542 96596 93594
rect 96620 93542 96650 93594
rect 96650 93542 96676 93594
rect 96380 93540 96436 93542
rect 96460 93540 96516 93542
rect 96540 93540 96596 93542
rect 96620 93540 96676 93542
rect 81020 93050 81076 93052
rect 81100 93050 81156 93052
rect 81180 93050 81236 93052
rect 81260 93050 81316 93052
rect 81020 92998 81046 93050
rect 81046 92998 81076 93050
rect 81100 92998 81110 93050
rect 81110 92998 81156 93050
rect 81180 92998 81226 93050
rect 81226 92998 81236 93050
rect 81260 92998 81290 93050
rect 81290 92998 81316 93050
rect 81020 92996 81076 92998
rect 81100 92996 81156 92998
rect 81180 92996 81236 92998
rect 81260 92996 81316 92998
rect 111740 93050 111796 93052
rect 111820 93050 111876 93052
rect 111900 93050 111956 93052
rect 111980 93050 112036 93052
rect 111740 92998 111766 93050
rect 111766 92998 111796 93050
rect 111820 92998 111830 93050
rect 111830 92998 111876 93050
rect 111900 92998 111946 93050
rect 111946 92998 111956 93050
rect 111980 92998 112010 93050
rect 112010 92998 112036 93050
rect 111740 92996 111796 92998
rect 111820 92996 111876 92998
rect 111900 92996 111956 92998
rect 111980 92996 112036 92998
rect 96380 92506 96436 92508
rect 96460 92506 96516 92508
rect 96540 92506 96596 92508
rect 96620 92506 96676 92508
rect 96380 92454 96406 92506
rect 96406 92454 96436 92506
rect 96460 92454 96470 92506
rect 96470 92454 96516 92506
rect 96540 92454 96586 92506
rect 96586 92454 96596 92506
rect 96620 92454 96650 92506
rect 96650 92454 96676 92506
rect 96380 92452 96436 92454
rect 96460 92452 96516 92454
rect 96540 92452 96596 92454
rect 96620 92452 96676 92454
rect 81020 91962 81076 91964
rect 81100 91962 81156 91964
rect 81180 91962 81236 91964
rect 81260 91962 81316 91964
rect 81020 91910 81046 91962
rect 81046 91910 81076 91962
rect 81100 91910 81110 91962
rect 81110 91910 81156 91962
rect 81180 91910 81226 91962
rect 81226 91910 81236 91962
rect 81260 91910 81290 91962
rect 81290 91910 81316 91962
rect 81020 91908 81076 91910
rect 81100 91908 81156 91910
rect 81180 91908 81236 91910
rect 81260 91908 81316 91910
rect 111740 91962 111796 91964
rect 111820 91962 111876 91964
rect 111900 91962 111956 91964
rect 111980 91962 112036 91964
rect 111740 91910 111766 91962
rect 111766 91910 111796 91962
rect 111820 91910 111830 91962
rect 111830 91910 111876 91962
rect 111900 91910 111946 91962
rect 111946 91910 111956 91962
rect 111980 91910 112010 91962
rect 112010 91910 112036 91962
rect 111740 91908 111796 91910
rect 111820 91908 111876 91910
rect 111900 91908 111956 91910
rect 111980 91908 112036 91910
rect 96380 91418 96436 91420
rect 96460 91418 96516 91420
rect 96540 91418 96596 91420
rect 96620 91418 96676 91420
rect 96380 91366 96406 91418
rect 96406 91366 96436 91418
rect 96460 91366 96470 91418
rect 96470 91366 96516 91418
rect 96540 91366 96586 91418
rect 96586 91366 96596 91418
rect 96620 91366 96650 91418
rect 96650 91366 96676 91418
rect 96380 91364 96436 91366
rect 96460 91364 96516 91366
rect 96540 91364 96596 91366
rect 96620 91364 96676 91366
rect 81020 90874 81076 90876
rect 81100 90874 81156 90876
rect 81180 90874 81236 90876
rect 81260 90874 81316 90876
rect 81020 90822 81046 90874
rect 81046 90822 81076 90874
rect 81100 90822 81110 90874
rect 81110 90822 81156 90874
rect 81180 90822 81226 90874
rect 81226 90822 81236 90874
rect 81260 90822 81290 90874
rect 81290 90822 81316 90874
rect 81020 90820 81076 90822
rect 81100 90820 81156 90822
rect 81180 90820 81236 90822
rect 81260 90820 81316 90822
rect 111740 90874 111796 90876
rect 111820 90874 111876 90876
rect 111900 90874 111956 90876
rect 111980 90874 112036 90876
rect 111740 90822 111766 90874
rect 111766 90822 111796 90874
rect 111820 90822 111830 90874
rect 111830 90822 111876 90874
rect 111900 90822 111946 90874
rect 111946 90822 111956 90874
rect 111980 90822 112010 90874
rect 112010 90822 112036 90874
rect 111740 90820 111796 90822
rect 111820 90820 111876 90822
rect 111900 90820 111956 90822
rect 111980 90820 112036 90822
rect 96380 90330 96436 90332
rect 96460 90330 96516 90332
rect 96540 90330 96596 90332
rect 96620 90330 96676 90332
rect 96380 90278 96406 90330
rect 96406 90278 96436 90330
rect 96460 90278 96470 90330
rect 96470 90278 96516 90330
rect 96540 90278 96586 90330
rect 96586 90278 96596 90330
rect 96620 90278 96650 90330
rect 96650 90278 96676 90330
rect 96380 90276 96436 90278
rect 96460 90276 96516 90278
rect 96540 90276 96596 90278
rect 96620 90276 96676 90278
rect 81020 89786 81076 89788
rect 81100 89786 81156 89788
rect 81180 89786 81236 89788
rect 81260 89786 81316 89788
rect 81020 89734 81046 89786
rect 81046 89734 81076 89786
rect 81100 89734 81110 89786
rect 81110 89734 81156 89786
rect 81180 89734 81226 89786
rect 81226 89734 81236 89786
rect 81260 89734 81290 89786
rect 81290 89734 81316 89786
rect 81020 89732 81076 89734
rect 81100 89732 81156 89734
rect 81180 89732 81236 89734
rect 81260 89732 81316 89734
rect 111740 89786 111796 89788
rect 111820 89786 111876 89788
rect 111900 89786 111956 89788
rect 111980 89786 112036 89788
rect 111740 89734 111766 89786
rect 111766 89734 111796 89786
rect 111820 89734 111830 89786
rect 111830 89734 111876 89786
rect 111900 89734 111946 89786
rect 111946 89734 111956 89786
rect 111980 89734 112010 89786
rect 112010 89734 112036 89786
rect 111740 89732 111796 89734
rect 111820 89732 111876 89734
rect 111900 89732 111956 89734
rect 111980 89732 112036 89734
rect 96380 89242 96436 89244
rect 96460 89242 96516 89244
rect 96540 89242 96596 89244
rect 96620 89242 96676 89244
rect 96380 89190 96406 89242
rect 96406 89190 96436 89242
rect 96460 89190 96470 89242
rect 96470 89190 96516 89242
rect 96540 89190 96586 89242
rect 96586 89190 96596 89242
rect 96620 89190 96650 89242
rect 96650 89190 96676 89242
rect 96380 89188 96436 89190
rect 96460 89188 96516 89190
rect 96540 89188 96596 89190
rect 96620 89188 96676 89190
rect 81020 88698 81076 88700
rect 81100 88698 81156 88700
rect 81180 88698 81236 88700
rect 81260 88698 81316 88700
rect 81020 88646 81046 88698
rect 81046 88646 81076 88698
rect 81100 88646 81110 88698
rect 81110 88646 81156 88698
rect 81180 88646 81226 88698
rect 81226 88646 81236 88698
rect 81260 88646 81290 88698
rect 81290 88646 81316 88698
rect 81020 88644 81076 88646
rect 81100 88644 81156 88646
rect 81180 88644 81236 88646
rect 81260 88644 81316 88646
rect 111740 88698 111796 88700
rect 111820 88698 111876 88700
rect 111900 88698 111956 88700
rect 111980 88698 112036 88700
rect 111740 88646 111766 88698
rect 111766 88646 111796 88698
rect 111820 88646 111830 88698
rect 111830 88646 111876 88698
rect 111900 88646 111946 88698
rect 111946 88646 111956 88698
rect 111980 88646 112010 88698
rect 112010 88646 112036 88698
rect 111740 88644 111796 88646
rect 111820 88644 111876 88646
rect 111900 88644 111956 88646
rect 111980 88644 112036 88646
rect 96380 88154 96436 88156
rect 96460 88154 96516 88156
rect 96540 88154 96596 88156
rect 96620 88154 96676 88156
rect 96380 88102 96406 88154
rect 96406 88102 96436 88154
rect 96460 88102 96470 88154
rect 96470 88102 96516 88154
rect 96540 88102 96586 88154
rect 96586 88102 96596 88154
rect 96620 88102 96650 88154
rect 96650 88102 96676 88154
rect 96380 88100 96436 88102
rect 96460 88100 96516 88102
rect 96540 88100 96596 88102
rect 96620 88100 96676 88102
rect 81020 87610 81076 87612
rect 81100 87610 81156 87612
rect 81180 87610 81236 87612
rect 81260 87610 81316 87612
rect 81020 87558 81046 87610
rect 81046 87558 81076 87610
rect 81100 87558 81110 87610
rect 81110 87558 81156 87610
rect 81180 87558 81226 87610
rect 81226 87558 81236 87610
rect 81260 87558 81290 87610
rect 81290 87558 81316 87610
rect 81020 87556 81076 87558
rect 81100 87556 81156 87558
rect 81180 87556 81236 87558
rect 81260 87556 81316 87558
rect 111740 87610 111796 87612
rect 111820 87610 111876 87612
rect 111900 87610 111956 87612
rect 111980 87610 112036 87612
rect 111740 87558 111766 87610
rect 111766 87558 111796 87610
rect 111820 87558 111830 87610
rect 111830 87558 111876 87610
rect 111900 87558 111946 87610
rect 111946 87558 111956 87610
rect 111980 87558 112010 87610
rect 112010 87558 112036 87610
rect 111740 87556 111796 87558
rect 111820 87556 111876 87558
rect 111900 87556 111956 87558
rect 111980 87556 112036 87558
rect 96380 87066 96436 87068
rect 96460 87066 96516 87068
rect 96540 87066 96596 87068
rect 96620 87066 96676 87068
rect 96380 87014 96406 87066
rect 96406 87014 96436 87066
rect 96460 87014 96470 87066
rect 96470 87014 96516 87066
rect 96540 87014 96586 87066
rect 96586 87014 96596 87066
rect 96620 87014 96650 87066
rect 96650 87014 96676 87066
rect 96380 87012 96436 87014
rect 96460 87012 96516 87014
rect 96540 87012 96596 87014
rect 96620 87012 96676 87014
rect 81020 86522 81076 86524
rect 81100 86522 81156 86524
rect 81180 86522 81236 86524
rect 81260 86522 81316 86524
rect 81020 86470 81046 86522
rect 81046 86470 81076 86522
rect 81100 86470 81110 86522
rect 81110 86470 81156 86522
rect 81180 86470 81226 86522
rect 81226 86470 81236 86522
rect 81260 86470 81290 86522
rect 81290 86470 81316 86522
rect 81020 86468 81076 86470
rect 81100 86468 81156 86470
rect 81180 86468 81236 86470
rect 81260 86468 81316 86470
rect 111740 86522 111796 86524
rect 111820 86522 111876 86524
rect 111900 86522 111956 86524
rect 111980 86522 112036 86524
rect 111740 86470 111766 86522
rect 111766 86470 111796 86522
rect 111820 86470 111830 86522
rect 111830 86470 111876 86522
rect 111900 86470 111946 86522
rect 111946 86470 111956 86522
rect 111980 86470 112010 86522
rect 112010 86470 112036 86522
rect 111740 86468 111796 86470
rect 111820 86468 111876 86470
rect 111900 86468 111956 86470
rect 111980 86468 112036 86470
rect 96380 85978 96436 85980
rect 96460 85978 96516 85980
rect 96540 85978 96596 85980
rect 96620 85978 96676 85980
rect 96380 85926 96406 85978
rect 96406 85926 96436 85978
rect 96460 85926 96470 85978
rect 96470 85926 96516 85978
rect 96540 85926 96586 85978
rect 96586 85926 96596 85978
rect 96620 85926 96650 85978
rect 96650 85926 96676 85978
rect 96380 85924 96436 85926
rect 96460 85924 96516 85926
rect 96540 85924 96596 85926
rect 96620 85924 96676 85926
rect 81020 85434 81076 85436
rect 81100 85434 81156 85436
rect 81180 85434 81236 85436
rect 81260 85434 81316 85436
rect 81020 85382 81046 85434
rect 81046 85382 81076 85434
rect 81100 85382 81110 85434
rect 81110 85382 81156 85434
rect 81180 85382 81226 85434
rect 81226 85382 81236 85434
rect 81260 85382 81290 85434
rect 81290 85382 81316 85434
rect 81020 85380 81076 85382
rect 81100 85380 81156 85382
rect 81180 85380 81236 85382
rect 81260 85380 81316 85382
rect 111740 85434 111796 85436
rect 111820 85434 111876 85436
rect 111900 85434 111956 85436
rect 111980 85434 112036 85436
rect 111740 85382 111766 85434
rect 111766 85382 111796 85434
rect 111820 85382 111830 85434
rect 111830 85382 111876 85434
rect 111900 85382 111946 85434
rect 111946 85382 111956 85434
rect 111980 85382 112010 85434
rect 112010 85382 112036 85434
rect 111740 85380 111796 85382
rect 111820 85380 111876 85382
rect 111900 85380 111956 85382
rect 111980 85380 112036 85382
rect 96380 84890 96436 84892
rect 96460 84890 96516 84892
rect 96540 84890 96596 84892
rect 96620 84890 96676 84892
rect 96380 84838 96406 84890
rect 96406 84838 96436 84890
rect 96460 84838 96470 84890
rect 96470 84838 96516 84890
rect 96540 84838 96586 84890
rect 96586 84838 96596 84890
rect 96620 84838 96650 84890
rect 96650 84838 96676 84890
rect 96380 84836 96436 84838
rect 96460 84836 96516 84838
rect 96540 84836 96596 84838
rect 96620 84836 96676 84838
rect 81020 84346 81076 84348
rect 81100 84346 81156 84348
rect 81180 84346 81236 84348
rect 81260 84346 81316 84348
rect 81020 84294 81046 84346
rect 81046 84294 81076 84346
rect 81100 84294 81110 84346
rect 81110 84294 81156 84346
rect 81180 84294 81226 84346
rect 81226 84294 81236 84346
rect 81260 84294 81290 84346
rect 81290 84294 81316 84346
rect 81020 84292 81076 84294
rect 81100 84292 81156 84294
rect 81180 84292 81236 84294
rect 81260 84292 81316 84294
rect 111740 84346 111796 84348
rect 111820 84346 111876 84348
rect 111900 84346 111956 84348
rect 111980 84346 112036 84348
rect 111740 84294 111766 84346
rect 111766 84294 111796 84346
rect 111820 84294 111830 84346
rect 111830 84294 111876 84346
rect 111900 84294 111946 84346
rect 111946 84294 111956 84346
rect 111980 84294 112010 84346
rect 112010 84294 112036 84346
rect 111740 84292 111796 84294
rect 111820 84292 111876 84294
rect 111900 84292 111956 84294
rect 111980 84292 112036 84294
rect 96380 83802 96436 83804
rect 96460 83802 96516 83804
rect 96540 83802 96596 83804
rect 96620 83802 96676 83804
rect 96380 83750 96406 83802
rect 96406 83750 96436 83802
rect 96460 83750 96470 83802
rect 96470 83750 96516 83802
rect 96540 83750 96586 83802
rect 96586 83750 96596 83802
rect 96620 83750 96650 83802
rect 96650 83750 96676 83802
rect 96380 83748 96436 83750
rect 96460 83748 96516 83750
rect 96540 83748 96596 83750
rect 96620 83748 96676 83750
rect 81020 83258 81076 83260
rect 81100 83258 81156 83260
rect 81180 83258 81236 83260
rect 81260 83258 81316 83260
rect 81020 83206 81046 83258
rect 81046 83206 81076 83258
rect 81100 83206 81110 83258
rect 81110 83206 81156 83258
rect 81180 83206 81226 83258
rect 81226 83206 81236 83258
rect 81260 83206 81290 83258
rect 81290 83206 81316 83258
rect 81020 83204 81076 83206
rect 81100 83204 81156 83206
rect 81180 83204 81236 83206
rect 81260 83204 81316 83206
rect 111740 83258 111796 83260
rect 111820 83258 111876 83260
rect 111900 83258 111956 83260
rect 111980 83258 112036 83260
rect 111740 83206 111766 83258
rect 111766 83206 111796 83258
rect 111820 83206 111830 83258
rect 111830 83206 111876 83258
rect 111900 83206 111946 83258
rect 111946 83206 111956 83258
rect 111980 83206 112010 83258
rect 112010 83206 112036 83258
rect 111740 83204 111796 83206
rect 111820 83204 111876 83206
rect 111900 83204 111956 83206
rect 111980 83204 112036 83206
rect 96380 82714 96436 82716
rect 96460 82714 96516 82716
rect 96540 82714 96596 82716
rect 96620 82714 96676 82716
rect 96380 82662 96406 82714
rect 96406 82662 96436 82714
rect 96460 82662 96470 82714
rect 96470 82662 96516 82714
rect 96540 82662 96586 82714
rect 96586 82662 96596 82714
rect 96620 82662 96650 82714
rect 96650 82662 96676 82714
rect 96380 82660 96436 82662
rect 96460 82660 96516 82662
rect 96540 82660 96596 82662
rect 96620 82660 96676 82662
rect 81020 82170 81076 82172
rect 81100 82170 81156 82172
rect 81180 82170 81236 82172
rect 81260 82170 81316 82172
rect 81020 82118 81046 82170
rect 81046 82118 81076 82170
rect 81100 82118 81110 82170
rect 81110 82118 81156 82170
rect 81180 82118 81226 82170
rect 81226 82118 81236 82170
rect 81260 82118 81290 82170
rect 81290 82118 81316 82170
rect 81020 82116 81076 82118
rect 81100 82116 81156 82118
rect 81180 82116 81236 82118
rect 81260 82116 81316 82118
rect 111740 82170 111796 82172
rect 111820 82170 111876 82172
rect 111900 82170 111956 82172
rect 111980 82170 112036 82172
rect 111740 82118 111766 82170
rect 111766 82118 111796 82170
rect 111820 82118 111830 82170
rect 111830 82118 111876 82170
rect 111900 82118 111946 82170
rect 111946 82118 111956 82170
rect 111980 82118 112010 82170
rect 112010 82118 112036 82170
rect 111740 82116 111796 82118
rect 111820 82116 111876 82118
rect 111900 82116 111956 82118
rect 111980 82116 112036 82118
rect 96380 81626 96436 81628
rect 96460 81626 96516 81628
rect 96540 81626 96596 81628
rect 96620 81626 96676 81628
rect 96380 81574 96406 81626
rect 96406 81574 96436 81626
rect 96460 81574 96470 81626
rect 96470 81574 96516 81626
rect 96540 81574 96586 81626
rect 96586 81574 96596 81626
rect 96620 81574 96650 81626
rect 96650 81574 96676 81626
rect 96380 81572 96436 81574
rect 96460 81572 96516 81574
rect 96540 81572 96596 81574
rect 96620 81572 96676 81574
rect 81020 81082 81076 81084
rect 81100 81082 81156 81084
rect 81180 81082 81236 81084
rect 81260 81082 81316 81084
rect 81020 81030 81046 81082
rect 81046 81030 81076 81082
rect 81100 81030 81110 81082
rect 81110 81030 81156 81082
rect 81180 81030 81226 81082
rect 81226 81030 81236 81082
rect 81260 81030 81290 81082
rect 81290 81030 81316 81082
rect 81020 81028 81076 81030
rect 81100 81028 81156 81030
rect 81180 81028 81236 81030
rect 81260 81028 81316 81030
rect 111740 81082 111796 81084
rect 111820 81082 111876 81084
rect 111900 81082 111956 81084
rect 111980 81082 112036 81084
rect 111740 81030 111766 81082
rect 111766 81030 111796 81082
rect 111820 81030 111830 81082
rect 111830 81030 111876 81082
rect 111900 81030 111946 81082
rect 111946 81030 111956 81082
rect 111980 81030 112010 81082
rect 112010 81030 112036 81082
rect 111740 81028 111796 81030
rect 111820 81028 111876 81030
rect 111900 81028 111956 81030
rect 111980 81028 112036 81030
rect 96380 80538 96436 80540
rect 96460 80538 96516 80540
rect 96540 80538 96596 80540
rect 96620 80538 96676 80540
rect 96380 80486 96406 80538
rect 96406 80486 96436 80538
rect 96460 80486 96470 80538
rect 96470 80486 96516 80538
rect 96540 80486 96586 80538
rect 96586 80486 96596 80538
rect 96620 80486 96650 80538
rect 96650 80486 96676 80538
rect 96380 80484 96436 80486
rect 96460 80484 96516 80486
rect 96540 80484 96596 80486
rect 96620 80484 96676 80486
rect 81020 79994 81076 79996
rect 81100 79994 81156 79996
rect 81180 79994 81236 79996
rect 81260 79994 81316 79996
rect 81020 79942 81046 79994
rect 81046 79942 81076 79994
rect 81100 79942 81110 79994
rect 81110 79942 81156 79994
rect 81180 79942 81226 79994
rect 81226 79942 81236 79994
rect 81260 79942 81290 79994
rect 81290 79942 81316 79994
rect 81020 79940 81076 79942
rect 81100 79940 81156 79942
rect 81180 79940 81236 79942
rect 81260 79940 81316 79942
rect 111740 79994 111796 79996
rect 111820 79994 111876 79996
rect 111900 79994 111956 79996
rect 111980 79994 112036 79996
rect 111740 79942 111766 79994
rect 111766 79942 111796 79994
rect 111820 79942 111830 79994
rect 111830 79942 111876 79994
rect 111900 79942 111946 79994
rect 111946 79942 111956 79994
rect 111980 79942 112010 79994
rect 112010 79942 112036 79994
rect 111740 79940 111796 79942
rect 111820 79940 111876 79942
rect 111900 79940 111956 79942
rect 111980 79940 112036 79942
rect 96380 79450 96436 79452
rect 96460 79450 96516 79452
rect 96540 79450 96596 79452
rect 96620 79450 96676 79452
rect 96380 79398 96406 79450
rect 96406 79398 96436 79450
rect 96460 79398 96470 79450
rect 96470 79398 96516 79450
rect 96540 79398 96586 79450
rect 96586 79398 96596 79450
rect 96620 79398 96650 79450
rect 96650 79398 96676 79450
rect 96380 79396 96436 79398
rect 96460 79396 96516 79398
rect 96540 79396 96596 79398
rect 96620 79396 96676 79398
rect 81020 78906 81076 78908
rect 81100 78906 81156 78908
rect 81180 78906 81236 78908
rect 81260 78906 81316 78908
rect 81020 78854 81046 78906
rect 81046 78854 81076 78906
rect 81100 78854 81110 78906
rect 81110 78854 81156 78906
rect 81180 78854 81226 78906
rect 81226 78854 81236 78906
rect 81260 78854 81290 78906
rect 81290 78854 81316 78906
rect 81020 78852 81076 78854
rect 81100 78852 81156 78854
rect 81180 78852 81236 78854
rect 81260 78852 81316 78854
rect 111740 78906 111796 78908
rect 111820 78906 111876 78908
rect 111900 78906 111956 78908
rect 111980 78906 112036 78908
rect 111740 78854 111766 78906
rect 111766 78854 111796 78906
rect 111820 78854 111830 78906
rect 111830 78854 111876 78906
rect 111900 78854 111946 78906
rect 111946 78854 111956 78906
rect 111980 78854 112010 78906
rect 112010 78854 112036 78906
rect 111740 78852 111796 78854
rect 111820 78852 111876 78854
rect 111900 78852 111956 78854
rect 111980 78852 112036 78854
rect 96380 78362 96436 78364
rect 96460 78362 96516 78364
rect 96540 78362 96596 78364
rect 96620 78362 96676 78364
rect 96380 78310 96406 78362
rect 96406 78310 96436 78362
rect 96460 78310 96470 78362
rect 96470 78310 96516 78362
rect 96540 78310 96586 78362
rect 96586 78310 96596 78362
rect 96620 78310 96650 78362
rect 96650 78310 96676 78362
rect 96380 78308 96436 78310
rect 96460 78308 96516 78310
rect 96540 78308 96596 78310
rect 96620 78308 96676 78310
rect 81020 77818 81076 77820
rect 81100 77818 81156 77820
rect 81180 77818 81236 77820
rect 81260 77818 81316 77820
rect 81020 77766 81046 77818
rect 81046 77766 81076 77818
rect 81100 77766 81110 77818
rect 81110 77766 81156 77818
rect 81180 77766 81226 77818
rect 81226 77766 81236 77818
rect 81260 77766 81290 77818
rect 81290 77766 81316 77818
rect 81020 77764 81076 77766
rect 81100 77764 81156 77766
rect 81180 77764 81236 77766
rect 81260 77764 81316 77766
rect 111740 77818 111796 77820
rect 111820 77818 111876 77820
rect 111900 77818 111956 77820
rect 111980 77818 112036 77820
rect 111740 77766 111766 77818
rect 111766 77766 111796 77818
rect 111820 77766 111830 77818
rect 111830 77766 111876 77818
rect 111900 77766 111946 77818
rect 111946 77766 111956 77818
rect 111980 77766 112010 77818
rect 112010 77766 112036 77818
rect 111740 77764 111796 77766
rect 111820 77764 111876 77766
rect 111900 77764 111956 77766
rect 111980 77764 112036 77766
rect 96380 77274 96436 77276
rect 96460 77274 96516 77276
rect 96540 77274 96596 77276
rect 96620 77274 96676 77276
rect 96380 77222 96406 77274
rect 96406 77222 96436 77274
rect 96460 77222 96470 77274
rect 96470 77222 96516 77274
rect 96540 77222 96586 77274
rect 96586 77222 96596 77274
rect 96620 77222 96650 77274
rect 96650 77222 96676 77274
rect 96380 77220 96436 77222
rect 96460 77220 96516 77222
rect 96540 77220 96596 77222
rect 96620 77220 96676 77222
rect 81020 76730 81076 76732
rect 81100 76730 81156 76732
rect 81180 76730 81236 76732
rect 81260 76730 81316 76732
rect 81020 76678 81046 76730
rect 81046 76678 81076 76730
rect 81100 76678 81110 76730
rect 81110 76678 81156 76730
rect 81180 76678 81226 76730
rect 81226 76678 81236 76730
rect 81260 76678 81290 76730
rect 81290 76678 81316 76730
rect 81020 76676 81076 76678
rect 81100 76676 81156 76678
rect 81180 76676 81236 76678
rect 81260 76676 81316 76678
rect 111740 76730 111796 76732
rect 111820 76730 111876 76732
rect 111900 76730 111956 76732
rect 111980 76730 112036 76732
rect 111740 76678 111766 76730
rect 111766 76678 111796 76730
rect 111820 76678 111830 76730
rect 111830 76678 111876 76730
rect 111900 76678 111946 76730
rect 111946 76678 111956 76730
rect 111980 76678 112010 76730
rect 112010 76678 112036 76730
rect 111740 76676 111796 76678
rect 111820 76676 111876 76678
rect 111900 76676 111956 76678
rect 111980 76676 112036 76678
rect 96380 76186 96436 76188
rect 96460 76186 96516 76188
rect 96540 76186 96596 76188
rect 96620 76186 96676 76188
rect 96380 76134 96406 76186
rect 96406 76134 96436 76186
rect 96460 76134 96470 76186
rect 96470 76134 96516 76186
rect 96540 76134 96586 76186
rect 96586 76134 96596 76186
rect 96620 76134 96650 76186
rect 96650 76134 96676 76186
rect 96380 76132 96436 76134
rect 96460 76132 96516 76134
rect 96540 76132 96596 76134
rect 96620 76132 96676 76134
rect 81020 75642 81076 75644
rect 81100 75642 81156 75644
rect 81180 75642 81236 75644
rect 81260 75642 81316 75644
rect 81020 75590 81046 75642
rect 81046 75590 81076 75642
rect 81100 75590 81110 75642
rect 81110 75590 81156 75642
rect 81180 75590 81226 75642
rect 81226 75590 81236 75642
rect 81260 75590 81290 75642
rect 81290 75590 81316 75642
rect 81020 75588 81076 75590
rect 81100 75588 81156 75590
rect 81180 75588 81236 75590
rect 81260 75588 81316 75590
rect 111740 75642 111796 75644
rect 111820 75642 111876 75644
rect 111900 75642 111956 75644
rect 111980 75642 112036 75644
rect 111740 75590 111766 75642
rect 111766 75590 111796 75642
rect 111820 75590 111830 75642
rect 111830 75590 111876 75642
rect 111900 75590 111946 75642
rect 111946 75590 111956 75642
rect 111980 75590 112010 75642
rect 112010 75590 112036 75642
rect 111740 75588 111796 75590
rect 111820 75588 111876 75590
rect 111900 75588 111956 75590
rect 111980 75588 112036 75590
rect 96380 75098 96436 75100
rect 96460 75098 96516 75100
rect 96540 75098 96596 75100
rect 96620 75098 96676 75100
rect 96380 75046 96406 75098
rect 96406 75046 96436 75098
rect 96460 75046 96470 75098
rect 96470 75046 96516 75098
rect 96540 75046 96586 75098
rect 96586 75046 96596 75098
rect 96620 75046 96650 75098
rect 96650 75046 96676 75098
rect 96380 75044 96436 75046
rect 96460 75044 96516 75046
rect 96540 75044 96596 75046
rect 96620 75044 96676 75046
rect 81020 74554 81076 74556
rect 81100 74554 81156 74556
rect 81180 74554 81236 74556
rect 81260 74554 81316 74556
rect 81020 74502 81046 74554
rect 81046 74502 81076 74554
rect 81100 74502 81110 74554
rect 81110 74502 81156 74554
rect 81180 74502 81226 74554
rect 81226 74502 81236 74554
rect 81260 74502 81290 74554
rect 81290 74502 81316 74554
rect 81020 74500 81076 74502
rect 81100 74500 81156 74502
rect 81180 74500 81236 74502
rect 81260 74500 81316 74502
rect 111740 74554 111796 74556
rect 111820 74554 111876 74556
rect 111900 74554 111956 74556
rect 111980 74554 112036 74556
rect 111740 74502 111766 74554
rect 111766 74502 111796 74554
rect 111820 74502 111830 74554
rect 111830 74502 111876 74554
rect 111900 74502 111946 74554
rect 111946 74502 111956 74554
rect 111980 74502 112010 74554
rect 112010 74502 112036 74554
rect 111740 74500 111796 74502
rect 111820 74500 111876 74502
rect 111900 74500 111956 74502
rect 111980 74500 112036 74502
rect 96380 74010 96436 74012
rect 96460 74010 96516 74012
rect 96540 74010 96596 74012
rect 96620 74010 96676 74012
rect 96380 73958 96406 74010
rect 96406 73958 96436 74010
rect 96460 73958 96470 74010
rect 96470 73958 96516 74010
rect 96540 73958 96586 74010
rect 96586 73958 96596 74010
rect 96620 73958 96650 74010
rect 96650 73958 96676 74010
rect 96380 73956 96436 73958
rect 96460 73956 96516 73958
rect 96540 73956 96596 73958
rect 96620 73956 96676 73958
rect 81020 73466 81076 73468
rect 81100 73466 81156 73468
rect 81180 73466 81236 73468
rect 81260 73466 81316 73468
rect 81020 73414 81046 73466
rect 81046 73414 81076 73466
rect 81100 73414 81110 73466
rect 81110 73414 81156 73466
rect 81180 73414 81226 73466
rect 81226 73414 81236 73466
rect 81260 73414 81290 73466
rect 81290 73414 81316 73466
rect 81020 73412 81076 73414
rect 81100 73412 81156 73414
rect 81180 73412 81236 73414
rect 81260 73412 81316 73414
rect 111740 73466 111796 73468
rect 111820 73466 111876 73468
rect 111900 73466 111956 73468
rect 111980 73466 112036 73468
rect 111740 73414 111766 73466
rect 111766 73414 111796 73466
rect 111820 73414 111830 73466
rect 111830 73414 111876 73466
rect 111900 73414 111946 73466
rect 111946 73414 111956 73466
rect 111980 73414 112010 73466
rect 112010 73414 112036 73466
rect 111740 73412 111796 73414
rect 111820 73412 111876 73414
rect 111900 73412 111956 73414
rect 111980 73412 112036 73414
rect 96380 72922 96436 72924
rect 96460 72922 96516 72924
rect 96540 72922 96596 72924
rect 96620 72922 96676 72924
rect 96380 72870 96406 72922
rect 96406 72870 96436 72922
rect 96460 72870 96470 72922
rect 96470 72870 96516 72922
rect 96540 72870 96586 72922
rect 96586 72870 96596 72922
rect 96620 72870 96650 72922
rect 96650 72870 96676 72922
rect 96380 72868 96436 72870
rect 96460 72868 96516 72870
rect 96540 72868 96596 72870
rect 96620 72868 96676 72870
rect 81020 72378 81076 72380
rect 81100 72378 81156 72380
rect 81180 72378 81236 72380
rect 81260 72378 81316 72380
rect 81020 72326 81046 72378
rect 81046 72326 81076 72378
rect 81100 72326 81110 72378
rect 81110 72326 81156 72378
rect 81180 72326 81226 72378
rect 81226 72326 81236 72378
rect 81260 72326 81290 72378
rect 81290 72326 81316 72378
rect 81020 72324 81076 72326
rect 81100 72324 81156 72326
rect 81180 72324 81236 72326
rect 81260 72324 81316 72326
rect 111740 72378 111796 72380
rect 111820 72378 111876 72380
rect 111900 72378 111956 72380
rect 111980 72378 112036 72380
rect 111740 72326 111766 72378
rect 111766 72326 111796 72378
rect 111820 72326 111830 72378
rect 111830 72326 111876 72378
rect 111900 72326 111946 72378
rect 111946 72326 111956 72378
rect 111980 72326 112010 72378
rect 112010 72326 112036 72378
rect 111740 72324 111796 72326
rect 111820 72324 111876 72326
rect 111900 72324 111956 72326
rect 111980 72324 112036 72326
rect 96380 71834 96436 71836
rect 96460 71834 96516 71836
rect 96540 71834 96596 71836
rect 96620 71834 96676 71836
rect 96380 71782 96406 71834
rect 96406 71782 96436 71834
rect 96460 71782 96470 71834
rect 96470 71782 96516 71834
rect 96540 71782 96586 71834
rect 96586 71782 96596 71834
rect 96620 71782 96650 71834
rect 96650 71782 96676 71834
rect 96380 71780 96436 71782
rect 96460 71780 96516 71782
rect 96540 71780 96596 71782
rect 96620 71780 96676 71782
rect 81020 71290 81076 71292
rect 81100 71290 81156 71292
rect 81180 71290 81236 71292
rect 81260 71290 81316 71292
rect 81020 71238 81046 71290
rect 81046 71238 81076 71290
rect 81100 71238 81110 71290
rect 81110 71238 81156 71290
rect 81180 71238 81226 71290
rect 81226 71238 81236 71290
rect 81260 71238 81290 71290
rect 81290 71238 81316 71290
rect 81020 71236 81076 71238
rect 81100 71236 81156 71238
rect 81180 71236 81236 71238
rect 81260 71236 81316 71238
rect 111740 71290 111796 71292
rect 111820 71290 111876 71292
rect 111900 71290 111956 71292
rect 111980 71290 112036 71292
rect 111740 71238 111766 71290
rect 111766 71238 111796 71290
rect 111820 71238 111830 71290
rect 111830 71238 111876 71290
rect 111900 71238 111946 71290
rect 111946 71238 111956 71290
rect 111980 71238 112010 71290
rect 112010 71238 112036 71290
rect 111740 71236 111796 71238
rect 111820 71236 111876 71238
rect 111900 71236 111956 71238
rect 111980 71236 112036 71238
rect 96380 70746 96436 70748
rect 96460 70746 96516 70748
rect 96540 70746 96596 70748
rect 96620 70746 96676 70748
rect 96380 70694 96406 70746
rect 96406 70694 96436 70746
rect 96460 70694 96470 70746
rect 96470 70694 96516 70746
rect 96540 70694 96586 70746
rect 96586 70694 96596 70746
rect 96620 70694 96650 70746
rect 96650 70694 96676 70746
rect 96380 70692 96436 70694
rect 96460 70692 96516 70694
rect 96540 70692 96596 70694
rect 96620 70692 96676 70694
rect 81020 70202 81076 70204
rect 81100 70202 81156 70204
rect 81180 70202 81236 70204
rect 81260 70202 81316 70204
rect 81020 70150 81046 70202
rect 81046 70150 81076 70202
rect 81100 70150 81110 70202
rect 81110 70150 81156 70202
rect 81180 70150 81226 70202
rect 81226 70150 81236 70202
rect 81260 70150 81290 70202
rect 81290 70150 81316 70202
rect 81020 70148 81076 70150
rect 81100 70148 81156 70150
rect 81180 70148 81236 70150
rect 81260 70148 81316 70150
rect 111740 70202 111796 70204
rect 111820 70202 111876 70204
rect 111900 70202 111956 70204
rect 111980 70202 112036 70204
rect 111740 70150 111766 70202
rect 111766 70150 111796 70202
rect 111820 70150 111830 70202
rect 111830 70150 111876 70202
rect 111900 70150 111946 70202
rect 111946 70150 111956 70202
rect 111980 70150 112010 70202
rect 112010 70150 112036 70202
rect 111740 70148 111796 70150
rect 111820 70148 111876 70150
rect 111900 70148 111956 70150
rect 111980 70148 112036 70150
rect 96380 69658 96436 69660
rect 96460 69658 96516 69660
rect 96540 69658 96596 69660
rect 96620 69658 96676 69660
rect 96380 69606 96406 69658
rect 96406 69606 96436 69658
rect 96460 69606 96470 69658
rect 96470 69606 96516 69658
rect 96540 69606 96586 69658
rect 96586 69606 96596 69658
rect 96620 69606 96650 69658
rect 96650 69606 96676 69658
rect 96380 69604 96436 69606
rect 96460 69604 96516 69606
rect 96540 69604 96596 69606
rect 96620 69604 96676 69606
rect 81020 69114 81076 69116
rect 81100 69114 81156 69116
rect 81180 69114 81236 69116
rect 81260 69114 81316 69116
rect 81020 69062 81046 69114
rect 81046 69062 81076 69114
rect 81100 69062 81110 69114
rect 81110 69062 81156 69114
rect 81180 69062 81226 69114
rect 81226 69062 81236 69114
rect 81260 69062 81290 69114
rect 81290 69062 81316 69114
rect 81020 69060 81076 69062
rect 81100 69060 81156 69062
rect 81180 69060 81236 69062
rect 81260 69060 81316 69062
rect 111740 69114 111796 69116
rect 111820 69114 111876 69116
rect 111900 69114 111956 69116
rect 111980 69114 112036 69116
rect 111740 69062 111766 69114
rect 111766 69062 111796 69114
rect 111820 69062 111830 69114
rect 111830 69062 111876 69114
rect 111900 69062 111946 69114
rect 111946 69062 111956 69114
rect 111980 69062 112010 69114
rect 112010 69062 112036 69114
rect 111740 69060 111796 69062
rect 111820 69060 111876 69062
rect 111900 69060 111956 69062
rect 111980 69060 112036 69062
rect 96380 68570 96436 68572
rect 96460 68570 96516 68572
rect 96540 68570 96596 68572
rect 96620 68570 96676 68572
rect 96380 68518 96406 68570
rect 96406 68518 96436 68570
rect 96460 68518 96470 68570
rect 96470 68518 96516 68570
rect 96540 68518 96586 68570
rect 96586 68518 96596 68570
rect 96620 68518 96650 68570
rect 96650 68518 96676 68570
rect 96380 68516 96436 68518
rect 96460 68516 96516 68518
rect 96540 68516 96596 68518
rect 96620 68516 96676 68518
rect 81020 68026 81076 68028
rect 81100 68026 81156 68028
rect 81180 68026 81236 68028
rect 81260 68026 81316 68028
rect 81020 67974 81046 68026
rect 81046 67974 81076 68026
rect 81100 67974 81110 68026
rect 81110 67974 81156 68026
rect 81180 67974 81226 68026
rect 81226 67974 81236 68026
rect 81260 67974 81290 68026
rect 81290 67974 81316 68026
rect 81020 67972 81076 67974
rect 81100 67972 81156 67974
rect 81180 67972 81236 67974
rect 81260 67972 81316 67974
rect 111740 68026 111796 68028
rect 111820 68026 111876 68028
rect 111900 68026 111956 68028
rect 111980 68026 112036 68028
rect 111740 67974 111766 68026
rect 111766 67974 111796 68026
rect 111820 67974 111830 68026
rect 111830 67974 111876 68026
rect 111900 67974 111946 68026
rect 111946 67974 111956 68026
rect 111980 67974 112010 68026
rect 112010 67974 112036 68026
rect 111740 67972 111796 67974
rect 111820 67972 111876 67974
rect 111900 67972 111956 67974
rect 111980 67972 112036 67974
rect 96380 67482 96436 67484
rect 96460 67482 96516 67484
rect 96540 67482 96596 67484
rect 96620 67482 96676 67484
rect 96380 67430 96406 67482
rect 96406 67430 96436 67482
rect 96460 67430 96470 67482
rect 96470 67430 96516 67482
rect 96540 67430 96586 67482
rect 96586 67430 96596 67482
rect 96620 67430 96650 67482
rect 96650 67430 96676 67482
rect 96380 67428 96436 67430
rect 96460 67428 96516 67430
rect 96540 67428 96596 67430
rect 96620 67428 96676 67430
rect 81020 66938 81076 66940
rect 81100 66938 81156 66940
rect 81180 66938 81236 66940
rect 81260 66938 81316 66940
rect 81020 66886 81046 66938
rect 81046 66886 81076 66938
rect 81100 66886 81110 66938
rect 81110 66886 81156 66938
rect 81180 66886 81226 66938
rect 81226 66886 81236 66938
rect 81260 66886 81290 66938
rect 81290 66886 81316 66938
rect 81020 66884 81076 66886
rect 81100 66884 81156 66886
rect 81180 66884 81236 66886
rect 81260 66884 81316 66886
rect 111740 66938 111796 66940
rect 111820 66938 111876 66940
rect 111900 66938 111956 66940
rect 111980 66938 112036 66940
rect 111740 66886 111766 66938
rect 111766 66886 111796 66938
rect 111820 66886 111830 66938
rect 111830 66886 111876 66938
rect 111900 66886 111946 66938
rect 111946 66886 111956 66938
rect 111980 66886 112010 66938
rect 112010 66886 112036 66938
rect 111740 66884 111796 66886
rect 111820 66884 111876 66886
rect 111900 66884 111956 66886
rect 111980 66884 112036 66886
rect 96380 66394 96436 66396
rect 96460 66394 96516 66396
rect 96540 66394 96596 66396
rect 96620 66394 96676 66396
rect 96380 66342 96406 66394
rect 96406 66342 96436 66394
rect 96460 66342 96470 66394
rect 96470 66342 96516 66394
rect 96540 66342 96586 66394
rect 96586 66342 96596 66394
rect 96620 66342 96650 66394
rect 96650 66342 96676 66394
rect 96380 66340 96436 66342
rect 96460 66340 96516 66342
rect 96540 66340 96596 66342
rect 96620 66340 96676 66342
rect 81020 65850 81076 65852
rect 81100 65850 81156 65852
rect 81180 65850 81236 65852
rect 81260 65850 81316 65852
rect 81020 65798 81046 65850
rect 81046 65798 81076 65850
rect 81100 65798 81110 65850
rect 81110 65798 81156 65850
rect 81180 65798 81226 65850
rect 81226 65798 81236 65850
rect 81260 65798 81290 65850
rect 81290 65798 81316 65850
rect 81020 65796 81076 65798
rect 81100 65796 81156 65798
rect 81180 65796 81236 65798
rect 81260 65796 81316 65798
rect 111740 65850 111796 65852
rect 111820 65850 111876 65852
rect 111900 65850 111956 65852
rect 111980 65850 112036 65852
rect 111740 65798 111766 65850
rect 111766 65798 111796 65850
rect 111820 65798 111830 65850
rect 111830 65798 111876 65850
rect 111900 65798 111946 65850
rect 111946 65798 111956 65850
rect 111980 65798 112010 65850
rect 112010 65798 112036 65850
rect 111740 65796 111796 65798
rect 111820 65796 111876 65798
rect 111900 65796 111956 65798
rect 111980 65796 112036 65798
rect 96380 65306 96436 65308
rect 96460 65306 96516 65308
rect 96540 65306 96596 65308
rect 96620 65306 96676 65308
rect 96380 65254 96406 65306
rect 96406 65254 96436 65306
rect 96460 65254 96470 65306
rect 96470 65254 96516 65306
rect 96540 65254 96586 65306
rect 96586 65254 96596 65306
rect 96620 65254 96650 65306
rect 96650 65254 96676 65306
rect 96380 65252 96436 65254
rect 96460 65252 96516 65254
rect 96540 65252 96596 65254
rect 96620 65252 96676 65254
rect 81020 64762 81076 64764
rect 81100 64762 81156 64764
rect 81180 64762 81236 64764
rect 81260 64762 81316 64764
rect 81020 64710 81046 64762
rect 81046 64710 81076 64762
rect 81100 64710 81110 64762
rect 81110 64710 81156 64762
rect 81180 64710 81226 64762
rect 81226 64710 81236 64762
rect 81260 64710 81290 64762
rect 81290 64710 81316 64762
rect 81020 64708 81076 64710
rect 81100 64708 81156 64710
rect 81180 64708 81236 64710
rect 81260 64708 81316 64710
rect 111740 64762 111796 64764
rect 111820 64762 111876 64764
rect 111900 64762 111956 64764
rect 111980 64762 112036 64764
rect 111740 64710 111766 64762
rect 111766 64710 111796 64762
rect 111820 64710 111830 64762
rect 111830 64710 111876 64762
rect 111900 64710 111946 64762
rect 111946 64710 111956 64762
rect 111980 64710 112010 64762
rect 112010 64710 112036 64762
rect 111740 64708 111796 64710
rect 111820 64708 111876 64710
rect 111900 64708 111956 64710
rect 111980 64708 112036 64710
rect 96380 64218 96436 64220
rect 96460 64218 96516 64220
rect 96540 64218 96596 64220
rect 96620 64218 96676 64220
rect 96380 64166 96406 64218
rect 96406 64166 96436 64218
rect 96460 64166 96470 64218
rect 96470 64166 96516 64218
rect 96540 64166 96586 64218
rect 96586 64166 96596 64218
rect 96620 64166 96650 64218
rect 96650 64166 96676 64218
rect 96380 64164 96436 64166
rect 96460 64164 96516 64166
rect 96540 64164 96596 64166
rect 96620 64164 96676 64166
rect 81020 63674 81076 63676
rect 81100 63674 81156 63676
rect 81180 63674 81236 63676
rect 81260 63674 81316 63676
rect 81020 63622 81046 63674
rect 81046 63622 81076 63674
rect 81100 63622 81110 63674
rect 81110 63622 81156 63674
rect 81180 63622 81226 63674
rect 81226 63622 81236 63674
rect 81260 63622 81290 63674
rect 81290 63622 81316 63674
rect 81020 63620 81076 63622
rect 81100 63620 81156 63622
rect 81180 63620 81236 63622
rect 81260 63620 81316 63622
rect 111740 63674 111796 63676
rect 111820 63674 111876 63676
rect 111900 63674 111956 63676
rect 111980 63674 112036 63676
rect 111740 63622 111766 63674
rect 111766 63622 111796 63674
rect 111820 63622 111830 63674
rect 111830 63622 111876 63674
rect 111900 63622 111946 63674
rect 111946 63622 111956 63674
rect 111980 63622 112010 63674
rect 112010 63622 112036 63674
rect 111740 63620 111796 63622
rect 111820 63620 111876 63622
rect 111900 63620 111956 63622
rect 111980 63620 112036 63622
rect 96380 63130 96436 63132
rect 96460 63130 96516 63132
rect 96540 63130 96596 63132
rect 96620 63130 96676 63132
rect 96380 63078 96406 63130
rect 96406 63078 96436 63130
rect 96460 63078 96470 63130
rect 96470 63078 96516 63130
rect 96540 63078 96586 63130
rect 96586 63078 96596 63130
rect 96620 63078 96650 63130
rect 96650 63078 96676 63130
rect 96380 63076 96436 63078
rect 96460 63076 96516 63078
rect 96540 63076 96596 63078
rect 96620 63076 96676 63078
rect 81020 62586 81076 62588
rect 81100 62586 81156 62588
rect 81180 62586 81236 62588
rect 81260 62586 81316 62588
rect 81020 62534 81046 62586
rect 81046 62534 81076 62586
rect 81100 62534 81110 62586
rect 81110 62534 81156 62586
rect 81180 62534 81226 62586
rect 81226 62534 81236 62586
rect 81260 62534 81290 62586
rect 81290 62534 81316 62586
rect 81020 62532 81076 62534
rect 81100 62532 81156 62534
rect 81180 62532 81236 62534
rect 81260 62532 81316 62534
rect 111740 62586 111796 62588
rect 111820 62586 111876 62588
rect 111900 62586 111956 62588
rect 111980 62586 112036 62588
rect 111740 62534 111766 62586
rect 111766 62534 111796 62586
rect 111820 62534 111830 62586
rect 111830 62534 111876 62586
rect 111900 62534 111946 62586
rect 111946 62534 111956 62586
rect 111980 62534 112010 62586
rect 112010 62534 112036 62586
rect 111740 62532 111796 62534
rect 111820 62532 111876 62534
rect 111900 62532 111956 62534
rect 111980 62532 112036 62534
rect 96380 62042 96436 62044
rect 96460 62042 96516 62044
rect 96540 62042 96596 62044
rect 96620 62042 96676 62044
rect 96380 61990 96406 62042
rect 96406 61990 96436 62042
rect 96460 61990 96470 62042
rect 96470 61990 96516 62042
rect 96540 61990 96586 62042
rect 96586 61990 96596 62042
rect 96620 61990 96650 62042
rect 96650 61990 96676 62042
rect 96380 61988 96436 61990
rect 96460 61988 96516 61990
rect 96540 61988 96596 61990
rect 96620 61988 96676 61990
rect 81020 61498 81076 61500
rect 81100 61498 81156 61500
rect 81180 61498 81236 61500
rect 81260 61498 81316 61500
rect 81020 61446 81046 61498
rect 81046 61446 81076 61498
rect 81100 61446 81110 61498
rect 81110 61446 81156 61498
rect 81180 61446 81226 61498
rect 81226 61446 81236 61498
rect 81260 61446 81290 61498
rect 81290 61446 81316 61498
rect 81020 61444 81076 61446
rect 81100 61444 81156 61446
rect 81180 61444 81236 61446
rect 81260 61444 81316 61446
rect 111740 61498 111796 61500
rect 111820 61498 111876 61500
rect 111900 61498 111956 61500
rect 111980 61498 112036 61500
rect 111740 61446 111766 61498
rect 111766 61446 111796 61498
rect 111820 61446 111830 61498
rect 111830 61446 111876 61498
rect 111900 61446 111946 61498
rect 111946 61446 111956 61498
rect 111980 61446 112010 61498
rect 112010 61446 112036 61498
rect 111740 61444 111796 61446
rect 111820 61444 111876 61446
rect 111900 61444 111956 61446
rect 111980 61444 112036 61446
rect 96380 60954 96436 60956
rect 96460 60954 96516 60956
rect 96540 60954 96596 60956
rect 96620 60954 96676 60956
rect 96380 60902 96406 60954
rect 96406 60902 96436 60954
rect 96460 60902 96470 60954
rect 96470 60902 96516 60954
rect 96540 60902 96586 60954
rect 96586 60902 96596 60954
rect 96620 60902 96650 60954
rect 96650 60902 96676 60954
rect 96380 60900 96436 60902
rect 96460 60900 96516 60902
rect 96540 60900 96596 60902
rect 96620 60900 96676 60902
rect 81020 60410 81076 60412
rect 81100 60410 81156 60412
rect 81180 60410 81236 60412
rect 81260 60410 81316 60412
rect 81020 60358 81046 60410
rect 81046 60358 81076 60410
rect 81100 60358 81110 60410
rect 81110 60358 81156 60410
rect 81180 60358 81226 60410
rect 81226 60358 81236 60410
rect 81260 60358 81290 60410
rect 81290 60358 81316 60410
rect 81020 60356 81076 60358
rect 81100 60356 81156 60358
rect 81180 60356 81236 60358
rect 81260 60356 81316 60358
rect 111740 60410 111796 60412
rect 111820 60410 111876 60412
rect 111900 60410 111956 60412
rect 111980 60410 112036 60412
rect 111740 60358 111766 60410
rect 111766 60358 111796 60410
rect 111820 60358 111830 60410
rect 111830 60358 111876 60410
rect 111900 60358 111946 60410
rect 111946 60358 111956 60410
rect 111980 60358 112010 60410
rect 112010 60358 112036 60410
rect 111740 60356 111796 60358
rect 111820 60356 111876 60358
rect 111900 60356 111956 60358
rect 111980 60356 112036 60358
rect 96380 59866 96436 59868
rect 96460 59866 96516 59868
rect 96540 59866 96596 59868
rect 96620 59866 96676 59868
rect 96380 59814 96406 59866
rect 96406 59814 96436 59866
rect 96460 59814 96470 59866
rect 96470 59814 96516 59866
rect 96540 59814 96586 59866
rect 96586 59814 96596 59866
rect 96620 59814 96650 59866
rect 96650 59814 96676 59866
rect 96380 59812 96436 59814
rect 96460 59812 96516 59814
rect 96540 59812 96596 59814
rect 96620 59812 96676 59814
rect 81020 59322 81076 59324
rect 81100 59322 81156 59324
rect 81180 59322 81236 59324
rect 81260 59322 81316 59324
rect 81020 59270 81046 59322
rect 81046 59270 81076 59322
rect 81100 59270 81110 59322
rect 81110 59270 81156 59322
rect 81180 59270 81226 59322
rect 81226 59270 81236 59322
rect 81260 59270 81290 59322
rect 81290 59270 81316 59322
rect 81020 59268 81076 59270
rect 81100 59268 81156 59270
rect 81180 59268 81236 59270
rect 81260 59268 81316 59270
rect 111740 59322 111796 59324
rect 111820 59322 111876 59324
rect 111900 59322 111956 59324
rect 111980 59322 112036 59324
rect 111740 59270 111766 59322
rect 111766 59270 111796 59322
rect 111820 59270 111830 59322
rect 111830 59270 111876 59322
rect 111900 59270 111946 59322
rect 111946 59270 111956 59322
rect 111980 59270 112010 59322
rect 112010 59270 112036 59322
rect 111740 59268 111796 59270
rect 111820 59268 111876 59270
rect 111900 59268 111956 59270
rect 111980 59268 112036 59270
rect 96380 58778 96436 58780
rect 96460 58778 96516 58780
rect 96540 58778 96596 58780
rect 96620 58778 96676 58780
rect 96380 58726 96406 58778
rect 96406 58726 96436 58778
rect 96460 58726 96470 58778
rect 96470 58726 96516 58778
rect 96540 58726 96586 58778
rect 96586 58726 96596 58778
rect 96620 58726 96650 58778
rect 96650 58726 96676 58778
rect 96380 58724 96436 58726
rect 96460 58724 96516 58726
rect 96540 58724 96596 58726
rect 96620 58724 96676 58726
rect 81020 58234 81076 58236
rect 81100 58234 81156 58236
rect 81180 58234 81236 58236
rect 81260 58234 81316 58236
rect 81020 58182 81046 58234
rect 81046 58182 81076 58234
rect 81100 58182 81110 58234
rect 81110 58182 81156 58234
rect 81180 58182 81226 58234
rect 81226 58182 81236 58234
rect 81260 58182 81290 58234
rect 81290 58182 81316 58234
rect 81020 58180 81076 58182
rect 81100 58180 81156 58182
rect 81180 58180 81236 58182
rect 81260 58180 81316 58182
rect 111740 58234 111796 58236
rect 111820 58234 111876 58236
rect 111900 58234 111956 58236
rect 111980 58234 112036 58236
rect 111740 58182 111766 58234
rect 111766 58182 111796 58234
rect 111820 58182 111830 58234
rect 111830 58182 111876 58234
rect 111900 58182 111946 58234
rect 111946 58182 111956 58234
rect 111980 58182 112010 58234
rect 112010 58182 112036 58234
rect 111740 58180 111796 58182
rect 111820 58180 111876 58182
rect 111900 58180 111956 58182
rect 111980 58180 112036 58182
rect 96380 57690 96436 57692
rect 96460 57690 96516 57692
rect 96540 57690 96596 57692
rect 96620 57690 96676 57692
rect 96380 57638 96406 57690
rect 96406 57638 96436 57690
rect 96460 57638 96470 57690
rect 96470 57638 96516 57690
rect 96540 57638 96586 57690
rect 96586 57638 96596 57690
rect 96620 57638 96650 57690
rect 96650 57638 96676 57690
rect 96380 57636 96436 57638
rect 96460 57636 96516 57638
rect 96540 57636 96596 57638
rect 96620 57636 96676 57638
rect 81020 57146 81076 57148
rect 81100 57146 81156 57148
rect 81180 57146 81236 57148
rect 81260 57146 81316 57148
rect 81020 57094 81046 57146
rect 81046 57094 81076 57146
rect 81100 57094 81110 57146
rect 81110 57094 81156 57146
rect 81180 57094 81226 57146
rect 81226 57094 81236 57146
rect 81260 57094 81290 57146
rect 81290 57094 81316 57146
rect 81020 57092 81076 57094
rect 81100 57092 81156 57094
rect 81180 57092 81236 57094
rect 81260 57092 81316 57094
rect 111740 57146 111796 57148
rect 111820 57146 111876 57148
rect 111900 57146 111956 57148
rect 111980 57146 112036 57148
rect 111740 57094 111766 57146
rect 111766 57094 111796 57146
rect 111820 57094 111830 57146
rect 111830 57094 111876 57146
rect 111900 57094 111946 57146
rect 111946 57094 111956 57146
rect 111980 57094 112010 57146
rect 112010 57094 112036 57146
rect 111740 57092 111796 57094
rect 111820 57092 111876 57094
rect 111900 57092 111956 57094
rect 111980 57092 112036 57094
rect 96380 56602 96436 56604
rect 96460 56602 96516 56604
rect 96540 56602 96596 56604
rect 96620 56602 96676 56604
rect 96380 56550 96406 56602
rect 96406 56550 96436 56602
rect 96460 56550 96470 56602
rect 96470 56550 96516 56602
rect 96540 56550 96586 56602
rect 96586 56550 96596 56602
rect 96620 56550 96650 56602
rect 96650 56550 96676 56602
rect 96380 56548 96436 56550
rect 96460 56548 96516 56550
rect 96540 56548 96596 56550
rect 96620 56548 96676 56550
rect 81020 56058 81076 56060
rect 81100 56058 81156 56060
rect 81180 56058 81236 56060
rect 81260 56058 81316 56060
rect 81020 56006 81046 56058
rect 81046 56006 81076 56058
rect 81100 56006 81110 56058
rect 81110 56006 81156 56058
rect 81180 56006 81226 56058
rect 81226 56006 81236 56058
rect 81260 56006 81290 56058
rect 81290 56006 81316 56058
rect 81020 56004 81076 56006
rect 81100 56004 81156 56006
rect 81180 56004 81236 56006
rect 81260 56004 81316 56006
rect 111740 56058 111796 56060
rect 111820 56058 111876 56060
rect 111900 56058 111956 56060
rect 111980 56058 112036 56060
rect 111740 56006 111766 56058
rect 111766 56006 111796 56058
rect 111820 56006 111830 56058
rect 111830 56006 111876 56058
rect 111900 56006 111946 56058
rect 111946 56006 111956 56058
rect 111980 56006 112010 56058
rect 112010 56006 112036 56058
rect 111740 56004 111796 56006
rect 111820 56004 111876 56006
rect 111900 56004 111956 56006
rect 111980 56004 112036 56006
rect 96380 55514 96436 55516
rect 96460 55514 96516 55516
rect 96540 55514 96596 55516
rect 96620 55514 96676 55516
rect 96380 55462 96406 55514
rect 96406 55462 96436 55514
rect 96460 55462 96470 55514
rect 96470 55462 96516 55514
rect 96540 55462 96586 55514
rect 96586 55462 96596 55514
rect 96620 55462 96650 55514
rect 96650 55462 96676 55514
rect 96380 55460 96436 55462
rect 96460 55460 96516 55462
rect 96540 55460 96596 55462
rect 96620 55460 96676 55462
rect 81020 54970 81076 54972
rect 81100 54970 81156 54972
rect 81180 54970 81236 54972
rect 81260 54970 81316 54972
rect 81020 54918 81046 54970
rect 81046 54918 81076 54970
rect 81100 54918 81110 54970
rect 81110 54918 81156 54970
rect 81180 54918 81226 54970
rect 81226 54918 81236 54970
rect 81260 54918 81290 54970
rect 81290 54918 81316 54970
rect 81020 54916 81076 54918
rect 81100 54916 81156 54918
rect 81180 54916 81236 54918
rect 81260 54916 81316 54918
rect 111740 54970 111796 54972
rect 111820 54970 111876 54972
rect 111900 54970 111956 54972
rect 111980 54970 112036 54972
rect 111740 54918 111766 54970
rect 111766 54918 111796 54970
rect 111820 54918 111830 54970
rect 111830 54918 111876 54970
rect 111900 54918 111946 54970
rect 111946 54918 111956 54970
rect 111980 54918 112010 54970
rect 112010 54918 112036 54970
rect 111740 54916 111796 54918
rect 111820 54916 111876 54918
rect 111900 54916 111956 54918
rect 111980 54916 112036 54918
rect 96380 54426 96436 54428
rect 96460 54426 96516 54428
rect 96540 54426 96596 54428
rect 96620 54426 96676 54428
rect 96380 54374 96406 54426
rect 96406 54374 96436 54426
rect 96460 54374 96470 54426
rect 96470 54374 96516 54426
rect 96540 54374 96586 54426
rect 96586 54374 96596 54426
rect 96620 54374 96650 54426
rect 96650 54374 96676 54426
rect 96380 54372 96436 54374
rect 96460 54372 96516 54374
rect 96540 54372 96596 54374
rect 96620 54372 96676 54374
rect 81020 53882 81076 53884
rect 81100 53882 81156 53884
rect 81180 53882 81236 53884
rect 81260 53882 81316 53884
rect 81020 53830 81046 53882
rect 81046 53830 81076 53882
rect 81100 53830 81110 53882
rect 81110 53830 81156 53882
rect 81180 53830 81226 53882
rect 81226 53830 81236 53882
rect 81260 53830 81290 53882
rect 81290 53830 81316 53882
rect 81020 53828 81076 53830
rect 81100 53828 81156 53830
rect 81180 53828 81236 53830
rect 81260 53828 81316 53830
rect 111740 53882 111796 53884
rect 111820 53882 111876 53884
rect 111900 53882 111956 53884
rect 111980 53882 112036 53884
rect 111740 53830 111766 53882
rect 111766 53830 111796 53882
rect 111820 53830 111830 53882
rect 111830 53830 111876 53882
rect 111900 53830 111946 53882
rect 111946 53830 111956 53882
rect 111980 53830 112010 53882
rect 112010 53830 112036 53882
rect 111740 53828 111796 53830
rect 111820 53828 111876 53830
rect 111900 53828 111956 53830
rect 111980 53828 112036 53830
rect 96380 53338 96436 53340
rect 96460 53338 96516 53340
rect 96540 53338 96596 53340
rect 96620 53338 96676 53340
rect 96380 53286 96406 53338
rect 96406 53286 96436 53338
rect 96460 53286 96470 53338
rect 96470 53286 96516 53338
rect 96540 53286 96586 53338
rect 96586 53286 96596 53338
rect 96620 53286 96650 53338
rect 96650 53286 96676 53338
rect 96380 53284 96436 53286
rect 96460 53284 96516 53286
rect 96540 53284 96596 53286
rect 96620 53284 96676 53286
rect 81020 52794 81076 52796
rect 81100 52794 81156 52796
rect 81180 52794 81236 52796
rect 81260 52794 81316 52796
rect 81020 52742 81046 52794
rect 81046 52742 81076 52794
rect 81100 52742 81110 52794
rect 81110 52742 81156 52794
rect 81180 52742 81226 52794
rect 81226 52742 81236 52794
rect 81260 52742 81290 52794
rect 81290 52742 81316 52794
rect 81020 52740 81076 52742
rect 81100 52740 81156 52742
rect 81180 52740 81236 52742
rect 81260 52740 81316 52742
rect 111740 52794 111796 52796
rect 111820 52794 111876 52796
rect 111900 52794 111956 52796
rect 111980 52794 112036 52796
rect 111740 52742 111766 52794
rect 111766 52742 111796 52794
rect 111820 52742 111830 52794
rect 111830 52742 111876 52794
rect 111900 52742 111946 52794
rect 111946 52742 111956 52794
rect 111980 52742 112010 52794
rect 112010 52742 112036 52794
rect 111740 52740 111796 52742
rect 111820 52740 111876 52742
rect 111900 52740 111956 52742
rect 111980 52740 112036 52742
rect 96380 52250 96436 52252
rect 96460 52250 96516 52252
rect 96540 52250 96596 52252
rect 96620 52250 96676 52252
rect 96380 52198 96406 52250
rect 96406 52198 96436 52250
rect 96460 52198 96470 52250
rect 96470 52198 96516 52250
rect 96540 52198 96586 52250
rect 96586 52198 96596 52250
rect 96620 52198 96650 52250
rect 96650 52198 96676 52250
rect 96380 52196 96436 52198
rect 96460 52196 96516 52198
rect 96540 52196 96596 52198
rect 96620 52196 96676 52198
rect 81020 51706 81076 51708
rect 81100 51706 81156 51708
rect 81180 51706 81236 51708
rect 81260 51706 81316 51708
rect 81020 51654 81046 51706
rect 81046 51654 81076 51706
rect 81100 51654 81110 51706
rect 81110 51654 81156 51706
rect 81180 51654 81226 51706
rect 81226 51654 81236 51706
rect 81260 51654 81290 51706
rect 81290 51654 81316 51706
rect 81020 51652 81076 51654
rect 81100 51652 81156 51654
rect 81180 51652 81236 51654
rect 81260 51652 81316 51654
rect 111740 51706 111796 51708
rect 111820 51706 111876 51708
rect 111900 51706 111956 51708
rect 111980 51706 112036 51708
rect 111740 51654 111766 51706
rect 111766 51654 111796 51706
rect 111820 51654 111830 51706
rect 111830 51654 111876 51706
rect 111900 51654 111946 51706
rect 111946 51654 111956 51706
rect 111980 51654 112010 51706
rect 112010 51654 112036 51706
rect 111740 51652 111796 51654
rect 111820 51652 111876 51654
rect 111900 51652 111956 51654
rect 111980 51652 112036 51654
rect 96380 51162 96436 51164
rect 96460 51162 96516 51164
rect 96540 51162 96596 51164
rect 96620 51162 96676 51164
rect 96380 51110 96406 51162
rect 96406 51110 96436 51162
rect 96460 51110 96470 51162
rect 96470 51110 96516 51162
rect 96540 51110 96586 51162
rect 96586 51110 96596 51162
rect 96620 51110 96650 51162
rect 96650 51110 96676 51162
rect 96380 51108 96436 51110
rect 96460 51108 96516 51110
rect 96540 51108 96596 51110
rect 96620 51108 96676 51110
rect 81020 50618 81076 50620
rect 81100 50618 81156 50620
rect 81180 50618 81236 50620
rect 81260 50618 81316 50620
rect 81020 50566 81046 50618
rect 81046 50566 81076 50618
rect 81100 50566 81110 50618
rect 81110 50566 81156 50618
rect 81180 50566 81226 50618
rect 81226 50566 81236 50618
rect 81260 50566 81290 50618
rect 81290 50566 81316 50618
rect 81020 50564 81076 50566
rect 81100 50564 81156 50566
rect 81180 50564 81236 50566
rect 81260 50564 81316 50566
rect 111740 50618 111796 50620
rect 111820 50618 111876 50620
rect 111900 50618 111956 50620
rect 111980 50618 112036 50620
rect 111740 50566 111766 50618
rect 111766 50566 111796 50618
rect 111820 50566 111830 50618
rect 111830 50566 111876 50618
rect 111900 50566 111946 50618
rect 111946 50566 111956 50618
rect 111980 50566 112010 50618
rect 112010 50566 112036 50618
rect 111740 50564 111796 50566
rect 111820 50564 111876 50566
rect 111900 50564 111956 50566
rect 111980 50564 112036 50566
rect 96380 50074 96436 50076
rect 96460 50074 96516 50076
rect 96540 50074 96596 50076
rect 96620 50074 96676 50076
rect 96380 50022 96406 50074
rect 96406 50022 96436 50074
rect 96460 50022 96470 50074
rect 96470 50022 96516 50074
rect 96540 50022 96586 50074
rect 96586 50022 96596 50074
rect 96620 50022 96650 50074
rect 96650 50022 96676 50074
rect 96380 50020 96436 50022
rect 96460 50020 96516 50022
rect 96540 50020 96596 50022
rect 96620 50020 96676 50022
rect 81020 49530 81076 49532
rect 81100 49530 81156 49532
rect 81180 49530 81236 49532
rect 81260 49530 81316 49532
rect 81020 49478 81046 49530
rect 81046 49478 81076 49530
rect 81100 49478 81110 49530
rect 81110 49478 81156 49530
rect 81180 49478 81226 49530
rect 81226 49478 81236 49530
rect 81260 49478 81290 49530
rect 81290 49478 81316 49530
rect 81020 49476 81076 49478
rect 81100 49476 81156 49478
rect 81180 49476 81236 49478
rect 81260 49476 81316 49478
rect 111740 49530 111796 49532
rect 111820 49530 111876 49532
rect 111900 49530 111956 49532
rect 111980 49530 112036 49532
rect 111740 49478 111766 49530
rect 111766 49478 111796 49530
rect 111820 49478 111830 49530
rect 111830 49478 111876 49530
rect 111900 49478 111946 49530
rect 111946 49478 111956 49530
rect 111980 49478 112010 49530
rect 112010 49478 112036 49530
rect 111740 49476 111796 49478
rect 111820 49476 111876 49478
rect 111900 49476 111956 49478
rect 111980 49476 112036 49478
rect 96380 48986 96436 48988
rect 96460 48986 96516 48988
rect 96540 48986 96596 48988
rect 96620 48986 96676 48988
rect 96380 48934 96406 48986
rect 96406 48934 96436 48986
rect 96460 48934 96470 48986
rect 96470 48934 96516 48986
rect 96540 48934 96586 48986
rect 96586 48934 96596 48986
rect 96620 48934 96650 48986
rect 96650 48934 96676 48986
rect 96380 48932 96436 48934
rect 96460 48932 96516 48934
rect 96540 48932 96596 48934
rect 96620 48932 96676 48934
rect 81020 48442 81076 48444
rect 81100 48442 81156 48444
rect 81180 48442 81236 48444
rect 81260 48442 81316 48444
rect 81020 48390 81046 48442
rect 81046 48390 81076 48442
rect 81100 48390 81110 48442
rect 81110 48390 81156 48442
rect 81180 48390 81226 48442
rect 81226 48390 81236 48442
rect 81260 48390 81290 48442
rect 81290 48390 81316 48442
rect 81020 48388 81076 48390
rect 81100 48388 81156 48390
rect 81180 48388 81236 48390
rect 81260 48388 81316 48390
rect 111740 48442 111796 48444
rect 111820 48442 111876 48444
rect 111900 48442 111956 48444
rect 111980 48442 112036 48444
rect 111740 48390 111766 48442
rect 111766 48390 111796 48442
rect 111820 48390 111830 48442
rect 111830 48390 111876 48442
rect 111900 48390 111946 48442
rect 111946 48390 111956 48442
rect 111980 48390 112010 48442
rect 112010 48390 112036 48442
rect 111740 48388 111796 48390
rect 111820 48388 111876 48390
rect 111900 48388 111956 48390
rect 111980 48388 112036 48390
rect 96380 47898 96436 47900
rect 96460 47898 96516 47900
rect 96540 47898 96596 47900
rect 96620 47898 96676 47900
rect 96380 47846 96406 47898
rect 96406 47846 96436 47898
rect 96460 47846 96470 47898
rect 96470 47846 96516 47898
rect 96540 47846 96586 47898
rect 96586 47846 96596 47898
rect 96620 47846 96650 47898
rect 96650 47846 96676 47898
rect 96380 47844 96436 47846
rect 96460 47844 96516 47846
rect 96540 47844 96596 47846
rect 96620 47844 96676 47846
rect 81020 47354 81076 47356
rect 81100 47354 81156 47356
rect 81180 47354 81236 47356
rect 81260 47354 81316 47356
rect 81020 47302 81046 47354
rect 81046 47302 81076 47354
rect 81100 47302 81110 47354
rect 81110 47302 81156 47354
rect 81180 47302 81226 47354
rect 81226 47302 81236 47354
rect 81260 47302 81290 47354
rect 81290 47302 81316 47354
rect 81020 47300 81076 47302
rect 81100 47300 81156 47302
rect 81180 47300 81236 47302
rect 81260 47300 81316 47302
rect 111740 47354 111796 47356
rect 111820 47354 111876 47356
rect 111900 47354 111956 47356
rect 111980 47354 112036 47356
rect 111740 47302 111766 47354
rect 111766 47302 111796 47354
rect 111820 47302 111830 47354
rect 111830 47302 111876 47354
rect 111900 47302 111946 47354
rect 111946 47302 111956 47354
rect 111980 47302 112010 47354
rect 112010 47302 112036 47354
rect 111740 47300 111796 47302
rect 111820 47300 111876 47302
rect 111900 47300 111956 47302
rect 111980 47300 112036 47302
rect 96380 46810 96436 46812
rect 96460 46810 96516 46812
rect 96540 46810 96596 46812
rect 96620 46810 96676 46812
rect 96380 46758 96406 46810
rect 96406 46758 96436 46810
rect 96460 46758 96470 46810
rect 96470 46758 96516 46810
rect 96540 46758 96586 46810
rect 96586 46758 96596 46810
rect 96620 46758 96650 46810
rect 96650 46758 96676 46810
rect 96380 46756 96436 46758
rect 96460 46756 96516 46758
rect 96540 46756 96596 46758
rect 96620 46756 96676 46758
rect 81020 46266 81076 46268
rect 81100 46266 81156 46268
rect 81180 46266 81236 46268
rect 81260 46266 81316 46268
rect 81020 46214 81046 46266
rect 81046 46214 81076 46266
rect 81100 46214 81110 46266
rect 81110 46214 81156 46266
rect 81180 46214 81226 46266
rect 81226 46214 81236 46266
rect 81260 46214 81290 46266
rect 81290 46214 81316 46266
rect 81020 46212 81076 46214
rect 81100 46212 81156 46214
rect 81180 46212 81236 46214
rect 81260 46212 81316 46214
rect 111740 46266 111796 46268
rect 111820 46266 111876 46268
rect 111900 46266 111956 46268
rect 111980 46266 112036 46268
rect 111740 46214 111766 46266
rect 111766 46214 111796 46266
rect 111820 46214 111830 46266
rect 111830 46214 111876 46266
rect 111900 46214 111946 46266
rect 111946 46214 111956 46266
rect 111980 46214 112010 46266
rect 112010 46214 112036 46266
rect 111740 46212 111796 46214
rect 111820 46212 111876 46214
rect 111900 46212 111956 46214
rect 111980 46212 112036 46214
rect 96380 45722 96436 45724
rect 96460 45722 96516 45724
rect 96540 45722 96596 45724
rect 96620 45722 96676 45724
rect 96380 45670 96406 45722
rect 96406 45670 96436 45722
rect 96460 45670 96470 45722
rect 96470 45670 96516 45722
rect 96540 45670 96586 45722
rect 96586 45670 96596 45722
rect 96620 45670 96650 45722
rect 96650 45670 96676 45722
rect 96380 45668 96436 45670
rect 96460 45668 96516 45670
rect 96540 45668 96596 45670
rect 96620 45668 96676 45670
rect 81020 45178 81076 45180
rect 81100 45178 81156 45180
rect 81180 45178 81236 45180
rect 81260 45178 81316 45180
rect 81020 45126 81046 45178
rect 81046 45126 81076 45178
rect 81100 45126 81110 45178
rect 81110 45126 81156 45178
rect 81180 45126 81226 45178
rect 81226 45126 81236 45178
rect 81260 45126 81290 45178
rect 81290 45126 81316 45178
rect 81020 45124 81076 45126
rect 81100 45124 81156 45126
rect 81180 45124 81236 45126
rect 81260 45124 81316 45126
rect 111740 45178 111796 45180
rect 111820 45178 111876 45180
rect 111900 45178 111956 45180
rect 111980 45178 112036 45180
rect 111740 45126 111766 45178
rect 111766 45126 111796 45178
rect 111820 45126 111830 45178
rect 111830 45126 111876 45178
rect 111900 45126 111946 45178
rect 111946 45126 111956 45178
rect 111980 45126 112010 45178
rect 112010 45126 112036 45178
rect 111740 45124 111796 45126
rect 111820 45124 111876 45126
rect 111900 45124 111956 45126
rect 111980 45124 112036 45126
rect 96380 44634 96436 44636
rect 96460 44634 96516 44636
rect 96540 44634 96596 44636
rect 96620 44634 96676 44636
rect 96380 44582 96406 44634
rect 96406 44582 96436 44634
rect 96460 44582 96470 44634
rect 96470 44582 96516 44634
rect 96540 44582 96586 44634
rect 96586 44582 96596 44634
rect 96620 44582 96650 44634
rect 96650 44582 96676 44634
rect 96380 44580 96436 44582
rect 96460 44580 96516 44582
rect 96540 44580 96596 44582
rect 96620 44580 96676 44582
rect 81020 44090 81076 44092
rect 81100 44090 81156 44092
rect 81180 44090 81236 44092
rect 81260 44090 81316 44092
rect 81020 44038 81046 44090
rect 81046 44038 81076 44090
rect 81100 44038 81110 44090
rect 81110 44038 81156 44090
rect 81180 44038 81226 44090
rect 81226 44038 81236 44090
rect 81260 44038 81290 44090
rect 81290 44038 81316 44090
rect 81020 44036 81076 44038
rect 81100 44036 81156 44038
rect 81180 44036 81236 44038
rect 81260 44036 81316 44038
rect 111740 44090 111796 44092
rect 111820 44090 111876 44092
rect 111900 44090 111956 44092
rect 111980 44090 112036 44092
rect 111740 44038 111766 44090
rect 111766 44038 111796 44090
rect 111820 44038 111830 44090
rect 111830 44038 111876 44090
rect 111900 44038 111946 44090
rect 111946 44038 111956 44090
rect 111980 44038 112010 44090
rect 112010 44038 112036 44090
rect 111740 44036 111796 44038
rect 111820 44036 111876 44038
rect 111900 44036 111956 44038
rect 111980 44036 112036 44038
rect 96380 43546 96436 43548
rect 96460 43546 96516 43548
rect 96540 43546 96596 43548
rect 96620 43546 96676 43548
rect 96380 43494 96406 43546
rect 96406 43494 96436 43546
rect 96460 43494 96470 43546
rect 96470 43494 96516 43546
rect 96540 43494 96586 43546
rect 96586 43494 96596 43546
rect 96620 43494 96650 43546
rect 96650 43494 96676 43546
rect 96380 43492 96436 43494
rect 96460 43492 96516 43494
rect 96540 43492 96596 43494
rect 96620 43492 96676 43494
rect 81020 43002 81076 43004
rect 81100 43002 81156 43004
rect 81180 43002 81236 43004
rect 81260 43002 81316 43004
rect 81020 42950 81046 43002
rect 81046 42950 81076 43002
rect 81100 42950 81110 43002
rect 81110 42950 81156 43002
rect 81180 42950 81226 43002
rect 81226 42950 81236 43002
rect 81260 42950 81290 43002
rect 81290 42950 81316 43002
rect 81020 42948 81076 42950
rect 81100 42948 81156 42950
rect 81180 42948 81236 42950
rect 81260 42948 81316 42950
rect 111740 43002 111796 43004
rect 111820 43002 111876 43004
rect 111900 43002 111956 43004
rect 111980 43002 112036 43004
rect 111740 42950 111766 43002
rect 111766 42950 111796 43002
rect 111820 42950 111830 43002
rect 111830 42950 111876 43002
rect 111900 42950 111946 43002
rect 111946 42950 111956 43002
rect 111980 42950 112010 43002
rect 112010 42950 112036 43002
rect 111740 42948 111796 42950
rect 111820 42948 111876 42950
rect 111900 42948 111956 42950
rect 111980 42948 112036 42950
rect 96380 42458 96436 42460
rect 96460 42458 96516 42460
rect 96540 42458 96596 42460
rect 96620 42458 96676 42460
rect 96380 42406 96406 42458
rect 96406 42406 96436 42458
rect 96460 42406 96470 42458
rect 96470 42406 96516 42458
rect 96540 42406 96586 42458
rect 96586 42406 96596 42458
rect 96620 42406 96650 42458
rect 96650 42406 96676 42458
rect 96380 42404 96436 42406
rect 96460 42404 96516 42406
rect 96540 42404 96596 42406
rect 96620 42404 96676 42406
rect 81020 41914 81076 41916
rect 81100 41914 81156 41916
rect 81180 41914 81236 41916
rect 81260 41914 81316 41916
rect 81020 41862 81046 41914
rect 81046 41862 81076 41914
rect 81100 41862 81110 41914
rect 81110 41862 81156 41914
rect 81180 41862 81226 41914
rect 81226 41862 81236 41914
rect 81260 41862 81290 41914
rect 81290 41862 81316 41914
rect 81020 41860 81076 41862
rect 81100 41860 81156 41862
rect 81180 41860 81236 41862
rect 81260 41860 81316 41862
rect 111740 41914 111796 41916
rect 111820 41914 111876 41916
rect 111900 41914 111956 41916
rect 111980 41914 112036 41916
rect 111740 41862 111766 41914
rect 111766 41862 111796 41914
rect 111820 41862 111830 41914
rect 111830 41862 111876 41914
rect 111900 41862 111946 41914
rect 111946 41862 111956 41914
rect 111980 41862 112010 41914
rect 112010 41862 112036 41914
rect 111740 41860 111796 41862
rect 111820 41860 111876 41862
rect 111900 41860 111956 41862
rect 111980 41860 112036 41862
rect 96380 41370 96436 41372
rect 96460 41370 96516 41372
rect 96540 41370 96596 41372
rect 96620 41370 96676 41372
rect 96380 41318 96406 41370
rect 96406 41318 96436 41370
rect 96460 41318 96470 41370
rect 96470 41318 96516 41370
rect 96540 41318 96586 41370
rect 96586 41318 96596 41370
rect 96620 41318 96650 41370
rect 96650 41318 96676 41370
rect 96380 41316 96436 41318
rect 96460 41316 96516 41318
rect 96540 41316 96596 41318
rect 96620 41316 96676 41318
rect 81020 40826 81076 40828
rect 81100 40826 81156 40828
rect 81180 40826 81236 40828
rect 81260 40826 81316 40828
rect 81020 40774 81046 40826
rect 81046 40774 81076 40826
rect 81100 40774 81110 40826
rect 81110 40774 81156 40826
rect 81180 40774 81226 40826
rect 81226 40774 81236 40826
rect 81260 40774 81290 40826
rect 81290 40774 81316 40826
rect 81020 40772 81076 40774
rect 81100 40772 81156 40774
rect 81180 40772 81236 40774
rect 81260 40772 81316 40774
rect 111740 40826 111796 40828
rect 111820 40826 111876 40828
rect 111900 40826 111956 40828
rect 111980 40826 112036 40828
rect 111740 40774 111766 40826
rect 111766 40774 111796 40826
rect 111820 40774 111830 40826
rect 111830 40774 111876 40826
rect 111900 40774 111946 40826
rect 111946 40774 111956 40826
rect 111980 40774 112010 40826
rect 112010 40774 112036 40826
rect 111740 40772 111796 40774
rect 111820 40772 111876 40774
rect 111900 40772 111956 40774
rect 111980 40772 112036 40774
rect 96380 40282 96436 40284
rect 96460 40282 96516 40284
rect 96540 40282 96596 40284
rect 96620 40282 96676 40284
rect 96380 40230 96406 40282
rect 96406 40230 96436 40282
rect 96460 40230 96470 40282
rect 96470 40230 96516 40282
rect 96540 40230 96586 40282
rect 96586 40230 96596 40282
rect 96620 40230 96650 40282
rect 96650 40230 96676 40282
rect 96380 40228 96436 40230
rect 96460 40228 96516 40230
rect 96540 40228 96596 40230
rect 96620 40228 96676 40230
rect 81020 39738 81076 39740
rect 81100 39738 81156 39740
rect 81180 39738 81236 39740
rect 81260 39738 81316 39740
rect 81020 39686 81046 39738
rect 81046 39686 81076 39738
rect 81100 39686 81110 39738
rect 81110 39686 81156 39738
rect 81180 39686 81226 39738
rect 81226 39686 81236 39738
rect 81260 39686 81290 39738
rect 81290 39686 81316 39738
rect 81020 39684 81076 39686
rect 81100 39684 81156 39686
rect 81180 39684 81236 39686
rect 81260 39684 81316 39686
rect 111740 39738 111796 39740
rect 111820 39738 111876 39740
rect 111900 39738 111956 39740
rect 111980 39738 112036 39740
rect 111740 39686 111766 39738
rect 111766 39686 111796 39738
rect 111820 39686 111830 39738
rect 111830 39686 111876 39738
rect 111900 39686 111946 39738
rect 111946 39686 111956 39738
rect 111980 39686 112010 39738
rect 112010 39686 112036 39738
rect 111740 39684 111796 39686
rect 111820 39684 111876 39686
rect 111900 39684 111956 39686
rect 111980 39684 112036 39686
rect 96380 39194 96436 39196
rect 96460 39194 96516 39196
rect 96540 39194 96596 39196
rect 96620 39194 96676 39196
rect 96380 39142 96406 39194
rect 96406 39142 96436 39194
rect 96460 39142 96470 39194
rect 96470 39142 96516 39194
rect 96540 39142 96586 39194
rect 96586 39142 96596 39194
rect 96620 39142 96650 39194
rect 96650 39142 96676 39194
rect 96380 39140 96436 39142
rect 96460 39140 96516 39142
rect 96540 39140 96596 39142
rect 96620 39140 96676 39142
rect 81020 38650 81076 38652
rect 81100 38650 81156 38652
rect 81180 38650 81236 38652
rect 81260 38650 81316 38652
rect 81020 38598 81046 38650
rect 81046 38598 81076 38650
rect 81100 38598 81110 38650
rect 81110 38598 81156 38650
rect 81180 38598 81226 38650
rect 81226 38598 81236 38650
rect 81260 38598 81290 38650
rect 81290 38598 81316 38650
rect 81020 38596 81076 38598
rect 81100 38596 81156 38598
rect 81180 38596 81236 38598
rect 81260 38596 81316 38598
rect 111740 38650 111796 38652
rect 111820 38650 111876 38652
rect 111900 38650 111956 38652
rect 111980 38650 112036 38652
rect 111740 38598 111766 38650
rect 111766 38598 111796 38650
rect 111820 38598 111830 38650
rect 111830 38598 111876 38650
rect 111900 38598 111946 38650
rect 111946 38598 111956 38650
rect 111980 38598 112010 38650
rect 112010 38598 112036 38650
rect 111740 38596 111796 38598
rect 111820 38596 111876 38598
rect 111900 38596 111956 38598
rect 111980 38596 112036 38598
rect 96380 38106 96436 38108
rect 96460 38106 96516 38108
rect 96540 38106 96596 38108
rect 96620 38106 96676 38108
rect 96380 38054 96406 38106
rect 96406 38054 96436 38106
rect 96460 38054 96470 38106
rect 96470 38054 96516 38106
rect 96540 38054 96586 38106
rect 96586 38054 96596 38106
rect 96620 38054 96650 38106
rect 96650 38054 96676 38106
rect 96380 38052 96436 38054
rect 96460 38052 96516 38054
rect 96540 38052 96596 38054
rect 96620 38052 96676 38054
rect 81020 37562 81076 37564
rect 81100 37562 81156 37564
rect 81180 37562 81236 37564
rect 81260 37562 81316 37564
rect 81020 37510 81046 37562
rect 81046 37510 81076 37562
rect 81100 37510 81110 37562
rect 81110 37510 81156 37562
rect 81180 37510 81226 37562
rect 81226 37510 81236 37562
rect 81260 37510 81290 37562
rect 81290 37510 81316 37562
rect 81020 37508 81076 37510
rect 81100 37508 81156 37510
rect 81180 37508 81236 37510
rect 81260 37508 81316 37510
rect 111740 37562 111796 37564
rect 111820 37562 111876 37564
rect 111900 37562 111956 37564
rect 111980 37562 112036 37564
rect 111740 37510 111766 37562
rect 111766 37510 111796 37562
rect 111820 37510 111830 37562
rect 111830 37510 111876 37562
rect 111900 37510 111946 37562
rect 111946 37510 111956 37562
rect 111980 37510 112010 37562
rect 112010 37510 112036 37562
rect 111740 37508 111796 37510
rect 111820 37508 111876 37510
rect 111900 37508 111956 37510
rect 111980 37508 112036 37510
rect 96380 37018 96436 37020
rect 96460 37018 96516 37020
rect 96540 37018 96596 37020
rect 96620 37018 96676 37020
rect 96380 36966 96406 37018
rect 96406 36966 96436 37018
rect 96460 36966 96470 37018
rect 96470 36966 96516 37018
rect 96540 36966 96586 37018
rect 96586 36966 96596 37018
rect 96620 36966 96650 37018
rect 96650 36966 96676 37018
rect 96380 36964 96436 36966
rect 96460 36964 96516 36966
rect 96540 36964 96596 36966
rect 96620 36964 96676 36966
rect 81020 36474 81076 36476
rect 81100 36474 81156 36476
rect 81180 36474 81236 36476
rect 81260 36474 81316 36476
rect 81020 36422 81046 36474
rect 81046 36422 81076 36474
rect 81100 36422 81110 36474
rect 81110 36422 81156 36474
rect 81180 36422 81226 36474
rect 81226 36422 81236 36474
rect 81260 36422 81290 36474
rect 81290 36422 81316 36474
rect 81020 36420 81076 36422
rect 81100 36420 81156 36422
rect 81180 36420 81236 36422
rect 81260 36420 81316 36422
rect 111740 36474 111796 36476
rect 111820 36474 111876 36476
rect 111900 36474 111956 36476
rect 111980 36474 112036 36476
rect 111740 36422 111766 36474
rect 111766 36422 111796 36474
rect 111820 36422 111830 36474
rect 111830 36422 111876 36474
rect 111900 36422 111946 36474
rect 111946 36422 111956 36474
rect 111980 36422 112010 36474
rect 112010 36422 112036 36474
rect 111740 36420 111796 36422
rect 111820 36420 111876 36422
rect 111900 36420 111956 36422
rect 111980 36420 112036 36422
rect 96380 35930 96436 35932
rect 96460 35930 96516 35932
rect 96540 35930 96596 35932
rect 96620 35930 96676 35932
rect 96380 35878 96406 35930
rect 96406 35878 96436 35930
rect 96460 35878 96470 35930
rect 96470 35878 96516 35930
rect 96540 35878 96586 35930
rect 96586 35878 96596 35930
rect 96620 35878 96650 35930
rect 96650 35878 96676 35930
rect 96380 35876 96436 35878
rect 96460 35876 96516 35878
rect 96540 35876 96596 35878
rect 96620 35876 96676 35878
rect 81020 35386 81076 35388
rect 81100 35386 81156 35388
rect 81180 35386 81236 35388
rect 81260 35386 81316 35388
rect 81020 35334 81046 35386
rect 81046 35334 81076 35386
rect 81100 35334 81110 35386
rect 81110 35334 81156 35386
rect 81180 35334 81226 35386
rect 81226 35334 81236 35386
rect 81260 35334 81290 35386
rect 81290 35334 81316 35386
rect 81020 35332 81076 35334
rect 81100 35332 81156 35334
rect 81180 35332 81236 35334
rect 81260 35332 81316 35334
rect 111740 35386 111796 35388
rect 111820 35386 111876 35388
rect 111900 35386 111956 35388
rect 111980 35386 112036 35388
rect 111740 35334 111766 35386
rect 111766 35334 111796 35386
rect 111820 35334 111830 35386
rect 111830 35334 111876 35386
rect 111900 35334 111946 35386
rect 111946 35334 111956 35386
rect 111980 35334 112010 35386
rect 112010 35334 112036 35386
rect 111740 35332 111796 35334
rect 111820 35332 111876 35334
rect 111900 35332 111956 35334
rect 111980 35332 112036 35334
rect 96380 34842 96436 34844
rect 96460 34842 96516 34844
rect 96540 34842 96596 34844
rect 96620 34842 96676 34844
rect 96380 34790 96406 34842
rect 96406 34790 96436 34842
rect 96460 34790 96470 34842
rect 96470 34790 96516 34842
rect 96540 34790 96586 34842
rect 96586 34790 96596 34842
rect 96620 34790 96650 34842
rect 96650 34790 96676 34842
rect 96380 34788 96436 34790
rect 96460 34788 96516 34790
rect 96540 34788 96596 34790
rect 96620 34788 96676 34790
rect 81020 34298 81076 34300
rect 81100 34298 81156 34300
rect 81180 34298 81236 34300
rect 81260 34298 81316 34300
rect 81020 34246 81046 34298
rect 81046 34246 81076 34298
rect 81100 34246 81110 34298
rect 81110 34246 81156 34298
rect 81180 34246 81226 34298
rect 81226 34246 81236 34298
rect 81260 34246 81290 34298
rect 81290 34246 81316 34298
rect 81020 34244 81076 34246
rect 81100 34244 81156 34246
rect 81180 34244 81236 34246
rect 81260 34244 81316 34246
rect 111740 34298 111796 34300
rect 111820 34298 111876 34300
rect 111900 34298 111956 34300
rect 111980 34298 112036 34300
rect 111740 34246 111766 34298
rect 111766 34246 111796 34298
rect 111820 34246 111830 34298
rect 111830 34246 111876 34298
rect 111900 34246 111946 34298
rect 111946 34246 111956 34298
rect 111980 34246 112010 34298
rect 112010 34246 112036 34298
rect 111740 34244 111796 34246
rect 111820 34244 111876 34246
rect 111900 34244 111956 34246
rect 111980 34244 112036 34246
rect 96380 33754 96436 33756
rect 96460 33754 96516 33756
rect 96540 33754 96596 33756
rect 96620 33754 96676 33756
rect 96380 33702 96406 33754
rect 96406 33702 96436 33754
rect 96460 33702 96470 33754
rect 96470 33702 96516 33754
rect 96540 33702 96586 33754
rect 96586 33702 96596 33754
rect 96620 33702 96650 33754
rect 96650 33702 96676 33754
rect 96380 33700 96436 33702
rect 96460 33700 96516 33702
rect 96540 33700 96596 33702
rect 96620 33700 96676 33702
rect 81020 33210 81076 33212
rect 81100 33210 81156 33212
rect 81180 33210 81236 33212
rect 81260 33210 81316 33212
rect 81020 33158 81046 33210
rect 81046 33158 81076 33210
rect 81100 33158 81110 33210
rect 81110 33158 81156 33210
rect 81180 33158 81226 33210
rect 81226 33158 81236 33210
rect 81260 33158 81290 33210
rect 81290 33158 81316 33210
rect 81020 33156 81076 33158
rect 81100 33156 81156 33158
rect 81180 33156 81236 33158
rect 81260 33156 81316 33158
rect 111740 33210 111796 33212
rect 111820 33210 111876 33212
rect 111900 33210 111956 33212
rect 111980 33210 112036 33212
rect 111740 33158 111766 33210
rect 111766 33158 111796 33210
rect 111820 33158 111830 33210
rect 111830 33158 111876 33210
rect 111900 33158 111946 33210
rect 111946 33158 111956 33210
rect 111980 33158 112010 33210
rect 112010 33158 112036 33210
rect 111740 33156 111796 33158
rect 111820 33156 111876 33158
rect 111900 33156 111956 33158
rect 111980 33156 112036 33158
rect 96380 32666 96436 32668
rect 96460 32666 96516 32668
rect 96540 32666 96596 32668
rect 96620 32666 96676 32668
rect 96380 32614 96406 32666
rect 96406 32614 96436 32666
rect 96460 32614 96470 32666
rect 96470 32614 96516 32666
rect 96540 32614 96586 32666
rect 96586 32614 96596 32666
rect 96620 32614 96650 32666
rect 96650 32614 96676 32666
rect 96380 32612 96436 32614
rect 96460 32612 96516 32614
rect 96540 32612 96596 32614
rect 96620 32612 96676 32614
rect 81020 32122 81076 32124
rect 81100 32122 81156 32124
rect 81180 32122 81236 32124
rect 81260 32122 81316 32124
rect 81020 32070 81046 32122
rect 81046 32070 81076 32122
rect 81100 32070 81110 32122
rect 81110 32070 81156 32122
rect 81180 32070 81226 32122
rect 81226 32070 81236 32122
rect 81260 32070 81290 32122
rect 81290 32070 81316 32122
rect 81020 32068 81076 32070
rect 81100 32068 81156 32070
rect 81180 32068 81236 32070
rect 81260 32068 81316 32070
rect 111740 32122 111796 32124
rect 111820 32122 111876 32124
rect 111900 32122 111956 32124
rect 111980 32122 112036 32124
rect 111740 32070 111766 32122
rect 111766 32070 111796 32122
rect 111820 32070 111830 32122
rect 111830 32070 111876 32122
rect 111900 32070 111946 32122
rect 111946 32070 111956 32122
rect 111980 32070 112010 32122
rect 112010 32070 112036 32122
rect 111740 32068 111796 32070
rect 111820 32068 111876 32070
rect 111900 32068 111956 32070
rect 111980 32068 112036 32070
rect 96380 31578 96436 31580
rect 96460 31578 96516 31580
rect 96540 31578 96596 31580
rect 96620 31578 96676 31580
rect 96380 31526 96406 31578
rect 96406 31526 96436 31578
rect 96460 31526 96470 31578
rect 96470 31526 96516 31578
rect 96540 31526 96586 31578
rect 96586 31526 96596 31578
rect 96620 31526 96650 31578
rect 96650 31526 96676 31578
rect 96380 31524 96436 31526
rect 96460 31524 96516 31526
rect 96540 31524 96596 31526
rect 96620 31524 96676 31526
rect 81020 31034 81076 31036
rect 81100 31034 81156 31036
rect 81180 31034 81236 31036
rect 81260 31034 81316 31036
rect 81020 30982 81046 31034
rect 81046 30982 81076 31034
rect 81100 30982 81110 31034
rect 81110 30982 81156 31034
rect 81180 30982 81226 31034
rect 81226 30982 81236 31034
rect 81260 30982 81290 31034
rect 81290 30982 81316 31034
rect 81020 30980 81076 30982
rect 81100 30980 81156 30982
rect 81180 30980 81236 30982
rect 81260 30980 81316 30982
rect 111740 31034 111796 31036
rect 111820 31034 111876 31036
rect 111900 31034 111956 31036
rect 111980 31034 112036 31036
rect 111740 30982 111766 31034
rect 111766 30982 111796 31034
rect 111820 30982 111830 31034
rect 111830 30982 111876 31034
rect 111900 30982 111946 31034
rect 111946 30982 111956 31034
rect 111980 30982 112010 31034
rect 112010 30982 112036 31034
rect 111740 30980 111796 30982
rect 111820 30980 111876 30982
rect 111900 30980 111956 30982
rect 111980 30980 112036 30982
rect 96380 30490 96436 30492
rect 96460 30490 96516 30492
rect 96540 30490 96596 30492
rect 96620 30490 96676 30492
rect 96380 30438 96406 30490
rect 96406 30438 96436 30490
rect 96460 30438 96470 30490
rect 96470 30438 96516 30490
rect 96540 30438 96586 30490
rect 96586 30438 96596 30490
rect 96620 30438 96650 30490
rect 96650 30438 96676 30490
rect 96380 30436 96436 30438
rect 96460 30436 96516 30438
rect 96540 30436 96596 30438
rect 96620 30436 96676 30438
rect 81020 29946 81076 29948
rect 81100 29946 81156 29948
rect 81180 29946 81236 29948
rect 81260 29946 81316 29948
rect 81020 29894 81046 29946
rect 81046 29894 81076 29946
rect 81100 29894 81110 29946
rect 81110 29894 81156 29946
rect 81180 29894 81226 29946
rect 81226 29894 81236 29946
rect 81260 29894 81290 29946
rect 81290 29894 81316 29946
rect 81020 29892 81076 29894
rect 81100 29892 81156 29894
rect 81180 29892 81236 29894
rect 81260 29892 81316 29894
rect 111740 29946 111796 29948
rect 111820 29946 111876 29948
rect 111900 29946 111956 29948
rect 111980 29946 112036 29948
rect 111740 29894 111766 29946
rect 111766 29894 111796 29946
rect 111820 29894 111830 29946
rect 111830 29894 111876 29946
rect 111900 29894 111946 29946
rect 111946 29894 111956 29946
rect 111980 29894 112010 29946
rect 112010 29894 112036 29946
rect 111740 29892 111796 29894
rect 111820 29892 111876 29894
rect 111900 29892 111956 29894
rect 111980 29892 112036 29894
rect 96380 29402 96436 29404
rect 96460 29402 96516 29404
rect 96540 29402 96596 29404
rect 96620 29402 96676 29404
rect 96380 29350 96406 29402
rect 96406 29350 96436 29402
rect 96460 29350 96470 29402
rect 96470 29350 96516 29402
rect 96540 29350 96586 29402
rect 96586 29350 96596 29402
rect 96620 29350 96650 29402
rect 96650 29350 96676 29402
rect 96380 29348 96436 29350
rect 96460 29348 96516 29350
rect 96540 29348 96596 29350
rect 96620 29348 96676 29350
rect 81020 28858 81076 28860
rect 81100 28858 81156 28860
rect 81180 28858 81236 28860
rect 81260 28858 81316 28860
rect 81020 28806 81046 28858
rect 81046 28806 81076 28858
rect 81100 28806 81110 28858
rect 81110 28806 81156 28858
rect 81180 28806 81226 28858
rect 81226 28806 81236 28858
rect 81260 28806 81290 28858
rect 81290 28806 81316 28858
rect 81020 28804 81076 28806
rect 81100 28804 81156 28806
rect 81180 28804 81236 28806
rect 81260 28804 81316 28806
rect 111740 28858 111796 28860
rect 111820 28858 111876 28860
rect 111900 28858 111956 28860
rect 111980 28858 112036 28860
rect 111740 28806 111766 28858
rect 111766 28806 111796 28858
rect 111820 28806 111830 28858
rect 111830 28806 111876 28858
rect 111900 28806 111946 28858
rect 111946 28806 111956 28858
rect 111980 28806 112010 28858
rect 112010 28806 112036 28858
rect 111740 28804 111796 28806
rect 111820 28804 111876 28806
rect 111900 28804 111956 28806
rect 111980 28804 112036 28806
rect 96380 28314 96436 28316
rect 96460 28314 96516 28316
rect 96540 28314 96596 28316
rect 96620 28314 96676 28316
rect 96380 28262 96406 28314
rect 96406 28262 96436 28314
rect 96460 28262 96470 28314
rect 96470 28262 96516 28314
rect 96540 28262 96586 28314
rect 96586 28262 96596 28314
rect 96620 28262 96650 28314
rect 96650 28262 96676 28314
rect 96380 28260 96436 28262
rect 96460 28260 96516 28262
rect 96540 28260 96596 28262
rect 96620 28260 96676 28262
rect 81020 27770 81076 27772
rect 81100 27770 81156 27772
rect 81180 27770 81236 27772
rect 81260 27770 81316 27772
rect 81020 27718 81046 27770
rect 81046 27718 81076 27770
rect 81100 27718 81110 27770
rect 81110 27718 81156 27770
rect 81180 27718 81226 27770
rect 81226 27718 81236 27770
rect 81260 27718 81290 27770
rect 81290 27718 81316 27770
rect 81020 27716 81076 27718
rect 81100 27716 81156 27718
rect 81180 27716 81236 27718
rect 81260 27716 81316 27718
rect 111740 27770 111796 27772
rect 111820 27770 111876 27772
rect 111900 27770 111956 27772
rect 111980 27770 112036 27772
rect 111740 27718 111766 27770
rect 111766 27718 111796 27770
rect 111820 27718 111830 27770
rect 111830 27718 111876 27770
rect 111900 27718 111946 27770
rect 111946 27718 111956 27770
rect 111980 27718 112010 27770
rect 112010 27718 112036 27770
rect 111740 27716 111796 27718
rect 111820 27716 111876 27718
rect 111900 27716 111956 27718
rect 111980 27716 112036 27718
rect 96380 27226 96436 27228
rect 96460 27226 96516 27228
rect 96540 27226 96596 27228
rect 96620 27226 96676 27228
rect 96380 27174 96406 27226
rect 96406 27174 96436 27226
rect 96460 27174 96470 27226
rect 96470 27174 96516 27226
rect 96540 27174 96586 27226
rect 96586 27174 96596 27226
rect 96620 27174 96650 27226
rect 96650 27174 96676 27226
rect 96380 27172 96436 27174
rect 96460 27172 96516 27174
rect 96540 27172 96596 27174
rect 96620 27172 96676 27174
rect 81020 26682 81076 26684
rect 81100 26682 81156 26684
rect 81180 26682 81236 26684
rect 81260 26682 81316 26684
rect 81020 26630 81046 26682
rect 81046 26630 81076 26682
rect 81100 26630 81110 26682
rect 81110 26630 81156 26682
rect 81180 26630 81226 26682
rect 81226 26630 81236 26682
rect 81260 26630 81290 26682
rect 81290 26630 81316 26682
rect 81020 26628 81076 26630
rect 81100 26628 81156 26630
rect 81180 26628 81236 26630
rect 81260 26628 81316 26630
rect 111740 26682 111796 26684
rect 111820 26682 111876 26684
rect 111900 26682 111956 26684
rect 111980 26682 112036 26684
rect 111740 26630 111766 26682
rect 111766 26630 111796 26682
rect 111820 26630 111830 26682
rect 111830 26630 111876 26682
rect 111900 26630 111946 26682
rect 111946 26630 111956 26682
rect 111980 26630 112010 26682
rect 112010 26630 112036 26682
rect 111740 26628 111796 26630
rect 111820 26628 111876 26630
rect 111900 26628 111956 26630
rect 111980 26628 112036 26630
rect 96380 26138 96436 26140
rect 96460 26138 96516 26140
rect 96540 26138 96596 26140
rect 96620 26138 96676 26140
rect 96380 26086 96406 26138
rect 96406 26086 96436 26138
rect 96460 26086 96470 26138
rect 96470 26086 96516 26138
rect 96540 26086 96586 26138
rect 96586 26086 96596 26138
rect 96620 26086 96650 26138
rect 96650 26086 96676 26138
rect 96380 26084 96436 26086
rect 96460 26084 96516 26086
rect 96540 26084 96596 26086
rect 96620 26084 96676 26086
rect 81020 25594 81076 25596
rect 81100 25594 81156 25596
rect 81180 25594 81236 25596
rect 81260 25594 81316 25596
rect 81020 25542 81046 25594
rect 81046 25542 81076 25594
rect 81100 25542 81110 25594
rect 81110 25542 81156 25594
rect 81180 25542 81226 25594
rect 81226 25542 81236 25594
rect 81260 25542 81290 25594
rect 81290 25542 81316 25594
rect 81020 25540 81076 25542
rect 81100 25540 81156 25542
rect 81180 25540 81236 25542
rect 81260 25540 81316 25542
rect 111740 25594 111796 25596
rect 111820 25594 111876 25596
rect 111900 25594 111956 25596
rect 111980 25594 112036 25596
rect 111740 25542 111766 25594
rect 111766 25542 111796 25594
rect 111820 25542 111830 25594
rect 111830 25542 111876 25594
rect 111900 25542 111946 25594
rect 111946 25542 111956 25594
rect 111980 25542 112010 25594
rect 112010 25542 112036 25594
rect 111740 25540 111796 25542
rect 111820 25540 111876 25542
rect 111900 25540 111956 25542
rect 111980 25540 112036 25542
rect 96380 25050 96436 25052
rect 96460 25050 96516 25052
rect 96540 25050 96596 25052
rect 96620 25050 96676 25052
rect 96380 24998 96406 25050
rect 96406 24998 96436 25050
rect 96460 24998 96470 25050
rect 96470 24998 96516 25050
rect 96540 24998 96586 25050
rect 96586 24998 96596 25050
rect 96620 24998 96650 25050
rect 96650 24998 96676 25050
rect 96380 24996 96436 24998
rect 96460 24996 96516 24998
rect 96540 24996 96596 24998
rect 96620 24996 96676 24998
rect 81020 24506 81076 24508
rect 81100 24506 81156 24508
rect 81180 24506 81236 24508
rect 81260 24506 81316 24508
rect 81020 24454 81046 24506
rect 81046 24454 81076 24506
rect 81100 24454 81110 24506
rect 81110 24454 81156 24506
rect 81180 24454 81226 24506
rect 81226 24454 81236 24506
rect 81260 24454 81290 24506
rect 81290 24454 81316 24506
rect 81020 24452 81076 24454
rect 81100 24452 81156 24454
rect 81180 24452 81236 24454
rect 81260 24452 81316 24454
rect 111740 24506 111796 24508
rect 111820 24506 111876 24508
rect 111900 24506 111956 24508
rect 111980 24506 112036 24508
rect 111740 24454 111766 24506
rect 111766 24454 111796 24506
rect 111820 24454 111830 24506
rect 111830 24454 111876 24506
rect 111900 24454 111946 24506
rect 111946 24454 111956 24506
rect 111980 24454 112010 24506
rect 112010 24454 112036 24506
rect 111740 24452 111796 24454
rect 111820 24452 111876 24454
rect 111900 24452 111956 24454
rect 111980 24452 112036 24454
rect 96380 23962 96436 23964
rect 96460 23962 96516 23964
rect 96540 23962 96596 23964
rect 96620 23962 96676 23964
rect 96380 23910 96406 23962
rect 96406 23910 96436 23962
rect 96460 23910 96470 23962
rect 96470 23910 96516 23962
rect 96540 23910 96586 23962
rect 96586 23910 96596 23962
rect 96620 23910 96650 23962
rect 96650 23910 96676 23962
rect 96380 23908 96436 23910
rect 96460 23908 96516 23910
rect 96540 23908 96596 23910
rect 96620 23908 96676 23910
rect 81020 23418 81076 23420
rect 81100 23418 81156 23420
rect 81180 23418 81236 23420
rect 81260 23418 81316 23420
rect 81020 23366 81046 23418
rect 81046 23366 81076 23418
rect 81100 23366 81110 23418
rect 81110 23366 81156 23418
rect 81180 23366 81226 23418
rect 81226 23366 81236 23418
rect 81260 23366 81290 23418
rect 81290 23366 81316 23418
rect 81020 23364 81076 23366
rect 81100 23364 81156 23366
rect 81180 23364 81236 23366
rect 81260 23364 81316 23366
rect 111740 23418 111796 23420
rect 111820 23418 111876 23420
rect 111900 23418 111956 23420
rect 111980 23418 112036 23420
rect 111740 23366 111766 23418
rect 111766 23366 111796 23418
rect 111820 23366 111830 23418
rect 111830 23366 111876 23418
rect 111900 23366 111946 23418
rect 111946 23366 111956 23418
rect 111980 23366 112010 23418
rect 112010 23366 112036 23418
rect 111740 23364 111796 23366
rect 111820 23364 111876 23366
rect 111900 23364 111956 23366
rect 111980 23364 112036 23366
rect 96380 22874 96436 22876
rect 96460 22874 96516 22876
rect 96540 22874 96596 22876
rect 96620 22874 96676 22876
rect 96380 22822 96406 22874
rect 96406 22822 96436 22874
rect 96460 22822 96470 22874
rect 96470 22822 96516 22874
rect 96540 22822 96586 22874
rect 96586 22822 96596 22874
rect 96620 22822 96650 22874
rect 96650 22822 96676 22874
rect 96380 22820 96436 22822
rect 96460 22820 96516 22822
rect 96540 22820 96596 22822
rect 96620 22820 96676 22822
rect 81020 22330 81076 22332
rect 81100 22330 81156 22332
rect 81180 22330 81236 22332
rect 81260 22330 81316 22332
rect 81020 22278 81046 22330
rect 81046 22278 81076 22330
rect 81100 22278 81110 22330
rect 81110 22278 81156 22330
rect 81180 22278 81226 22330
rect 81226 22278 81236 22330
rect 81260 22278 81290 22330
rect 81290 22278 81316 22330
rect 81020 22276 81076 22278
rect 81100 22276 81156 22278
rect 81180 22276 81236 22278
rect 81260 22276 81316 22278
rect 111740 22330 111796 22332
rect 111820 22330 111876 22332
rect 111900 22330 111956 22332
rect 111980 22330 112036 22332
rect 111740 22278 111766 22330
rect 111766 22278 111796 22330
rect 111820 22278 111830 22330
rect 111830 22278 111876 22330
rect 111900 22278 111946 22330
rect 111946 22278 111956 22330
rect 111980 22278 112010 22330
rect 112010 22278 112036 22330
rect 111740 22276 111796 22278
rect 111820 22276 111876 22278
rect 111900 22276 111956 22278
rect 111980 22276 112036 22278
rect 96380 21786 96436 21788
rect 96460 21786 96516 21788
rect 96540 21786 96596 21788
rect 96620 21786 96676 21788
rect 96380 21734 96406 21786
rect 96406 21734 96436 21786
rect 96460 21734 96470 21786
rect 96470 21734 96516 21786
rect 96540 21734 96586 21786
rect 96586 21734 96596 21786
rect 96620 21734 96650 21786
rect 96650 21734 96676 21786
rect 96380 21732 96436 21734
rect 96460 21732 96516 21734
rect 96540 21732 96596 21734
rect 96620 21732 96676 21734
rect 81020 21242 81076 21244
rect 81100 21242 81156 21244
rect 81180 21242 81236 21244
rect 81260 21242 81316 21244
rect 81020 21190 81046 21242
rect 81046 21190 81076 21242
rect 81100 21190 81110 21242
rect 81110 21190 81156 21242
rect 81180 21190 81226 21242
rect 81226 21190 81236 21242
rect 81260 21190 81290 21242
rect 81290 21190 81316 21242
rect 81020 21188 81076 21190
rect 81100 21188 81156 21190
rect 81180 21188 81236 21190
rect 81260 21188 81316 21190
rect 111740 21242 111796 21244
rect 111820 21242 111876 21244
rect 111900 21242 111956 21244
rect 111980 21242 112036 21244
rect 111740 21190 111766 21242
rect 111766 21190 111796 21242
rect 111820 21190 111830 21242
rect 111830 21190 111876 21242
rect 111900 21190 111946 21242
rect 111946 21190 111956 21242
rect 111980 21190 112010 21242
rect 112010 21190 112036 21242
rect 111740 21188 111796 21190
rect 111820 21188 111876 21190
rect 111900 21188 111956 21190
rect 111980 21188 112036 21190
rect 96380 20698 96436 20700
rect 96460 20698 96516 20700
rect 96540 20698 96596 20700
rect 96620 20698 96676 20700
rect 96380 20646 96406 20698
rect 96406 20646 96436 20698
rect 96460 20646 96470 20698
rect 96470 20646 96516 20698
rect 96540 20646 96586 20698
rect 96586 20646 96596 20698
rect 96620 20646 96650 20698
rect 96650 20646 96676 20698
rect 96380 20644 96436 20646
rect 96460 20644 96516 20646
rect 96540 20644 96596 20646
rect 96620 20644 96676 20646
rect 69386 4664 69442 4720
rect 69754 3440 69810 3496
rect 81020 20154 81076 20156
rect 81100 20154 81156 20156
rect 81180 20154 81236 20156
rect 81260 20154 81316 20156
rect 81020 20102 81046 20154
rect 81046 20102 81076 20154
rect 81100 20102 81110 20154
rect 81110 20102 81156 20154
rect 81180 20102 81226 20154
rect 81226 20102 81236 20154
rect 81260 20102 81290 20154
rect 81290 20102 81316 20154
rect 81020 20100 81076 20102
rect 81100 20100 81156 20102
rect 81180 20100 81236 20102
rect 81260 20100 81316 20102
rect 111740 20154 111796 20156
rect 111820 20154 111876 20156
rect 111900 20154 111956 20156
rect 111980 20154 112036 20156
rect 111740 20102 111766 20154
rect 111766 20102 111796 20154
rect 111820 20102 111830 20154
rect 111830 20102 111876 20154
rect 111900 20102 111946 20154
rect 111946 20102 111956 20154
rect 111980 20102 112010 20154
rect 112010 20102 112036 20154
rect 111740 20100 111796 20102
rect 111820 20100 111876 20102
rect 111900 20100 111956 20102
rect 111980 20100 112036 20102
rect 127100 116442 127156 116444
rect 127180 116442 127236 116444
rect 127260 116442 127316 116444
rect 127340 116442 127396 116444
rect 127100 116390 127126 116442
rect 127126 116390 127156 116442
rect 127180 116390 127190 116442
rect 127190 116390 127236 116442
rect 127260 116390 127306 116442
rect 127306 116390 127316 116442
rect 127340 116390 127370 116442
rect 127370 116390 127396 116442
rect 127100 116388 127156 116390
rect 127180 116388 127236 116390
rect 127260 116388 127316 116390
rect 127340 116388 127396 116390
rect 127100 115354 127156 115356
rect 127180 115354 127236 115356
rect 127260 115354 127316 115356
rect 127340 115354 127396 115356
rect 127100 115302 127126 115354
rect 127126 115302 127156 115354
rect 127180 115302 127190 115354
rect 127190 115302 127236 115354
rect 127260 115302 127306 115354
rect 127306 115302 127316 115354
rect 127340 115302 127370 115354
rect 127370 115302 127396 115354
rect 127100 115300 127156 115302
rect 127180 115300 127236 115302
rect 127260 115300 127316 115302
rect 127340 115300 127396 115302
rect 127100 114266 127156 114268
rect 127180 114266 127236 114268
rect 127260 114266 127316 114268
rect 127340 114266 127396 114268
rect 127100 114214 127126 114266
rect 127126 114214 127156 114266
rect 127180 114214 127190 114266
rect 127190 114214 127236 114266
rect 127260 114214 127306 114266
rect 127306 114214 127316 114266
rect 127340 114214 127370 114266
rect 127370 114214 127396 114266
rect 127100 114212 127156 114214
rect 127180 114212 127236 114214
rect 127260 114212 127316 114214
rect 127340 114212 127396 114214
rect 127100 113178 127156 113180
rect 127180 113178 127236 113180
rect 127260 113178 127316 113180
rect 127340 113178 127396 113180
rect 127100 113126 127126 113178
rect 127126 113126 127156 113178
rect 127180 113126 127190 113178
rect 127190 113126 127236 113178
rect 127260 113126 127306 113178
rect 127306 113126 127316 113178
rect 127340 113126 127370 113178
rect 127370 113126 127396 113178
rect 127100 113124 127156 113126
rect 127180 113124 127236 113126
rect 127260 113124 127316 113126
rect 127340 113124 127396 113126
rect 127100 112090 127156 112092
rect 127180 112090 127236 112092
rect 127260 112090 127316 112092
rect 127340 112090 127396 112092
rect 127100 112038 127126 112090
rect 127126 112038 127156 112090
rect 127180 112038 127190 112090
rect 127190 112038 127236 112090
rect 127260 112038 127306 112090
rect 127306 112038 127316 112090
rect 127340 112038 127370 112090
rect 127370 112038 127396 112090
rect 127100 112036 127156 112038
rect 127180 112036 127236 112038
rect 127260 112036 127316 112038
rect 127340 112036 127396 112038
rect 127100 111002 127156 111004
rect 127180 111002 127236 111004
rect 127260 111002 127316 111004
rect 127340 111002 127396 111004
rect 127100 110950 127126 111002
rect 127126 110950 127156 111002
rect 127180 110950 127190 111002
rect 127190 110950 127236 111002
rect 127260 110950 127306 111002
rect 127306 110950 127316 111002
rect 127340 110950 127370 111002
rect 127370 110950 127396 111002
rect 127100 110948 127156 110950
rect 127180 110948 127236 110950
rect 127260 110948 127316 110950
rect 127340 110948 127396 110950
rect 127100 109914 127156 109916
rect 127180 109914 127236 109916
rect 127260 109914 127316 109916
rect 127340 109914 127396 109916
rect 127100 109862 127126 109914
rect 127126 109862 127156 109914
rect 127180 109862 127190 109914
rect 127190 109862 127236 109914
rect 127260 109862 127306 109914
rect 127306 109862 127316 109914
rect 127340 109862 127370 109914
rect 127370 109862 127396 109914
rect 127100 109860 127156 109862
rect 127180 109860 127236 109862
rect 127260 109860 127316 109862
rect 127340 109860 127396 109862
rect 127100 108826 127156 108828
rect 127180 108826 127236 108828
rect 127260 108826 127316 108828
rect 127340 108826 127396 108828
rect 127100 108774 127126 108826
rect 127126 108774 127156 108826
rect 127180 108774 127190 108826
rect 127190 108774 127236 108826
rect 127260 108774 127306 108826
rect 127306 108774 127316 108826
rect 127340 108774 127370 108826
rect 127370 108774 127396 108826
rect 127100 108772 127156 108774
rect 127180 108772 127236 108774
rect 127260 108772 127316 108774
rect 127340 108772 127396 108774
rect 127100 107738 127156 107740
rect 127180 107738 127236 107740
rect 127260 107738 127316 107740
rect 127340 107738 127396 107740
rect 127100 107686 127126 107738
rect 127126 107686 127156 107738
rect 127180 107686 127190 107738
rect 127190 107686 127236 107738
rect 127260 107686 127306 107738
rect 127306 107686 127316 107738
rect 127340 107686 127370 107738
rect 127370 107686 127396 107738
rect 127100 107684 127156 107686
rect 127180 107684 127236 107686
rect 127260 107684 127316 107686
rect 127340 107684 127396 107686
rect 127100 106650 127156 106652
rect 127180 106650 127236 106652
rect 127260 106650 127316 106652
rect 127340 106650 127396 106652
rect 127100 106598 127126 106650
rect 127126 106598 127156 106650
rect 127180 106598 127190 106650
rect 127190 106598 127236 106650
rect 127260 106598 127306 106650
rect 127306 106598 127316 106650
rect 127340 106598 127370 106650
rect 127370 106598 127396 106650
rect 127100 106596 127156 106598
rect 127180 106596 127236 106598
rect 127260 106596 127316 106598
rect 127340 106596 127396 106598
rect 127100 105562 127156 105564
rect 127180 105562 127236 105564
rect 127260 105562 127316 105564
rect 127340 105562 127396 105564
rect 127100 105510 127126 105562
rect 127126 105510 127156 105562
rect 127180 105510 127190 105562
rect 127190 105510 127236 105562
rect 127260 105510 127306 105562
rect 127306 105510 127316 105562
rect 127340 105510 127370 105562
rect 127370 105510 127396 105562
rect 127100 105508 127156 105510
rect 127180 105508 127236 105510
rect 127260 105508 127316 105510
rect 127340 105508 127396 105510
rect 127100 104474 127156 104476
rect 127180 104474 127236 104476
rect 127260 104474 127316 104476
rect 127340 104474 127396 104476
rect 127100 104422 127126 104474
rect 127126 104422 127156 104474
rect 127180 104422 127190 104474
rect 127190 104422 127236 104474
rect 127260 104422 127306 104474
rect 127306 104422 127316 104474
rect 127340 104422 127370 104474
rect 127370 104422 127396 104474
rect 127100 104420 127156 104422
rect 127180 104420 127236 104422
rect 127260 104420 127316 104422
rect 127340 104420 127396 104422
rect 127100 103386 127156 103388
rect 127180 103386 127236 103388
rect 127260 103386 127316 103388
rect 127340 103386 127396 103388
rect 127100 103334 127126 103386
rect 127126 103334 127156 103386
rect 127180 103334 127190 103386
rect 127190 103334 127236 103386
rect 127260 103334 127306 103386
rect 127306 103334 127316 103386
rect 127340 103334 127370 103386
rect 127370 103334 127396 103386
rect 127100 103332 127156 103334
rect 127180 103332 127236 103334
rect 127260 103332 127316 103334
rect 127340 103332 127396 103334
rect 127100 102298 127156 102300
rect 127180 102298 127236 102300
rect 127260 102298 127316 102300
rect 127340 102298 127396 102300
rect 127100 102246 127126 102298
rect 127126 102246 127156 102298
rect 127180 102246 127190 102298
rect 127190 102246 127236 102298
rect 127260 102246 127306 102298
rect 127306 102246 127316 102298
rect 127340 102246 127370 102298
rect 127370 102246 127396 102298
rect 127100 102244 127156 102246
rect 127180 102244 127236 102246
rect 127260 102244 127316 102246
rect 127340 102244 127396 102246
rect 127100 101210 127156 101212
rect 127180 101210 127236 101212
rect 127260 101210 127316 101212
rect 127340 101210 127396 101212
rect 127100 101158 127126 101210
rect 127126 101158 127156 101210
rect 127180 101158 127190 101210
rect 127190 101158 127236 101210
rect 127260 101158 127306 101210
rect 127306 101158 127316 101210
rect 127340 101158 127370 101210
rect 127370 101158 127396 101210
rect 127100 101156 127156 101158
rect 127180 101156 127236 101158
rect 127260 101156 127316 101158
rect 127340 101156 127396 101158
rect 127100 100122 127156 100124
rect 127180 100122 127236 100124
rect 127260 100122 127316 100124
rect 127340 100122 127396 100124
rect 127100 100070 127126 100122
rect 127126 100070 127156 100122
rect 127180 100070 127190 100122
rect 127190 100070 127236 100122
rect 127260 100070 127306 100122
rect 127306 100070 127316 100122
rect 127340 100070 127370 100122
rect 127370 100070 127396 100122
rect 127100 100068 127156 100070
rect 127180 100068 127236 100070
rect 127260 100068 127316 100070
rect 127340 100068 127396 100070
rect 127100 99034 127156 99036
rect 127180 99034 127236 99036
rect 127260 99034 127316 99036
rect 127340 99034 127396 99036
rect 127100 98982 127126 99034
rect 127126 98982 127156 99034
rect 127180 98982 127190 99034
rect 127190 98982 127236 99034
rect 127260 98982 127306 99034
rect 127306 98982 127316 99034
rect 127340 98982 127370 99034
rect 127370 98982 127396 99034
rect 127100 98980 127156 98982
rect 127180 98980 127236 98982
rect 127260 98980 127316 98982
rect 127340 98980 127396 98982
rect 127100 97946 127156 97948
rect 127180 97946 127236 97948
rect 127260 97946 127316 97948
rect 127340 97946 127396 97948
rect 127100 97894 127126 97946
rect 127126 97894 127156 97946
rect 127180 97894 127190 97946
rect 127190 97894 127236 97946
rect 127260 97894 127306 97946
rect 127306 97894 127316 97946
rect 127340 97894 127370 97946
rect 127370 97894 127396 97946
rect 127100 97892 127156 97894
rect 127180 97892 127236 97894
rect 127260 97892 127316 97894
rect 127340 97892 127396 97894
rect 127100 96858 127156 96860
rect 127180 96858 127236 96860
rect 127260 96858 127316 96860
rect 127340 96858 127396 96860
rect 127100 96806 127126 96858
rect 127126 96806 127156 96858
rect 127180 96806 127190 96858
rect 127190 96806 127236 96858
rect 127260 96806 127306 96858
rect 127306 96806 127316 96858
rect 127340 96806 127370 96858
rect 127370 96806 127396 96858
rect 127100 96804 127156 96806
rect 127180 96804 127236 96806
rect 127260 96804 127316 96806
rect 127340 96804 127396 96806
rect 127100 95770 127156 95772
rect 127180 95770 127236 95772
rect 127260 95770 127316 95772
rect 127340 95770 127396 95772
rect 127100 95718 127126 95770
rect 127126 95718 127156 95770
rect 127180 95718 127190 95770
rect 127190 95718 127236 95770
rect 127260 95718 127306 95770
rect 127306 95718 127316 95770
rect 127340 95718 127370 95770
rect 127370 95718 127396 95770
rect 127100 95716 127156 95718
rect 127180 95716 127236 95718
rect 127260 95716 127316 95718
rect 127340 95716 127396 95718
rect 127100 94682 127156 94684
rect 127180 94682 127236 94684
rect 127260 94682 127316 94684
rect 127340 94682 127396 94684
rect 127100 94630 127126 94682
rect 127126 94630 127156 94682
rect 127180 94630 127190 94682
rect 127190 94630 127236 94682
rect 127260 94630 127306 94682
rect 127306 94630 127316 94682
rect 127340 94630 127370 94682
rect 127370 94630 127396 94682
rect 127100 94628 127156 94630
rect 127180 94628 127236 94630
rect 127260 94628 127316 94630
rect 127340 94628 127396 94630
rect 127100 93594 127156 93596
rect 127180 93594 127236 93596
rect 127260 93594 127316 93596
rect 127340 93594 127396 93596
rect 127100 93542 127126 93594
rect 127126 93542 127156 93594
rect 127180 93542 127190 93594
rect 127190 93542 127236 93594
rect 127260 93542 127306 93594
rect 127306 93542 127316 93594
rect 127340 93542 127370 93594
rect 127370 93542 127396 93594
rect 127100 93540 127156 93542
rect 127180 93540 127236 93542
rect 127260 93540 127316 93542
rect 127340 93540 127396 93542
rect 127100 92506 127156 92508
rect 127180 92506 127236 92508
rect 127260 92506 127316 92508
rect 127340 92506 127396 92508
rect 127100 92454 127126 92506
rect 127126 92454 127156 92506
rect 127180 92454 127190 92506
rect 127190 92454 127236 92506
rect 127260 92454 127306 92506
rect 127306 92454 127316 92506
rect 127340 92454 127370 92506
rect 127370 92454 127396 92506
rect 127100 92452 127156 92454
rect 127180 92452 127236 92454
rect 127260 92452 127316 92454
rect 127340 92452 127396 92454
rect 127100 91418 127156 91420
rect 127180 91418 127236 91420
rect 127260 91418 127316 91420
rect 127340 91418 127396 91420
rect 127100 91366 127126 91418
rect 127126 91366 127156 91418
rect 127180 91366 127190 91418
rect 127190 91366 127236 91418
rect 127260 91366 127306 91418
rect 127306 91366 127316 91418
rect 127340 91366 127370 91418
rect 127370 91366 127396 91418
rect 127100 91364 127156 91366
rect 127180 91364 127236 91366
rect 127260 91364 127316 91366
rect 127340 91364 127396 91366
rect 127100 90330 127156 90332
rect 127180 90330 127236 90332
rect 127260 90330 127316 90332
rect 127340 90330 127396 90332
rect 127100 90278 127126 90330
rect 127126 90278 127156 90330
rect 127180 90278 127190 90330
rect 127190 90278 127236 90330
rect 127260 90278 127306 90330
rect 127306 90278 127316 90330
rect 127340 90278 127370 90330
rect 127370 90278 127396 90330
rect 127100 90276 127156 90278
rect 127180 90276 127236 90278
rect 127260 90276 127316 90278
rect 127340 90276 127396 90278
rect 127100 89242 127156 89244
rect 127180 89242 127236 89244
rect 127260 89242 127316 89244
rect 127340 89242 127396 89244
rect 127100 89190 127126 89242
rect 127126 89190 127156 89242
rect 127180 89190 127190 89242
rect 127190 89190 127236 89242
rect 127260 89190 127306 89242
rect 127306 89190 127316 89242
rect 127340 89190 127370 89242
rect 127370 89190 127396 89242
rect 127100 89188 127156 89190
rect 127180 89188 127236 89190
rect 127260 89188 127316 89190
rect 127340 89188 127396 89190
rect 127100 88154 127156 88156
rect 127180 88154 127236 88156
rect 127260 88154 127316 88156
rect 127340 88154 127396 88156
rect 127100 88102 127126 88154
rect 127126 88102 127156 88154
rect 127180 88102 127190 88154
rect 127190 88102 127236 88154
rect 127260 88102 127306 88154
rect 127306 88102 127316 88154
rect 127340 88102 127370 88154
rect 127370 88102 127396 88154
rect 127100 88100 127156 88102
rect 127180 88100 127236 88102
rect 127260 88100 127316 88102
rect 127340 88100 127396 88102
rect 127100 87066 127156 87068
rect 127180 87066 127236 87068
rect 127260 87066 127316 87068
rect 127340 87066 127396 87068
rect 127100 87014 127126 87066
rect 127126 87014 127156 87066
rect 127180 87014 127190 87066
rect 127190 87014 127236 87066
rect 127260 87014 127306 87066
rect 127306 87014 127316 87066
rect 127340 87014 127370 87066
rect 127370 87014 127396 87066
rect 127100 87012 127156 87014
rect 127180 87012 127236 87014
rect 127260 87012 127316 87014
rect 127340 87012 127396 87014
rect 127100 85978 127156 85980
rect 127180 85978 127236 85980
rect 127260 85978 127316 85980
rect 127340 85978 127396 85980
rect 127100 85926 127126 85978
rect 127126 85926 127156 85978
rect 127180 85926 127190 85978
rect 127190 85926 127236 85978
rect 127260 85926 127306 85978
rect 127306 85926 127316 85978
rect 127340 85926 127370 85978
rect 127370 85926 127396 85978
rect 127100 85924 127156 85926
rect 127180 85924 127236 85926
rect 127260 85924 127316 85926
rect 127340 85924 127396 85926
rect 127100 84890 127156 84892
rect 127180 84890 127236 84892
rect 127260 84890 127316 84892
rect 127340 84890 127396 84892
rect 127100 84838 127126 84890
rect 127126 84838 127156 84890
rect 127180 84838 127190 84890
rect 127190 84838 127236 84890
rect 127260 84838 127306 84890
rect 127306 84838 127316 84890
rect 127340 84838 127370 84890
rect 127370 84838 127396 84890
rect 127100 84836 127156 84838
rect 127180 84836 127236 84838
rect 127260 84836 127316 84838
rect 127340 84836 127396 84838
rect 127100 83802 127156 83804
rect 127180 83802 127236 83804
rect 127260 83802 127316 83804
rect 127340 83802 127396 83804
rect 127100 83750 127126 83802
rect 127126 83750 127156 83802
rect 127180 83750 127190 83802
rect 127190 83750 127236 83802
rect 127260 83750 127306 83802
rect 127306 83750 127316 83802
rect 127340 83750 127370 83802
rect 127370 83750 127396 83802
rect 127100 83748 127156 83750
rect 127180 83748 127236 83750
rect 127260 83748 127316 83750
rect 127340 83748 127396 83750
rect 127100 82714 127156 82716
rect 127180 82714 127236 82716
rect 127260 82714 127316 82716
rect 127340 82714 127396 82716
rect 127100 82662 127126 82714
rect 127126 82662 127156 82714
rect 127180 82662 127190 82714
rect 127190 82662 127236 82714
rect 127260 82662 127306 82714
rect 127306 82662 127316 82714
rect 127340 82662 127370 82714
rect 127370 82662 127396 82714
rect 127100 82660 127156 82662
rect 127180 82660 127236 82662
rect 127260 82660 127316 82662
rect 127340 82660 127396 82662
rect 127100 81626 127156 81628
rect 127180 81626 127236 81628
rect 127260 81626 127316 81628
rect 127340 81626 127396 81628
rect 127100 81574 127126 81626
rect 127126 81574 127156 81626
rect 127180 81574 127190 81626
rect 127190 81574 127236 81626
rect 127260 81574 127306 81626
rect 127306 81574 127316 81626
rect 127340 81574 127370 81626
rect 127370 81574 127396 81626
rect 127100 81572 127156 81574
rect 127180 81572 127236 81574
rect 127260 81572 127316 81574
rect 127340 81572 127396 81574
rect 127100 80538 127156 80540
rect 127180 80538 127236 80540
rect 127260 80538 127316 80540
rect 127340 80538 127396 80540
rect 127100 80486 127126 80538
rect 127126 80486 127156 80538
rect 127180 80486 127190 80538
rect 127190 80486 127236 80538
rect 127260 80486 127306 80538
rect 127306 80486 127316 80538
rect 127340 80486 127370 80538
rect 127370 80486 127396 80538
rect 127100 80484 127156 80486
rect 127180 80484 127236 80486
rect 127260 80484 127316 80486
rect 127340 80484 127396 80486
rect 127100 79450 127156 79452
rect 127180 79450 127236 79452
rect 127260 79450 127316 79452
rect 127340 79450 127396 79452
rect 127100 79398 127126 79450
rect 127126 79398 127156 79450
rect 127180 79398 127190 79450
rect 127190 79398 127236 79450
rect 127260 79398 127306 79450
rect 127306 79398 127316 79450
rect 127340 79398 127370 79450
rect 127370 79398 127396 79450
rect 127100 79396 127156 79398
rect 127180 79396 127236 79398
rect 127260 79396 127316 79398
rect 127340 79396 127396 79398
rect 127100 78362 127156 78364
rect 127180 78362 127236 78364
rect 127260 78362 127316 78364
rect 127340 78362 127396 78364
rect 127100 78310 127126 78362
rect 127126 78310 127156 78362
rect 127180 78310 127190 78362
rect 127190 78310 127236 78362
rect 127260 78310 127306 78362
rect 127306 78310 127316 78362
rect 127340 78310 127370 78362
rect 127370 78310 127396 78362
rect 127100 78308 127156 78310
rect 127180 78308 127236 78310
rect 127260 78308 127316 78310
rect 127340 78308 127396 78310
rect 127100 77274 127156 77276
rect 127180 77274 127236 77276
rect 127260 77274 127316 77276
rect 127340 77274 127396 77276
rect 127100 77222 127126 77274
rect 127126 77222 127156 77274
rect 127180 77222 127190 77274
rect 127190 77222 127236 77274
rect 127260 77222 127306 77274
rect 127306 77222 127316 77274
rect 127340 77222 127370 77274
rect 127370 77222 127396 77274
rect 127100 77220 127156 77222
rect 127180 77220 127236 77222
rect 127260 77220 127316 77222
rect 127340 77220 127396 77222
rect 127100 76186 127156 76188
rect 127180 76186 127236 76188
rect 127260 76186 127316 76188
rect 127340 76186 127396 76188
rect 127100 76134 127126 76186
rect 127126 76134 127156 76186
rect 127180 76134 127190 76186
rect 127190 76134 127236 76186
rect 127260 76134 127306 76186
rect 127306 76134 127316 76186
rect 127340 76134 127370 76186
rect 127370 76134 127396 76186
rect 127100 76132 127156 76134
rect 127180 76132 127236 76134
rect 127260 76132 127316 76134
rect 127340 76132 127396 76134
rect 127100 75098 127156 75100
rect 127180 75098 127236 75100
rect 127260 75098 127316 75100
rect 127340 75098 127396 75100
rect 127100 75046 127126 75098
rect 127126 75046 127156 75098
rect 127180 75046 127190 75098
rect 127190 75046 127236 75098
rect 127260 75046 127306 75098
rect 127306 75046 127316 75098
rect 127340 75046 127370 75098
rect 127370 75046 127396 75098
rect 127100 75044 127156 75046
rect 127180 75044 127236 75046
rect 127260 75044 127316 75046
rect 127340 75044 127396 75046
rect 127100 74010 127156 74012
rect 127180 74010 127236 74012
rect 127260 74010 127316 74012
rect 127340 74010 127396 74012
rect 127100 73958 127126 74010
rect 127126 73958 127156 74010
rect 127180 73958 127190 74010
rect 127190 73958 127236 74010
rect 127260 73958 127306 74010
rect 127306 73958 127316 74010
rect 127340 73958 127370 74010
rect 127370 73958 127396 74010
rect 127100 73956 127156 73958
rect 127180 73956 127236 73958
rect 127260 73956 127316 73958
rect 127340 73956 127396 73958
rect 127100 72922 127156 72924
rect 127180 72922 127236 72924
rect 127260 72922 127316 72924
rect 127340 72922 127396 72924
rect 127100 72870 127126 72922
rect 127126 72870 127156 72922
rect 127180 72870 127190 72922
rect 127190 72870 127236 72922
rect 127260 72870 127306 72922
rect 127306 72870 127316 72922
rect 127340 72870 127370 72922
rect 127370 72870 127396 72922
rect 127100 72868 127156 72870
rect 127180 72868 127236 72870
rect 127260 72868 127316 72870
rect 127340 72868 127396 72870
rect 127100 71834 127156 71836
rect 127180 71834 127236 71836
rect 127260 71834 127316 71836
rect 127340 71834 127396 71836
rect 127100 71782 127126 71834
rect 127126 71782 127156 71834
rect 127180 71782 127190 71834
rect 127190 71782 127236 71834
rect 127260 71782 127306 71834
rect 127306 71782 127316 71834
rect 127340 71782 127370 71834
rect 127370 71782 127396 71834
rect 127100 71780 127156 71782
rect 127180 71780 127236 71782
rect 127260 71780 127316 71782
rect 127340 71780 127396 71782
rect 127100 70746 127156 70748
rect 127180 70746 127236 70748
rect 127260 70746 127316 70748
rect 127340 70746 127396 70748
rect 127100 70694 127126 70746
rect 127126 70694 127156 70746
rect 127180 70694 127190 70746
rect 127190 70694 127236 70746
rect 127260 70694 127306 70746
rect 127306 70694 127316 70746
rect 127340 70694 127370 70746
rect 127370 70694 127396 70746
rect 127100 70692 127156 70694
rect 127180 70692 127236 70694
rect 127260 70692 127316 70694
rect 127340 70692 127396 70694
rect 127100 69658 127156 69660
rect 127180 69658 127236 69660
rect 127260 69658 127316 69660
rect 127340 69658 127396 69660
rect 127100 69606 127126 69658
rect 127126 69606 127156 69658
rect 127180 69606 127190 69658
rect 127190 69606 127236 69658
rect 127260 69606 127306 69658
rect 127306 69606 127316 69658
rect 127340 69606 127370 69658
rect 127370 69606 127396 69658
rect 127100 69604 127156 69606
rect 127180 69604 127236 69606
rect 127260 69604 127316 69606
rect 127340 69604 127396 69606
rect 127100 68570 127156 68572
rect 127180 68570 127236 68572
rect 127260 68570 127316 68572
rect 127340 68570 127396 68572
rect 127100 68518 127126 68570
rect 127126 68518 127156 68570
rect 127180 68518 127190 68570
rect 127190 68518 127236 68570
rect 127260 68518 127306 68570
rect 127306 68518 127316 68570
rect 127340 68518 127370 68570
rect 127370 68518 127396 68570
rect 127100 68516 127156 68518
rect 127180 68516 127236 68518
rect 127260 68516 127316 68518
rect 127340 68516 127396 68518
rect 127100 67482 127156 67484
rect 127180 67482 127236 67484
rect 127260 67482 127316 67484
rect 127340 67482 127396 67484
rect 127100 67430 127126 67482
rect 127126 67430 127156 67482
rect 127180 67430 127190 67482
rect 127190 67430 127236 67482
rect 127260 67430 127306 67482
rect 127306 67430 127316 67482
rect 127340 67430 127370 67482
rect 127370 67430 127396 67482
rect 127100 67428 127156 67430
rect 127180 67428 127236 67430
rect 127260 67428 127316 67430
rect 127340 67428 127396 67430
rect 127100 66394 127156 66396
rect 127180 66394 127236 66396
rect 127260 66394 127316 66396
rect 127340 66394 127396 66396
rect 127100 66342 127126 66394
rect 127126 66342 127156 66394
rect 127180 66342 127190 66394
rect 127190 66342 127236 66394
rect 127260 66342 127306 66394
rect 127306 66342 127316 66394
rect 127340 66342 127370 66394
rect 127370 66342 127396 66394
rect 127100 66340 127156 66342
rect 127180 66340 127236 66342
rect 127260 66340 127316 66342
rect 127340 66340 127396 66342
rect 127100 65306 127156 65308
rect 127180 65306 127236 65308
rect 127260 65306 127316 65308
rect 127340 65306 127396 65308
rect 127100 65254 127126 65306
rect 127126 65254 127156 65306
rect 127180 65254 127190 65306
rect 127190 65254 127236 65306
rect 127260 65254 127306 65306
rect 127306 65254 127316 65306
rect 127340 65254 127370 65306
rect 127370 65254 127396 65306
rect 127100 65252 127156 65254
rect 127180 65252 127236 65254
rect 127260 65252 127316 65254
rect 127340 65252 127396 65254
rect 127100 64218 127156 64220
rect 127180 64218 127236 64220
rect 127260 64218 127316 64220
rect 127340 64218 127396 64220
rect 127100 64166 127126 64218
rect 127126 64166 127156 64218
rect 127180 64166 127190 64218
rect 127190 64166 127236 64218
rect 127260 64166 127306 64218
rect 127306 64166 127316 64218
rect 127340 64166 127370 64218
rect 127370 64166 127396 64218
rect 127100 64164 127156 64166
rect 127180 64164 127236 64166
rect 127260 64164 127316 64166
rect 127340 64164 127396 64166
rect 127100 63130 127156 63132
rect 127180 63130 127236 63132
rect 127260 63130 127316 63132
rect 127340 63130 127396 63132
rect 127100 63078 127126 63130
rect 127126 63078 127156 63130
rect 127180 63078 127190 63130
rect 127190 63078 127236 63130
rect 127260 63078 127306 63130
rect 127306 63078 127316 63130
rect 127340 63078 127370 63130
rect 127370 63078 127396 63130
rect 127100 63076 127156 63078
rect 127180 63076 127236 63078
rect 127260 63076 127316 63078
rect 127340 63076 127396 63078
rect 127100 62042 127156 62044
rect 127180 62042 127236 62044
rect 127260 62042 127316 62044
rect 127340 62042 127396 62044
rect 127100 61990 127126 62042
rect 127126 61990 127156 62042
rect 127180 61990 127190 62042
rect 127190 61990 127236 62042
rect 127260 61990 127306 62042
rect 127306 61990 127316 62042
rect 127340 61990 127370 62042
rect 127370 61990 127396 62042
rect 127100 61988 127156 61990
rect 127180 61988 127236 61990
rect 127260 61988 127316 61990
rect 127340 61988 127396 61990
rect 127100 60954 127156 60956
rect 127180 60954 127236 60956
rect 127260 60954 127316 60956
rect 127340 60954 127396 60956
rect 127100 60902 127126 60954
rect 127126 60902 127156 60954
rect 127180 60902 127190 60954
rect 127190 60902 127236 60954
rect 127260 60902 127306 60954
rect 127306 60902 127316 60954
rect 127340 60902 127370 60954
rect 127370 60902 127396 60954
rect 127100 60900 127156 60902
rect 127180 60900 127236 60902
rect 127260 60900 127316 60902
rect 127340 60900 127396 60902
rect 127100 59866 127156 59868
rect 127180 59866 127236 59868
rect 127260 59866 127316 59868
rect 127340 59866 127396 59868
rect 127100 59814 127126 59866
rect 127126 59814 127156 59866
rect 127180 59814 127190 59866
rect 127190 59814 127236 59866
rect 127260 59814 127306 59866
rect 127306 59814 127316 59866
rect 127340 59814 127370 59866
rect 127370 59814 127396 59866
rect 127100 59812 127156 59814
rect 127180 59812 127236 59814
rect 127260 59812 127316 59814
rect 127340 59812 127396 59814
rect 127100 58778 127156 58780
rect 127180 58778 127236 58780
rect 127260 58778 127316 58780
rect 127340 58778 127396 58780
rect 127100 58726 127126 58778
rect 127126 58726 127156 58778
rect 127180 58726 127190 58778
rect 127190 58726 127236 58778
rect 127260 58726 127306 58778
rect 127306 58726 127316 58778
rect 127340 58726 127370 58778
rect 127370 58726 127396 58778
rect 127100 58724 127156 58726
rect 127180 58724 127236 58726
rect 127260 58724 127316 58726
rect 127340 58724 127396 58726
rect 127100 57690 127156 57692
rect 127180 57690 127236 57692
rect 127260 57690 127316 57692
rect 127340 57690 127396 57692
rect 127100 57638 127126 57690
rect 127126 57638 127156 57690
rect 127180 57638 127190 57690
rect 127190 57638 127236 57690
rect 127260 57638 127306 57690
rect 127306 57638 127316 57690
rect 127340 57638 127370 57690
rect 127370 57638 127396 57690
rect 127100 57636 127156 57638
rect 127180 57636 127236 57638
rect 127260 57636 127316 57638
rect 127340 57636 127396 57638
rect 127100 56602 127156 56604
rect 127180 56602 127236 56604
rect 127260 56602 127316 56604
rect 127340 56602 127396 56604
rect 127100 56550 127126 56602
rect 127126 56550 127156 56602
rect 127180 56550 127190 56602
rect 127190 56550 127236 56602
rect 127260 56550 127306 56602
rect 127306 56550 127316 56602
rect 127340 56550 127370 56602
rect 127370 56550 127396 56602
rect 127100 56548 127156 56550
rect 127180 56548 127236 56550
rect 127260 56548 127316 56550
rect 127340 56548 127396 56550
rect 127100 55514 127156 55516
rect 127180 55514 127236 55516
rect 127260 55514 127316 55516
rect 127340 55514 127396 55516
rect 127100 55462 127126 55514
rect 127126 55462 127156 55514
rect 127180 55462 127190 55514
rect 127190 55462 127236 55514
rect 127260 55462 127306 55514
rect 127306 55462 127316 55514
rect 127340 55462 127370 55514
rect 127370 55462 127396 55514
rect 127100 55460 127156 55462
rect 127180 55460 127236 55462
rect 127260 55460 127316 55462
rect 127340 55460 127396 55462
rect 127100 54426 127156 54428
rect 127180 54426 127236 54428
rect 127260 54426 127316 54428
rect 127340 54426 127396 54428
rect 127100 54374 127126 54426
rect 127126 54374 127156 54426
rect 127180 54374 127190 54426
rect 127190 54374 127236 54426
rect 127260 54374 127306 54426
rect 127306 54374 127316 54426
rect 127340 54374 127370 54426
rect 127370 54374 127396 54426
rect 127100 54372 127156 54374
rect 127180 54372 127236 54374
rect 127260 54372 127316 54374
rect 127340 54372 127396 54374
rect 127100 53338 127156 53340
rect 127180 53338 127236 53340
rect 127260 53338 127316 53340
rect 127340 53338 127396 53340
rect 127100 53286 127126 53338
rect 127126 53286 127156 53338
rect 127180 53286 127190 53338
rect 127190 53286 127236 53338
rect 127260 53286 127306 53338
rect 127306 53286 127316 53338
rect 127340 53286 127370 53338
rect 127370 53286 127396 53338
rect 127100 53284 127156 53286
rect 127180 53284 127236 53286
rect 127260 53284 127316 53286
rect 127340 53284 127396 53286
rect 127100 52250 127156 52252
rect 127180 52250 127236 52252
rect 127260 52250 127316 52252
rect 127340 52250 127396 52252
rect 127100 52198 127126 52250
rect 127126 52198 127156 52250
rect 127180 52198 127190 52250
rect 127190 52198 127236 52250
rect 127260 52198 127306 52250
rect 127306 52198 127316 52250
rect 127340 52198 127370 52250
rect 127370 52198 127396 52250
rect 127100 52196 127156 52198
rect 127180 52196 127236 52198
rect 127260 52196 127316 52198
rect 127340 52196 127396 52198
rect 127100 51162 127156 51164
rect 127180 51162 127236 51164
rect 127260 51162 127316 51164
rect 127340 51162 127396 51164
rect 127100 51110 127126 51162
rect 127126 51110 127156 51162
rect 127180 51110 127190 51162
rect 127190 51110 127236 51162
rect 127260 51110 127306 51162
rect 127306 51110 127316 51162
rect 127340 51110 127370 51162
rect 127370 51110 127396 51162
rect 127100 51108 127156 51110
rect 127180 51108 127236 51110
rect 127260 51108 127316 51110
rect 127340 51108 127396 51110
rect 127100 50074 127156 50076
rect 127180 50074 127236 50076
rect 127260 50074 127316 50076
rect 127340 50074 127396 50076
rect 127100 50022 127126 50074
rect 127126 50022 127156 50074
rect 127180 50022 127190 50074
rect 127190 50022 127236 50074
rect 127260 50022 127306 50074
rect 127306 50022 127316 50074
rect 127340 50022 127370 50074
rect 127370 50022 127396 50074
rect 127100 50020 127156 50022
rect 127180 50020 127236 50022
rect 127260 50020 127316 50022
rect 127340 50020 127396 50022
rect 127100 48986 127156 48988
rect 127180 48986 127236 48988
rect 127260 48986 127316 48988
rect 127340 48986 127396 48988
rect 127100 48934 127126 48986
rect 127126 48934 127156 48986
rect 127180 48934 127190 48986
rect 127190 48934 127236 48986
rect 127260 48934 127306 48986
rect 127306 48934 127316 48986
rect 127340 48934 127370 48986
rect 127370 48934 127396 48986
rect 127100 48932 127156 48934
rect 127180 48932 127236 48934
rect 127260 48932 127316 48934
rect 127340 48932 127396 48934
rect 127100 47898 127156 47900
rect 127180 47898 127236 47900
rect 127260 47898 127316 47900
rect 127340 47898 127396 47900
rect 127100 47846 127126 47898
rect 127126 47846 127156 47898
rect 127180 47846 127190 47898
rect 127190 47846 127236 47898
rect 127260 47846 127306 47898
rect 127306 47846 127316 47898
rect 127340 47846 127370 47898
rect 127370 47846 127396 47898
rect 127100 47844 127156 47846
rect 127180 47844 127236 47846
rect 127260 47844 127316 47846
rect 127340 47844 127396 47846
rect 127100 46810 127156 46812
rect 127180 46810 127236 46812
rect 127260 46810 127316 46812
rect 127340 46810 127396 46812
rect 127100 46758 127126 46810
rect 127126 46758 127156 46810
rect 127180 46758 127190 46810
rect 127190 46758 127236 46810
rect 127260 46758 127306 46810
rect 127306 46758 127316 46810
rect 127340 46758 127370 46810
rect 127370 46758 127396 46810
rect 127100 46756 127156 46758
rect 127180 46756 127236 46758
rect 127260 46756 127316 46758
rect 127340 46756 127396 46758
rect 127100 45722 127156 45724
rect 127180 45722 127236 45724
rect 127260 45722 127316 45724
rect 127340 45722 127396 45724
rect 127100 45670 127126 45722
rect 127126 45670 127156 45722
rect 127180 45670 127190 45722
rect 127190 45670 127236 45722
rect 127260 45670 127306 45722
rect 127306 45670 127316 45722
rect 127340 45670 127370 45722
rect 127370 45670 127396 45722
rect 127100 45668 127156 45670
rect 127180 45668 127236 45670
rect 127260 45668 127316 45670
rect 127340 45668 127396 45670
rect 127100 44634 127156 44636
rect 127180 44634 127236 44636
rect 127260 44634 127316 44636
rect 127340 44634 127396 44636
rect 127100 44582 127126 44634
rect 127126 44582 127156 44634
rect 127180 44582 127190 44634
rect 127190 44582 127236 44634
rect 127260 44582 127306 44634
rect 127306 44582 127316 44634
rect 127340 44582 127370 44634
rect 127370 44582 127396 44634
rect 127100 44580 127156 44582
rect 127180 44580 127236 44582
rect 127260 44580 127316 44582
rect 127340 44580 127396 44582
rect 127100 43546 127156 43548
rect 127180 43546 127236 43548
rect 127260 43546 127316 43548
rect 127340 43546 127396 43548
rect 127100 43494 127126 43546
rect 127126 43494 127156 43546
rect 127180 43494 127190 43546
rect 127190 43494 127236 43546
rect 127260 43494 127306 43546
rect 127306 43494 127316 43546
rect 127340 43494 127370 43546
rect 127370 43494 127396 43546
rect 127100 43492 127156 43494
rect 127180 43492 127236 43494
rect 127260 43492 127316 43494
rect 127340 43492 127396 43494
rect 127100 42458 127156 42460
rect 127180 42458 127236 42460
rect 127260 42458 127316 42460
rect 127340 42458 127396 42460
rect 127100 42406 127126 42458
rect 127126 42406 127156 42458
rect 127180 42406 127190 42458
rect 127190 42406 127236 42458
rect 127260 42406 127306 42458
rect 127306 42406 127316 42458
rect 127340 42406 127370 42458
rect 127370 42406 127396 42458
rect 127100 42404 127156 42406
rect 127180 42404 127236 42406
rect 127260 42404 127316 42406
rect 127340 42404 127396 42406
rect 127100 41370 127156 41372
rect 127180 41370 127236 41372
rect 127260 41370 127316 41372
rect 127340 41370 127396 41372
rect 127100 41318 127126 41370
rect 127126 41318 127156 41370
rect 127180 41318 127190 41370
rect 127190 41318 127236 41370
rect 127260 41318 127306 41370
rect 127306 41318 127316 41370
rect 127340 41318 127370 41370
rect 127370 41318 127396 41370
rect 127100 41316 127156 41318
rect 127180 41316 127236 41318
rect 127260 41316 127316 41318
rect 127340 41316 127396 41318
rect 127100 40282 127156 40284
rect 127180 40282 127236 40284
rect 127260 40282 127316 40284
rect 127340 40282 127396 40284
rect 127100 40230 127126 40282
rect 127126 40230 127156 40282
rect 127180 40230 127190 40282
rect 127190 40230 127236 40282
rect 127260 40230 127306 40282
rect 127306 40230 127316 40282
rect 127340 40230 127370 40282
rect 127370 40230 127396 40282
rect 127100 40228 127156 40230
rect 127180 40228 127236 40230
rect 127260 40228 127316 40230
rect 127340 40228 127396 40230
rect 127100 39194 127156 39196
rect 127180 39194 127236 39196
rect 127260 39194 127316 39196
rect 127340 39194 127396 39196
rect 127100 39142 127126 39194
rect 127126 39142 127156 39194
rect 127180 39142 127190 39194
rect 127190 39142 127236 39194
rect 127260 39142 127306 39194
rect 127306 39142 127316 39194
rect 127340 39142 127370 39194
rect 127370 39142 127396 39194
rect 127100 39140 127156 39142
rect 127180 39140 127236 39142
rect 127260 39140 127316 39142
rect 127340 39140 127396 39142
rect 127100 38106 127156 38108
rect 127180 38106 127236 38108
rect 127260 38106 127316 38108
rect 127340 38106 127396 38108
rect 127100 38054 127126 38106
rect 127126 38054 127156 38106
rect 127180 38054 127190 38106
rect 127190 38054 127236 38106
rect 127260 38054 127306 38106
rect 127306 38054 127316 38106
rect 127340 38054 127370 38106
rect 127370 38054 127396 38106
rect 127100 38052 127156 38054
rect 127180 38052 127236 38054
rect 127260 38052 127316 38054
rect 127340 38052 127396 38054
rect 127100 37018 127156 37020
rect 127180 37018 127236 37020
rect 127260 37018 127316 37020
rect 127340 37018 127396 37020
rect 127100 36966 127126 37018
rect 127126 36966 127156 37018
rect 127180 36966 127190 37018
rect 127190 36966 127236 37018
rect 127260 36966 127306 37018
rect 127306 36966 127316 37018
rect 127340 36966 127370 37018
rect 127370 36966 127396 37018
rect 127100 36964 127156 36966
rect 127180 36964 127236 36966
rect 127260 36964 127316 36966
rect 127340 36964 127396 36966
rect 127100 35930 127156 35932
rect 127180 35930 127236 35932
rect 127260 35930 127316 35932
rect 127340 35930 127396 35932
rect 127100 35878 127126 35930
rect 127126 35878 127156 35930
rect 127180 35878 127190 35930
rect 127190 35878 127236 35930
rect 127260 35878 127306 35930
rect 127306 35878 127316 35930
rect 127340 35878 127370 35930
rect 127370 35878 127396 35930
rect 127100 35876 127156 35878
rect 127180 35876 127236 35878
rect 127260 35876 127316 35878
rect 127340 35876 127396 35878
rect 127100 34842 127156 34844
rect 127180 34842 127236 34844
rect 127260 34842 127316 34844
rect 127340 34842 127396 34844
rect 127100 34790 127126 34842
rect 127126 34790 127156 34842
rect 127180 34790 127190 34842
rect 127190 34790 127236 34842
rect 127260 34790 127306 34842
rect 127306 34790 127316 34842
rect 127340 34790 127370 34842
rect 127370 34790 127396 34842
rect 127100 34788 127156 34790
rect 127180 34788 127236 34790
rect 127260 34788 127316 34790
rect 127340 34788 127396 34790
rect 127100 33754 127156 33756
rect 127180 33754 127236 33756
rect 127260 33754 127316 33756
rect 127340 33754 127396 33756
rect 127100 33702 127126 33754
rect 127126 33702 127156 33754
rect 127180 33702 127190 33754
rect 127190 33702 127236 33754
rect 127260 33702 127306 33754
rect 127306 33702 127316 33754
rect 127340 33702 127370 33754
rect 127370 33702 127396 33754
rect 127100 33700 127156 33702
rect 127180 33700 127236 33702
rect 127260 33700 127316 33702
rect 127340 33700 127396 33702
rect 127100 32666 127156 32668
rect 127180 32666 127236 32668
rect 127260 32666 127316 32668
rect 127340 32666 127396 32668
rect 127100 32614 127126 32666
rect 127126 32614 127156 32666
rect 127180 32614 127190 32666
rect 127190 32614 127236 32666
rect 127260 32614 127306 32666
rect 127306 32614 127316 32666
rect 127340 32614 127370 32666
rect 127370 32614 127396 32666
rect 127100 32612 127156 32614
rect 127180 32612 127236 32614
rect 127260 32612 127316 32614
rect 127340 32612 127396 32614
rect 127100 31578 127156 31580
rect 127180 31578 127236 31580
rect 127260 31578 127316 31580
rect 127340 31578 127396 31580
rect 127100 31526 127126 31578
rect 127126 31526 127156 31578
rect 127180 31526 127190 31578
rect 127190 31526 127236 31578
rect 127260 31526 127306 31578
rect 127306 31526 127316 31578
rect 127340 31526 127370 31578
rect 127370 31526 127396 31578
rect 127100 31524 127156 31526
rect 127180 31524 127236 31526
rect 127260 31524 127316 31526
rect 127340 31524 127396 31526
rect 127100 30490 127156 30492
rect 127180 30490 127236 30492
rect 127260 30490 127316 30492
rect 127340 30490 127396 30492
rect 127100 30438 127126 30490
rect 127126 30438 127156 30490
rect 127180 30438 127190 30490
rect 127190 30438 127236 30490
rect 127260 30438 127306 30490
rect 127306 30438 127316 30490
rect 127340 30438 127370 30490
rect 127370 30438 127396 30490
rect 127100 30436 127156 30438
rect 127180 30436 127236 30438
rect 127260 30436 127316 30438
rect 127340 30436 127396 30438
rect 127100 29402 127156 29404
rect 127180 29402 127236 29404
rect 127260 29402 127316 29404
rect 127340 29402 127396 29404
rect 127100 29350 127126 29402
rect 127126 29350 127156 29402
rect 127180 29350 127190 29402
rect 127190 29350 127236 29402
rect 127260 29350 127306 29402
rect 127306 29350 127316 29402
rect 127340 29350 127370 29402
rect 127370 29350 127396 29402
rect 127100 29348 127156 29350
rect 127180 29348 127236 29350
rect 127260 29348 127316 29350
rect 127340 29348 127396 29350
rect 127100 28314 127156 28316
rect 127180 28314 127236 28316
rect 127260 28314 127316 28316
rect 127340 28314 127396 28316
rect 127100 28262 127126 28314
rect 127126 28262 127156 28314
rect 127180 28262 127190 28314
rect 127190 28262 127236 28314
rect 127260 28262 127306 28314
rect 127306 28262 127316 28314
rect 127340 28262 127370 28314
rect 127370 28262 127396 28314
rect 127100 28260 127156 28262
rect 127180 28260 127236 28262
rect 127260 28260 127316 28262
rect 127340 28260 127396 28262
rect 127100 27226 127156 27228
rect 127180 27226 127236 27228
rect 127260 27226 127316 27228
rect 127340 27226 127396 27228
rect 127100 27174 127126 27226
rect 127126 27174 127156 27226
rect 127180 27174 127190 27226
rect 127190 27174 127236 27226
rect 127260 27174 127306 27226
rect 127306 27174 127316 27226
rect 127340 27174 127370 27226
rect 127370 27174 127396 27226
rect 127100 27172 127156 27174
rect 127180 27172 127236 27174
rect 127260 27172 127316 27174
rect 127340 27172 127396 27174
rect 127100 26138 127156 26140
rect 127180 26138 127236 26140
rect 127260 26138 127316 26140
rect 127340 26138 127396 26140
rect 127100 26086 127126 26138
rect 127126 26086 127156 26138
rect 127180 26086 127190 26138
rect 127190 26086 127236 26138
rect 127260 26086 127306 26138
rect 127306 26086 127316 26138
rect 127340 26086 127370 26138
rect 127370 26086 127396 26138
rect 127100 26084 127156 26086
rect 127180 26084 127236 26086
rect 127260 26084 127316 26086
rect 127340 26084 127396 26086
rect 127100 25050 127156 25052
rect 127180 25050 127236 25052
rect 127260 25050 127316 25052
rect 127340 25050 127396 25052
rect 127100 24998 127126 25050
rect 127126 24998 127156 25050
rect 127180 24998 127190 25050
rect 127190 24998 127236 25050
rect 127260 24998 127306 25050
rect 127306 24998 127316 25050
rect 127340 24998 127370 25050
rect 127370 24998 127396 25050
rect 127100 24996 127156 24998
rect 127180 24996 127236 24998
rect 127260 24996 127316 24998
rect 127340 24996 127396 24998
rect 127100 23962 127156 23964
rect 127180 23962 127236 23964
rect 127260 23962 127316 23964
rect 127340 23962 127396 23964
rect 127100 23910 127126 23962
rect 127126 23910 127156 23962
rect 127180 23910 127190 23962
rect 127190 23910 127236 23962
rect 127260 23910 127306 23962
rect 127306 23910 127316 23962
rect 127340 23910 127370 23962
rect 127370 23910 127396 23962
rect 127100 23908 127156 23910
rect 127180 23908 127236 23910
rect 127260 23908 127316 23910
rect 127340 23908 127396 23910
rect 127100 22874 127156 22876
rect 127180 22874 127236 22876
rect 127260 22874 127316 22876
rect 127340 22874 127396 22876
rect 127100 22822 127126 22874
rect 127126 22822 127156 22874
rect 127180 22822 127190 22874
rect 127190 22822 127236 22874
rect 127260 22822 127306 22874
rect 127306 22822 127316 22874
rect 127340 22822 127370 22874
rect 127370 22822 127396 22874
rect 127100 22820 127156 22822
rect 127180 22820 127236 22822
rect 127260 22820 127316 22822
rect 127340 22820 127396 22822
rect 127100 21786 127156 21788
rect 127180 21786 127236 21788
rect 127260 21786 127316 21788
rect 127340 21786 127396 21788
rect 127100 21734 127126 21786
rect 127126 21734 127156 21786
rect 127180 21734 127190 21786
rect 127190 21734 127236 21786
rect 127260 21734 127306 21786
rect 127306 21734 127316 21786
rect 127340 21734 127370 21786
rect 127370 21734 127396 21786
rect 127100 21732 127156 21734
rect 127180 21732 127236 21734
rect 127260 21732 127316 21734
rect 127340 21732 127396 21734
rect 127100 20698 127156 20700
rect 127180 20698 127236 20700
rect 127260 20698 127316 20700
rect 127340 20698 127396 20700
rect 127100 20646 127126 20698
rect 127126 20646 127156 20698
rect 127180 20646 127190 20698
rect 127190 20646 127236 20698
rect 127260 20646 127306 20698
rect 127306 20646 127316 20698
rect 127340 20646 127370 20698
rect 127370 20646 127396 20698
rect 127100 20644 127156 20646
rect 127180 20644 127236 20646
rect 127260 20644 127316 20646
rect 127340 20644 127396 20646
rect 96380 19610 96436 19612
rect 96460 19610 96516 19612
rect 96540 19610 96596 19612
rect 96620 19610 96676 19612
rect 96380 19558 96406 19610
rect 96406 19558 96436 19610
rect 96460 19558 96470 19610
rect 96470 19558 96516 19610
rect 96540 19558 96586 19610
rect 96586 19558 96596 19610
rect 96620 19558 96650 19610
rect 96650 19558 96676 19610
rect 96380 19556 96436 19558
rect 96460 19556 96516 19558
rect 96540 19556 96596 19558
rect 96620 19556 96676 19558
rect 127100 19610 127156 19612
rect 127180 19610 127236 19612
rect 127260 19610 127316 19612
rect 127340 19610 127396 19612
rect 127100 19558 127126 19610
rect 127126 19558 127156 19610
rect 127180 19558 127190 19610
rect 127190 19558 127236 19610
rect 127260 19558 127306 19610
rect 127306 19558 127316 19610
rect 127340 19558 127370 19610
rect 127370 19558 127396 19610
rect 127100 19556 127156 19558
rect 127180 19556 127236 19558
rect 127260 19556 127316 19558
rect 127340 19556 127396 19558
rect 142460 116986 142516 116988
rect 142540 116986 142596 116988
rect 142620 116986 142676 116988
rect 142700 116986 142756 116988
rect 142460 116934 142486 116986
rect 142486 116934 142516 116986
rect 142540 116934 142550 116986
rect 142550 116934 142596 116986
rect 142620 116934 142666 116986
rect 142666 116934 142676 116986
rect 142700 116934 142730 116986
rect 142730 116934 142756 116986
rect 142460 116932 142516 116934
rect 142540 116932 142596 116934
rect 142620 116932 142676 116934
rect 142700 116932 142756 116934
rect 142460 115898 142516 115900
rect 142540 115898 142596 115900
rect 142620 115898 142676 115900
rect 142700 115898 142756 115900
rect 142460 115846 142486 115898
rect 142486 115846 142516 115898
rect 142540 115846 142550 115898
rect 142550 115846 142596 115898
rect 142620 115846 142666 115898
rect 142666 115846 142676 115898
rect 142700 115846 142730 115898
rect 142730 115846 142756 115898
rect 142460 115844 142516 115846
rect 142540 115844 142596 115846
rect 142620 115844 142676 115846
rect 142700 115844 142756 115846
rect 142460 114810 142516 114812
rect 142540 114810 142596 114812
rect 142620 114810 142676 114812
rect 142700 114810 142756 114812
rect 142460 114758 142486 114810
rect 142486 114758 142516 114810
rect 142540 114758 142550 114810
rect 142550 114758 142596 114810
rect 142620 114758 142666 114810
rect 142666 114758 142676 114810
rect 142700 114758 142730 114810
rect 142730 114758 142756 114810
rect 142460 114756 142516 114758
rect 142540 114756 142596 114758
rect 142620 114756 142676 114758
rect 142700 114756 142756 114758
rect 142460 113722 142516 113724
rect 142540 113722 142596 113724
rect 142620 113722 142676 113724
rect 142700 113722 142756 113724
rect 142460 113670 142486 113722
rect 142486 113670 142516 113722
rect 142540 113670 142550 113722
rect 142550 113670 142596 113722
rect 142620 113670 142666 113722
rect 142666 113670 142676 113722
rect 142700 113670 142730 113722
rect 142730 113670 142756 113722
rect 142460 113668 142516 113670
rect 142540 113668 142596 113670
rect 142620 113668 142676 113670
rect 142700 113668 142756 113670
rect 142460 112634 142516 112636
rect 142540 112634 142596 112636
rect 142620 112634 142676 112636
rect 142700 112634 142756 112636
rect 142460 112582 142486 112634
rect 142486 112582 142516 112634
rect 142540 112582 142550 112634
rect 142550 112582 142596 112634
rect 142620 112582 142666 112634
rect 142666 112582 142676 112634
rect 142700 112582 142730 112634
rect 142730 112582 142756 112634
rect 142460 112580 142516 112582
rect 142540 112580 142596 112582
rect 142620 112580 142676 112582
rect 142700 112580 142756 112582
rect 142460 111546 142516 111548
rect 142540 111546 142596 111548
rect 142620 111546 142676 111548
rect 142700 111546 142756 111548
rect 142460 111494 142486 111546
rect 142486 111494 142516 111546
rect 142540 111494 142550 111546
rect 142550 111494 142596 111546
rect 142620 111494 142666 111546
rect 142666 111494 142676 111546
rect 142700 111494 142730 111546
rect 142730 111494 142756 111546
rect 142460 111492 142516 111494
rect 142540 111492 142596 111494
rect 142620 111492 142676 111494
rect 142700 111492 142756 111494
rect 142460 110458 142516 110460
rect 142540 110458 142596 110460
rect 142620 110458 142676 110460
rect 142700 110458 142756 110460
rect 142460 110406 142486 110458
rect 142486 110406 142516 110458
rect 142540 110406 142550 110458
rect 142550 110406 142596 110458
rect 142620 110406 142666 110458
rect 142666 110406 142676 110458
rect 142700 110406 142730 110458
rect 142730 110406 142756 110458
rect 142460 110404 142516 110406
rect 142540 110404 142596 110406
rect 142620 110404 142676 110406
rect 142700 110404 142756 110406
rect 142460 109370 142516 109372
rect 142540 109370 142596 109372
rect 142620 109370 142676 109372
rect 142700 109370 142756 109372
rect 142460 109318 142486 109370
rect 142486 109318 142516 109370
rect 142540 109318 142550 109370
rect 142550 109318 142596 109370
rect 142620 109318 142666 109370
rect 142666 109318 142676 109370
rect 142700 109318 142730 109370
rect 142730 109318 142756 109370
rect 142460 109316 142516 109318
rect 142540 109316 142596 109318
rect 142620 109316 142676 109318
rect 142700 109316 142756 109318
rect 142460 108282 142516 108284
rect 142540 108282 142596 108284
rect 142620 108282 142676 108284
rect 142700 108282 142756 108284
rect 142460 108230 142486 108282
rect 142486 108230 142516 108282
rect 142540 108230 142550 108282
rect 142550 108230 142596 108282
rect 142620 108230 142666 108282
rect 142666 108230 142676 108282
rect 142700 108230 142730 108282
rect 142730 108230 142756 108282
rect 142460 108228 142516 108230
rect 142540 108228 142596 108230
rect 142620 108228 142676 108230
rect 142700 108228 142756 108230
rect 142460 107194 142516 107196
rect 142540 107194 142596 107196
rect 142620 107194 142676 107196
rect 142700 107194 142756 107196
rect 142460 107142 142486 107194
rect 142486 107142 142516 107194
rect 142540 107142 142550 107194
rect 142550 107142 142596 107194
rect 142620 107142 142666 107194
rect 142666 107142 142676 107194
rect 142700 107142 142730 107194
rect 142730 107142 142756 107194
rect 142460 107140 142516 107142
rect 142540 107140 142596 107142
rect 142620 107140 142676 107142
rect 142700 107140 142756 107142
rect 142460 106106 142516 106108
rect 142540 106106 142596 106108
rect 142620 106106 142676 106108
rect 142700 106106 142756 106108
rect 142460 106054 142486 106106
rect 142486 106054 142516 106106
rect 142540 106054 142550 106106
rect 142550 106054 142596 106106
rect 142620 106054 142666 106106
rect 142666 106054 142676 106106
rect 142700 106054 142730 106106
rect 142730 106054 142756 106106
rect 142460 106052 142516 106054
rect 142540 106052 142596 106054
rect 142620 106052 142676 106054
rect 142700 106052 142756 106054
rect 142460 105018 142516 105020
rect 142540 105018 142596 105020
rect 142620 105018 142676 105020
rect 142700 105018 142756 105020
rect 142460 104966 142486 105018
rect 142486 104966 142516 105018
rect 142540 104966 142550 105018
rect 142550 104966 142596 105018
rect 142620 104966 142666 105018
rect 142666 104966 142676 105018
rect 142700 104966 142730 105018
rect 142730 104966 142756 105018
rect 142460 104964 142516 104966
rect 142540 104964 142596 104966
rect 142620 104964 142676 104966
rect 142700 104964 142756 104966
rect 142460 103930 142516 103932
rect 142540 103930 142596 103932
rect 142620 103930 142676 103932
rect 142700 103930 142756 103932
rect 142460 103878 142486 103930
rect 142486 103878 142516 103930
rect 142540 103878 142550 103930
rect 142550 103878 142596 103930
rect 142620 103878 142666 103930
rect 142666 103878 142676 103930
rect 142700 103878 142730 103930
rect 142730 103878 142756 103930
rect 142460 103876 142516 103878
rect 142540 103876 142596 103878
rect 142620 103876 142676 103878
rect 142700 103876 142756 103878
rect 142460 102842 142516 102844
rect 142540 102842 142596 102844
rect 142620 102842 142676 102844
rect 142700 102842 142756 102844
rect 142460 102790 142486 102842
rect 142486 102790 142516 102842
rect 142540 102790 142550 102842
rect 142550 102790 142596 102842
rect 142620 102790 142666 102842
rect 142666 102790 142676 102842
rect 142700 102790 142730 102842
rect 142730 102790 142756 102842
rect 142460 102788 142516 102790
rect 142540 102788 142596 102790
rect 142620 102788 142676 102790
rect 142700 102788 142756 102790
rect 142460 101754 142516 101756
rect 142540 101754 142596 101756
rect 142620 101754 142676 101756
rect 142700 101754 142756 101756
rect 142460 101702 142486 101754
rect 142486 101702 142516 101754
rect 142540 101702 142550 101754
rect 142550 101702 142596 101754
rect 142620 101702 142666 101754
rect 142666 101702 142676 101754
rect 142700 101702 142730 101754
rect 142730 101702 142756 101754
rect 142460 101700 142516 101702
rect 142540 101700 142596 101702
rect 142620 101700 142676 101702
rect 142700 101700 142756 101702
rect 142460 100666 142516 100668
rect 142540 100666 142596 100668
rect 142620 100666 142676 100668
rect 142700 100666 142756 100668
rect 142460 100614 142486 100666
rect 142486 100614 142516 100666
rect 142540 100614 142550 100666
rect 142550 100614 142596 100666
rect 142620 100614 142666 100666
rect 142666 100614 142676 100666
rect 142700 100614 142730 100666
rect 142730 100614 142756 100666
rect 142460 100612 142516 100614
rect 142540 100612 142596 100614
rect 142620 100612 142676 100614
rect 142700 100612 142756 100614
rect 142460 99578 142516 99580
rect 142540 99578 142596 99580
rect 142620 99578 142676 99580
rect 142700 99578 142756 99580
rect 142460 99526 142486 99578
rect 142486 99526 142516 99578
rect 142540 99526 142550 99578
rect 142550 99526 142596 99578
rect 142620 99526 142666 99578
rect 142666 99526 142676 99578
rect 142700 99526 142730 99578
rect 142730 99526 142756 99578
rect 142460 99524 142516 99526
rect 142540 99524 142596 99526
rect 142620 99524 142676 99526
rect 142700 99524 142756 99526
rect 142460 98490 142516 98492
rect 142540 98490 142596 98492
rect 142620 98490 142676 98492
rect 142700 98490 142756 98492
rect 142460 98438 142486 98490
rect 142486 98438 142516 98490
rect 142540 98438 142550 98490
rect 142550 98438 142596 98490
rect 142620 98438 142666 98490
rect 142666 98438 142676 98490
rect 142700 98438 142730 98490
rect 142730 98438 142756 98490
rect 142460 98436 142516 98438
rect 142540 98436 142596 98438
rect 142620 98436 142676 98438
rect 142700 98436 142756 98438
rect 142460 97402 142516 97404
rect 142540 97402 142596 97404
rect 142620 97402 142676 97404
rect 142700 97402 142756 97404
rect 142460 97350 142486 97402
rect 142486 97350 142516 97402
rect 142540 97350 142550 97402
rect 142550 97350 142596 97402
rect 142620 97350 142666 97402
rect 142666 97350 142676 97402
rect 142700 97350 142730 97402
rect 142730 97350 142756 97402
rect 142460 97348 142516 97350
rect 142540 97348 142596 97350
rect 142620 97348 142676 97350
rect 142700 97348 142756 97350
rect 142460 96314 142516 96316
rect 142540 96314 142596 96316
rect 142620 96314 142676 96316
rect 142700 96314 142756 96316
rect 142460 96262 142486 96314
rect 142486 96262 142516 96314
rect 142540 96262 142550 96314
rect 142550 96262 142596 96314
rect 142620 96262 142666 96314
rect 142666 96262 142676 96314
rect 142700 96262 142730 96314
rect 142730 96262 142756 96314
rect 142460 96260 142516 96262
rect 142540 96260 142596 96262
rect 142620 96260 142676 96262
rect 142700 96260 142756 96262
rect 142460 95226 142516 95228
rect 142540 95226 142596 95228
rect 142620 95226 142676 95228
rect 142700 95226 142756 95228
rect 142460 95174 142486 95226
rect 142486 95174 142516 95226
rect 142540 95174 142550 95226
rect 142550 95174 142596 95226
rect 142620 95174 142666 95226
rect 142666 95174 142676 95226
rect 142700 95174 142730 95226
rect 142730 95174 142756 95226
rect 142460 95172 142516 95174
rect 142540 95172 142596 95174
rect 142620 95172 142676 95174
rect 142700 95172 142756 95174
rect 142460 94138 142516 94140
rect 142540 94138 142596 94140
rect 142620 94138 142676 94140
rect 142700 94138 142756 94140
rect 142460 94086 142486 94138
rect 142486 94086 142516 94138
rect 142540 94086 142550 94138
rect 142550 94086 142596 94138
rect 142620 94086 142666 94138
rect 142666 94086 142676 94138
rect 142700 94086 142730 94138
rect 142730 94086 142756 94138
rect 142460 94084 142516 94086
rect 142540 94084 142596 94086
rect 142620 94084 142676 94086
rect 142700 94084 142756 94086
rect 142460 93050 142516 93052
rect 142540 93050 142596 93052
rect 142620 93050 142676 93052
rect 142700 93050 142756 93052
rect 142460 92998 142486 93050
rect 142486 92998 142516 93050
rect 142540 92998 142550 93050
rect 142550 92998 142596 93050
rect 142620 92998 142666 93050
rect 142666 92998 142676 93050
rect 142700 92998 142730 93050
rect 142730 92998 142756 93050
rect 142460 92996 142516 92998
rect 142540 92996 142596 92998
rect 142620 92996 142676 92998
rect 142700 92996 142756 92998
rect 142460 91962 142516 91964
rect 142540 91962 142596 91964
rect 142620 91962 142676 91964
rect 142700 91962 142756 91964
rect 142460 91910 142486 91962
rect 142486 91910 142516 91962
rect 142540 91910 142550 91962
rect 142550 91910 142596 91962
rect 142620 91910 142666 91962
rect 142666 91910 142676 91962
rect 142700 91910 142730 91962
rect 142730 91910 142756 91962
rect 142460 91908 142516 91910
rect 142540 91908 142596 91910
rect 142620 91908 142676 91910
rect 142700 91908 142756 91910
rect 142460 90874 142516 90876
rect 142540 90874 142596 90876
rect 142620 90874 142676 90876
rect 142700 90874 142756 90876
rect 142460 90822 142486 90874
rect 142486 90822 142516 90874
rect 142540 90822 142550 90874
rect 142550 90822 142596 90874
rect 142620 90822 142666 90874
rect 142666 90822 142676 90874
rect 142700 90822 142730 90874
rect 142730 90822 142756 90874
rect 142460 90820 142516 90822
rect 142540 90820 142596 90822
rect 142620 90820 142676 90822
rect 142700 90820 142756 90822
rect 142460 89786 142516 89788
rect 142540 89786 142596 89788
rect 142620 89786 142676 89788
rect 142700 89786 142756 89788
rect 142460 89734 142486 89786
rect 142486 89734 142516 89786
rect 142540 89734 142550 89786
rect 142550 89734 142596 89786
rect 142620 89734 142666 89786
rect 142666 89734 142676 89786
rect 142700 89734 142730 89786
rect 142730 89734 142756 89786
rect 142460 89732 142516 89734
rect 142540 89732 142596 89734
rect 142620 89732 142676 89734
rect 142700 89732 142756 89734
rect 142460 88698 142516 88700
rect 142540 88698 142596 88700
rect 142620 88698 142676 88700
rect 142700 88698 142756 88700
rect 142460 88646 142486 88698
rect 142486 88646 142516 88698
rect 142540 88646 142550 88698
rect 142550 88646 142596 88698
rect 142620 88646 142666 88698
rect 142666 88646 142676 88698
rect 142700 88646 142730 88698
rect 142730 88646 142756 88698
rect 142460 88644 142516 88646
rect 142540 88644 142596 88646
rect 142620 88644 142676 88646
rect 142700 88644 142756 88646
rect 142460 87610 142516 87612
rect 142540 87610 142596 87612
rect 142620 87610 142676 87612
rect 142700 87610 142756 87612
rect 142460 87558 142486 87610
rect 142486 87558 142516 87610
rect 142540 87558 142550 87610
rect 142550 87558 142596 87610
rect 142620 87558 142666 87610
rect 142666 87558 142676 87610
rect 142700 87558 142730 87610
rect 142730 87558 142756 87610
rect 142460 87556 142516 87558
rect 142540 87556 142596 87558
rect 142620 87556 142676 87558
rect 142700 87556 142756 87558
rect 142460 86522 142516 86524
rect 142540 86522 142596 86524
rect 142620 86522 142676 86524
rect 142700 86522 142756 86524
rect 142460 86470 142486 86522
rect 142486 86470 142516 86522
rect 142540 86470 142550 86522
rect 142550 86470 142596 86522
rect 142620 86470 142666 86522
rect 142666 86470 142676 86522
rect 142700 86470 142730 86522
rect 142730 86470 142756 86522
rect 142460 86468 142516 86470
rect 142540 86468 142596 86470
rect 142620 86468 142676 86470
rect 142700 86468 142756 86470
rect 142460 85434 142516 85436
rect 142540 85434 142596 85436
rect 142620 85434 142676 85436
rect 142700 85434 142756 85436
rect 142460 85382 142486 85434
rect 142486 85382 142516 85434
rect 142540 85382 142550 85434
rect 142550 85382 142596 85434
rect 142620 85382 142666 85434
rect 142666 85382 142676 85434
rect 142700 85382 142730 85434
rect 142730 85382 142756 85434
rect 142460 85380 142516 85382
rect 142540 85380 142596 85382
rect 142620 85380 142676 85382
rect 142700 85380 142756 85382
rect 142460 84346 142516 84348
rect 142540 84346 142596 84348
rect 142620 84346 142676 84348
rect 142700 84346 142756 84348
rect 142460 84294 142486 84346
rect 142486 84294 142516 84346
rect 142540 84294 142550 84346
rect 142550 84294 142596 84346
rect 142620 84294 142666 84346
rect 142666 84294 142676 84346
rect 142700 84294 142730 84346
rect 142730 84294 142756 84346
rect 142460 84292 142516 84294
rect 142540 84292 142596 84294
rect 142620 84292 142676 84294
rect 142700 84292 142756 84294
rect 142460 83258 142516 83260
rect 142540 83258 142596 83260
rect 142620 83258 142676 83260
rect 142700 83258 142756 83260
rect 142460 83206 142486 83258
rect 142486 83206 142516 83258
rect 142540 83206 142550 83258
rect 142550 83206 142596 83258
rect 142620 83206 142666 83258
rect 142666 83206 142676 83258
rect 142700 83206 142730 83258
rect 142730 83206 142756 83258
rect 142460 83204 142516 83206
rect 142540 83204 142596 83206
rect 142620 83204 142676 83206
rect 142700 83204 142756 83206
rect 142460 82170 142516 82172
rect 142540 82170 142596 82172
rect 142620 82170 142676 82172
rect 142700 82170 142756 82172
rect 142460 82118 142486 82170
rect 142486 82118 142516 82170
rect 142540 82118 142550 82170
rect 142550 82118 142596 82170
rect 142620 82118 142666 82170
rect 142666 82118 142676 82170
rect 142700 82118 142730 82170
rect 142730 82118 142756 82170
rect 142460 82116 142516 82118
rect 142540 82116 142596 82118
rect 142620 82116 142676 82118
rect 142700 82116 142756 82118
rect 142460 81082 142516 81084
rect 142540 81082 142596 81084
rect 142620 81082 142676 81084
rect 142700 81082 142756 81084
rect 142460 81030 142486 81082
rect 142486 81030 142516 81082
rect 142540 81030 142550 81082
rect 142550 81030 142596 81082
rect 142620 81030 142666 81082
rect 142666 81030 142676 81082
rect 142700 81030 142730 81082
rect 142730 81030 142756 81082
rect 142460 81028 142516 81030
rect 142540 81028 142596 81030
rect 142620 81028 142676 81030
rect 142700 81028 142756 81030
rect 142460 79994 142516 79996
rect 142540 79994 142596 79996
rect 142620 79994 142676 79996
rect 142700 79994 142756 79996
rect 142460 79942 142486 79994
rect 142486 79942 142516 79994
rect 142540 79942 142550 79994
rect 142550 79942 142596 79994
rect 142620 79942 142666 79994
rect 142666 79942 142676 79994
rect 142700 79942 142730 79994
rect 142730 79942 142756 79994
rect 142460 79940 142516 79942
rect 142540 79940 142596 79942
rect 142620 79940 142676 79942
rect 142700 79940 142756 79942
rect 142460 78906 142516 78908
rect 142540 78906 142596 78908
rect 142620 78906 142676 78908
rect 142700 78906 142756 78908
rect 142460 78854 142486 78906
rect 142486 78854 142516 78906
rect 142540 78854 142550 78906
rect 142550 78854 142596 78906
rect 142620 78854 142666 78906
rect 142666 78854 142676 78906
rect 142700 78854 142730 78906
rect 142730 78854 142756 78906
rect 142460 78852 142516 78854
rect 142540 78852 142596 78854
rect 142620 78852 142676 78854
rect 142700 78852 142756 78854
rect 142460 77818 142516 77820
rect 142540 77818 142596 77820
rect 142620 77818 142676 77820
rect 142700 77818 142756 77820
rect 142460 77766 142486 77818
rect 142486 77766 142516 77818
rect 142540 77766 142550 77818
rect 142550 77766 142596 77818
rect 142620 77766 142666 77818
rect 142666 77766 142676 77818
rect 142700 77766 142730 77818
rect 142730 77766 142756 77818
rect 142460 77764 142516 77766
rect 142540 77764 142596 77766
rect 142620 77764 142676 77766
rect 142700 77764 142756 77766
rect 142460 76730 142516 76732
rect 142540 76730 142596 76732
rect 142620 76730 142676 76732
rect 142700 76730 142756 76732
rect 142460 76678 142486 76730
rect 142486 76678 142516 76730
rect 142540 76678 142550 76730
rect 142550 76678 142596 76730
rect 142620 76678 142666 76730
rect 142666 76678 142676 76730
rect 142700 76678 142730 76730
rect 142730 76678 142756 76730
rect 142460 76676 142516 76678
rect 142540 76676 142596 76678
rect 142620 76676 142676 76678
rect 142700 76676 142756 76678
rect 142460 75642 142516 75644
rect 142540 75642 142596 75644
rect 142620 75642 142676 75644
rect 142700 75642 142756 75644
rect 142460 75590 142486 75642
rect 142486 75590 142516 75642
rect 142540 75590 142550 75642
rect 142550 75590 142596 75642
rect 142620 75590 142666 75642
rect 142666 75590 142676 75642
rect 142700 75590 142730 75642
rect 142730 75590 142756 75642
rect 142460 75588 142516 75590
rect 142540 75588 142596 75590
rect 142620 75588 142676 75590
rect 142700 75588 142756 75590
rect 142460 74554 142516 74556
rect 142540 74554 142596 74556
rect 142620 74554 142676 74556
rect 142700 74554 142756 74556
rect 142460 74502 142486 74554
rect 142486 74502 142516 74554
rect 142540 74502 142550 74554
rect 142550 74502 142596 74554
rect 142620 74502 142666 74554
rect 142666 74502 142676 74554
rect 142700 74502 142730 74554
rect 142730 74502 142756 74554
rect 142460 74500 142516 74502
rect 142540 74500 142596 74502
rect 142620 74500 142676 74502
rect 142700 74500 142756 74502
rect 142460 73466 142516 73468
rect 142540 73466 142596 73468
rect 142620 73466 142676 73468
rect 142700 73466 142756 73468
rect 142460 73414 142486 73466
rect 142486 73414 142516 73466
rect 142540 73414 142550 73466
rect 142550 73414 142596 73466
rect 142620 73414 142666 73466
rect 142666 73414 142676 73466
rect 142700 73414 142730 73466
rect 142730 73414 142756 73466
rect 142460 73412 142516 73414
rect 142540 73412 142596 73414
rect 142620 73412 142676 73414
rect 142700 73412 142756 73414
rect 142460 72378 142516 72380
rect 142540 72378 142596 72380
rect 142620 72378 142676 72380
rect 142700 72378 142756 72380
rect 142460 72326 142486 72378
rect 142486 72326 142516 72378
rect 142540 72326 142550 72378
rect 142550 72326 142596 72378
rect 142620 72326 142666 72378
rect 142666 72326 142676 72378
rect 142700 72326 142730 72378
rect 142730 72326 142756 72378
rect 142460 72324 142516 72326
rect 142540 72324 142596 72326
rect 142620 72324 142676 72326
rect 142700 72324 142756 72326
rect 142460 71290 142516 71292
rect 142540 71290 142596 71292
rect 142620 71290 142676 71292
rect 142700 71290 142756 71292
rect 142460 71238 142486 71290
rect 142486 71238 142516 71290
rect 142540 71238 142550 71290
rect 142550 71238 142596 71290
rect 142620 71238 142666 71290
rect 142666 71238 142676 71290
rect 142700 71238 142730 71290
rect 142730 71238 142756 71290
rect 142460 71236 142516 71238
rect 142540 71236 142596 71238
rect 142620 71236 142676 71238
rect 142700 71236 142756 71238
rect 142460 70202 142516 70204
rect 142540 70202 142596 70204
rect 142620 70202 142676 70204
rect 142700 70202 142756 70204
rect 142460 70150 142486 70202
rect 142486 70150 142516 70202
rect 142540 70150 142550 70202
rect 142550 70150 142596 70202
rect 142620 70150 142666 70202
rect 142666 70150 142676 70202
rect 142700 70150 142730 70202
rect 142730 70150 142756 70202
rect 142460 70148 142516 70150
rect 142540 70148 142596 70150
rect 142620 70148 142676 70150
rect 142700 70148 142756 70150
rect 142460 69114 142516 69116
rect 142540 69114 142596 69116
rect 142620 69114 142676 69116
rect 142700 69114 142756 69116
rect 142460 69062 142486 69114
rect 142486 69062 142516 69114
rect 142540 69062 142550 69114
rect 142550 69062 142596 69114
rect 142620 69062 142666 69114
rect 142666 69062 142676 69114
rect 142700 69062 142730 69114
rect 142730 69062 142756 69114
rect 142460 69060 142516 69062
rect 142540 69060 142596 69062
rect 142620 69060 142676 69062
rect 142700 69060 142756 69062
rect 142460 68026 142516 68028
rect 142540 68026 142596 68028
rect 142620 68026 142676 68028
rect 142700 68026 142756 68028
rect 142460 67974 142486 68026
rect 142486 67974 142516 68026
rect 142540 67974 142550 68026
rect 142550 67974 142596 68026
rect 142620 67974 142666 68026
rect 142666 67974 142676 68026
rect 142700 67974 142730 68026
rect 142730 67974 142756 68026
rect 142460 67972 142516 67974
rect 142540 67972 142596 67974
rect 142620 67972 142676 67974
rect 142700 67972 142756 67974
rect 142460 66938 142516 66940
rect 142540 66938 142596 66940
rect 142620 66938 142676 66940
rect 142700 66938 142756 66940
rect 142460 66886 142486 66938
rect 142486 66886 142516 66938
rect 142540 66886 142550 66938
rect 142550 66886 142596 66938
rect 142620 66886 142666 66938
rect 142666 66886 142676 66938
rect 142700 66886 142730 66938
rect 142730 66886 142756 66938
rect 142460 66884 142516 66886
rect 142540 66884 142596 66886
rect 142620 66884 142676 66886
rect 142700 66884 142756 66886
rect 142460 65850 142516 65852
rect 142540 65850 142596 65852
rect 142620 65850 142676 65852
rect 142700 65850 142756 65852
rect 142460 65798 142486 65850
rect 142486 65798 142516 65850
rect 142540 65798 142550 65850
rect 142550 65798 142596 65850
rect 142620 65798 142666 65850
rect 142666 65798 142676 65850
rect 142700 65798 142730 65850
rect 142730 65798 142756 65850
rect 142460 65796 142516 65798
rect 142540 65796 142596 65798
rect 142620 65796 142676 65798
rect 142700 65796 142756 65798
rect 142460 64762 142516 64764
rect 142540 64762 142596 64764
rect 142620 64762 142676 64764
rect 142700 64762 142756 64764
rect 142460 64710 142486 64762
rect 142486 64710 142516 64762
rect 142540 64710 142550 64762
rect 142550 64710 142596 64762
rect 142620 64710 142666 64762
rect 142666 64710 142676 64762
rect 142700 64710 142730 64762
rect 142730 64710 142756 64762
rect 142460 64708 142516 64710
rect 142540 64708 142596 64710
rect 142620 64708 142676 64710
rect 142700 64708 142756 64710
rect 142460 63674 142516 63676
rect 142540 63674 142596 63676
rect 142620 63674 142676 63676
rect 142700 63674 142756 63676
rect 142460 63622 142486 63674
rect 142486 63622 142516 63674
rect 142540 63622 142550 63674
rect 142550 63622 142596 63674
rect 142620 63622 142666 63674
rect 142666 63622 142676 63674
rect 142700 63622 142730 63674
rect 142730 63622 142756 63674
rect 142460 63620 142516 63622
rect 142540 63620 142596 63622
rect 142620 63620 142676 63622
rect 142700 63620 142756 63622
rect 142460 62586 142516 62588
rect 142540 62586 142596 62588
rect 142620 62586 142676 62588
rect 142700 62586 142756 62588
rect 142460 62534 142486 62586
rect 142486 62534 142516 62586
rect 142540 62534 142550 62586
rect 142550 62534 142596 62586
rect 142620 62534 142666 62586
rect 142666 62534 142676 62586
rect 142700 62534 142730 62586
rect 142730 62534 142756 62586
rect 142460 62532 142516 62534
rect 142540 62532 142596 62534
rect 142620 62532 142676 62534
rect 142700 62532 142756 62534
rect 142460 61498 142516 61500
rect 142540 61498 142596 61500
rect 142620 61498 142676 61500
rect 142700 61498 142756 61500
rect 142460 61446 142486 61498
rect 142486 61446 142516 61498
rect 142540 61446 142550 61498
rect 142550 61446 142596 61498
rect 142620 61446 142666 61498
rect 142666 61446 142676 61498
rect 142700 61446 142730 61498
rect 142730 61446 142756 61498
rect 142460 61444 142516 61446
rect 142540 61444 142596 61446
rect 142620 61444 142676 61446
rect 142700 61444 142756 61446
rect 142460 60410 142516 60412
rect 142540 60410 142596 60412
rect 142620 60410 142676 60412
rect 142700 60410 142756 60412
rect 142460 60358 142486 60410
rect 142486 60358 142516 60410
rect 142540 60358 142550 60410
rect 142550 60358 142596 60410
rect 142620 60358 142666 60410
rect 142666 60358 142676 60410
rect 142700 60358 142730 60410
rect 142730 60358 142756 60410
rect 142460 60356 142516 60358
rect 142540 60356 142596 60358
rect 142620 60356 142676 60358
rect 142700 60356 142756 60358
rect 142460 59322 142516 59324
rect 142540 59322 142596 59324
rect 142620 59322 142676 59324
rect 142700 59322 142756 59324
rect 142460 59270 142486 59322
rect 142486 59270 142516 59322
rect 142540 59270 142550 59322
rect 142550 59270 142596 59322
rect 142620 59270 142666 59322
rect 142666 59270 142676 59322
rect 142700 59270 142730 59322
rect 142730 59270 142756 59322
rect 142460 59268 142516 59270
rect 142540 59268 142596 59270
rect 142620 59268 142676 59270
rect 142700 59268 142756 59270
rect 142460 58234 142516 58236
rect 142540 58234 142596 58236
rect 142620 58234 142676 58236
rect 142700 58234 142756 58236
rect 142460 58182 142486 58234
rect 142486 58182 142516 58234
rect 142540 58182 142550 58234
rect 142550 58182 142596 58234
rect 142620 58182 142666 58234
rect 142666 58182 142676 58234
rect 142700 58182 142730 58234
rect 142730 58182 142756 58234
rect 142460 58180 142516 58182
rect 142540 58180 142596 58182
rect 142620 58180 142676 58182
rect 142700 58180 142756 58182
rect 142460 57146 142516 57148
rect 142540 57146 142596 57148
rect 142620 57146 142676 57148
rect 142700 57146 142756 57148
rect 142460 57094 142486 57146
rect 142486 57094 142516 57146
rect 142540 57094 142550 57146
rect 142550 57094 142596 57146
rect 142620 57094 142666 57146
rect 142666 57094 142676 57146
rect 142700 57094 142730 57146
rect 142730 57094 142756 57146
rect 142460 57092 142516 57094
rect 142540 57092 142596 57094
rect 142620 57092 142676 57094
rect 142700 57092 142756 57094
rect 142460 56058 142516 56060
rect 142540 56058 142596 56060
rect 142620 56058 142676 56060
rect 142700 56058 142756 56060
rect 142460 56006 142486 56058
rect 142486 56006 142516 56058
rect 142540 56006 142550 56058
rect 142550 56006 142596 56058
rect 142620 56006 142666 56058
rect 142666 56006 142676 56058
rect 142700 56006 142730 56058
rect 142730 56006 142756 56058
rect 142460 56004 142516 56006
rect 142540 56004 142596 56006
rect 142620 56004 142676 56006
rect 142700 56004 142756 56006
rect 142460 54970 142516 54972
rect 142540 54970 142596 54972
rect 142620 54970 142676 54972
rect 142700 54970 142756 54972
rect 142460 54918 142486 54970
rect 142486 54918 142516 54970
rect 142540 54918 142550 54970
rect 142550 54918 142596 54970
rect 142620 54918 142666 54970
rect 142666 54918 142676 54970
rect 142700 54918 142730 54970
rect 142730 54918 142756 54970
rect 142460 54916 142516 54918
rect 142540 54916 142596 54918
rect 142620 54916 142676 54918
rect 142700 54916 142756 54918
rect 142460 53882 142516 53884
rect 142540 53882 142596 53884
rect 142620 53882 142676 53884
rect 142700 53882 142756 53884
rect 142460 53830 142486 53882
rect 142486 53830 142516 53882
rect 142540 53830 142550 53882
rect 142550 53830 142596 53882
rect 142620 53830 142666 53882
rect 142666 53830 142676 53882
rect 142700 53830 142730 53882
rect 142730 53830 142756 53882
rect 142460 53828 142516 53830
rect 142540 53828 142596 53830
rect 142620 53828 142676 53830
rect 142700 53828 142756 53830
rect 142460 52794 142516 52796
rect 142540 52794 142596 52796
rect 142620 52794 142676 52796
rect 142700 52794 142756 52796
rect 142460 52742 142486 52794
rect 142486 52742 142516 52794
rect 142540 52742 142550 52794
rect 142550 52742 142596 52794
rect 142620 52742 142666 52794
rect 142666 52742 142676 52794
rect 142700 52742 142730 52794
rect 142730 52742 142756 52794
rect 142460 52740 142516 52742
rect 142540 52740 142596 52742
rect 142620 52740 142676 52742
rect 142700 52740 142756 52742
rect 142460 51706 142516 51708
rect 142540 51706 142596 51708
rect 142620 51706 142676 51708
rect 142700 51706 142756 51708
rect 142460 51654 142486 51706
rect 142486 51654 142516 51706
rect 142540 51654 142550 51706
rect 142550 51654 142596 51706
rect 142620 51654 142666 51706
rect 142666 51654 142676 51706
rect 142700 51654 142730 51706
rect 142730 51654 142756 51706
rect 142460 51652 142516 51654
rect 142540 51652 142596 51654
rect 142620 51652 142676 51654
rect 142700 51652 142756 51654
rect 142460 50618 142516 50620
rect 142540 50618 142596 50620
rect 142620 50618 142676 50620
rect 142700 50618 142756 50620
rect 142460 50566 142486 50618
rect 142486 50566 142516 50618
rect 142540 50566 142550 50618
rect 142550 50566 142596 50618
rect 142620 50566 142666 50618
rect 142666 50566 142676 50618
rect 142700 50566 142730 50618
rect 142730 50566 142756 50618
rect 142460 50564 142516 50566
rect 142540 50564 142596 50566
rect 142620 50564 142676 50566
rect 142700 50564 142756 50566
rect 142460 49530 142516 49532
rect 142540 49530 142596 49532
rect 142620 49530 142676 49532
rect 142700 49530 142756 49532
rect 142460 49478 142486 49530
rect 142486 49478 142516 49530
rect 142540 49478 142550 49530
rect 142550 49478 142596 49530
rect 142620 49478 142666 49530
rect 142666 49478 142676 49530
rect 142700 49478 142730 49530
rect 142730 49478 142756 49530
rect 142460 49476 142516 49478
rect 142540 49476 142596 49478
rect 142620 49476 142676 49478
rect 142700 49476 142756 49478
rect 142460 48442 142516 48444
rect 142540 48442 142596 48444
rect 142620 48442 142676 48444
rect 142700 48442 142756 48444
rect 142460 48390 142486 48442
rect 142486 48390 142516 48442
rect 142540 48390 142550 48442
rect 142550 48390 142596 48442
rect 142620 48390 142666 48442
rect 142666 48390 142676 48442
rect 142700 48390 142730 48442
rect 142730 48390 142756 48442
rect 142460 48388 142516 48390
rect 142540 48388 142596 48390
rect 142620 48388 142676 48390
rect 142700 48388 142756 48390
rect 142460 47354 142516 47356
rect 142540 47354 142596 47356
rect 142620 47354 142676 47356
rect 142700 47354 142756 47356
rect 142460 47302 142486 47354
rect 142486 47302 142516 47354
rect 142540 47302 142550 47354
rect 142550 47302 142596 47354
rect 142620 47302 142666 47354
rect 142666 47302 142676 47354
rect 142700 47302 142730 47354
rect 142730 47302 142756 47354
rect 142460 47300 142516 47302
rect 142540 47300 142596 47302
rect 142620 47300 142676 47302
rect 142700 47300 142756 47302
rect 142460 46266 142516 46268
rect 142540 46266 142596 46268
rect 142620 46266 142676 46268
rect 142700 46266 142756 46268
rect 142460 46214 142486 46266
rect 142486 46214 142516 46266
rect 142540 46214 142550 46266
rect 142550 46214 142596 46266
rect 142620 46214 142666 46266
rect 142666 46214 142676 46266
rect 142700 46214 142730 46266
rect 142730 46214 142756 46266
rect 142460 46212 142516 46214
rect 142540 46212 142596 46214
rect 142620 46212 142676 46214
rect 142700 46212 142756 46214
rect 142460 45178 142516 45180
rect 142540 45178 142596 45180
rect 142620 45178 142676 45180
rect 142700 45178 142756 45180
rect 142460 45126 142486 45178
rect 142486 45126 142516 45178
rect 142540 45126 142550 45178
rect 142550 45126 142596 45178
rect 142620 45126 142666 45178
rect 142666 45126 142676 45178
rect 142700 45126 142730 45178
rect 142730 45126 142756 45178
rect 142460 45124 142516 45126
rect 142540 45124 142596 45126
rect 142620 45124 142676 45126
rect 142700 45124 142756 45126
rect 142460 44090 142516 44092
rect 142540 44090 142596 44092
rect 142620 44090 142676 44092
rect 142700 44090 142756 44092
rect 142460 44038 142486 44090
rect 142486 44038 142516 44090
rect 142540 44038 142550 44090
rect 142550 44038 142596 44090
rect 142620 44038 142666 44090
rect 142666 44038 142676 44090
rect 142700 44038 142730 44090
rect 142730 44038 142756 44090
rect 142460 44036 142516 44038
rect 142540 44036 142596 44038
rect 142620 44036 142676 44038
rect 142700 44036 142756 44038
rect 142460 43002 142516 43004
rect 142540 43002 142596 43004
rect 142620 43002 142676 43004
rect 142700 43002 142756 43004
rect 142460 42950 142486 43002
rect 142486 42950 142516 43002
rect 142540 42950 142550 43002
rect 142550 42950 142596 43002
rect 142620 42950 142666 43002
rect 142666 42950 142676 43002
rect 142700 42950 142730 43002
rect 142730 42950 142756 43002
rect 142460 42948 142516 42950
rect 142540 42948 142596 42950
rect 142620 42948 142676 42950
rect 142700 42948 142756 42950
rect 142460 41914 142516 41916
rect 142540 41914 142596 41916
rect 142620 41914 142676 41916
rect 142700 41914 142756 41916
rect 142460 41862 142486 41914
rect 142486 41862 142516 41914
rect 142540 41862 142550 41914
rect 142550 41862 142596 41914
rect 142620 41862 142666 41914
rect 142666 41862 142676 41914
rect 142700 41862 142730 41914
rect 142730 41862 142756 41914
rect 142460 41860 142516 41862
rect 142540 41860 142596 41862
rect 142620 41860 142676 41862
rect 142700 41860 142756 41862
rect 142460 40826 142516 40828
rect 142540 40826 142596 40828
rect 142620 40826 142676 40828
rect 142700 40826 142756 40828
rect 142460 40774 142486 40826
rect 142486 40774 142516 40826
rect 142540 40774 142550 40826
rect 142550 40774 142596 40826
rect 142620 40774 142666 40826
rect 142666 40774 142676 40826
rect 142700 40774 142730 40826
rect 142730 40774 142756 40826
rect 142460 40772 142516 40774
rect 142540 40772 142596 40774
rect 142620 40772 142676 40774
rect 142700 40772 142756 40774
rect 142460 39738 142516 39740
rect 142540 39738 142596 39740
rect 142620 39738 142676 39740
rect 142700 39738 142756 39740
rect 142460 39686 142486 39738
rect 142486 39686 142516 39738
rect 142540 39686 142550 39738
rect 142550 39686 142596 39738
rect 142620 39686 142666 39738
rect 142666 39686 142676 39738
rect 142700 39686 142730 39738
rect 142730 39686 142756 39738
rect 142460 39684 142516 39686
rect 142540 39684 142596 39686
rect 142620 39684 142676 39686
rect 142700 39684 142756 39686
rect 142460 38650 142516 38652
rect 142540 38650 142596 38652
rect 142620 38650 142676 38652
rect 142700 38650 142756 38652
rect 142460 38598 142486 38650
rect 142486 38598 142516 38650
rect 142540 38598 142550 38650
rect 142550 38598 142596 38650
rect 142620 38598 142666 38650
rect 142666 38598 142676 38650
rect 142700 38598 142730 38650
rect 142730 38598 142756 38650
rect 142460 38596 142516 38598
rect 142540 38596 142596 38598
rect 142620 38596 142676 38598
rect 142700 38596 142756 38598
rect 142460 37562 142516 37564
rect 142540 37562 142596 37564
rect 142620 37562 142676 37564
rect 142700 37562 142756 37564
rect 142460 37510 142486 37562
rect 142486 37510 142516 37562
rect 142540 37510 142550 37562
rect 142550 37510 142596 37562
rect 142620 37510 142666 37562
rect 142666 37510 142676 37562
rect 142700 37510 142730 37562
rect 142730 37510 142756 37562
rect 142460 37508 142516 37510
rect 142540 37508 142596 37510
rect 142620 37508 142676 37510
rect 142700 37508 142756 37510
rect 142460 36474 142516 36476
rect 142540 36474 142596 36476
rect 142620 36474 142676 36476
rect 142700 36474 142756 36476
rect 142460 36422 142486 36474
rect 142486 36422 142516 36474
rect 142540 36422 142550 36474
rect 142550 36422 142596 36474
rect 142620 36422 142666 36474
rect 142666 36422 142676 36474
rect 142700 36422 142730 36474
rect 142730 36422 142756 36474
rect 142460 36420 142516 36422
rect 142540 36420 142596 36422
rect 142620 36420 142676 36422
rect 142700 36420 142756 36422
rect 142460 35386 142516 35388
rect 142540 35386 142596 35388
rect 142620 35386 142676 35388
rect 142700 35386 142756 35388
rect 142460 35334 142486 35386
rect 142486 35334 142516 35386
rect 142540 35334 142550 35386
rect 142550 35334 142596 35386
rect 142620 35334 142666 35386
rect 142666 35334 142676 35386
rect 142700 35334 142730 35386
rect 142730 35334 142756 35386
rect 142460 35332 142516 35334
rect 142540 35332 142596 35334
rect 142620 35332 142676 35334
rect 142700 35332 142756 35334
rect 142460 34298 142516 34300
rect 142540 34298 142596 34300
rect 142620 34298 142676 34300
rect 142700 34298 142756 34300
rect 142460 34246 142486 34298
rect 142486 34246 142516 34298
rect 142540 34246 142550 34298
rect 142550 34246 142596 34298
rect 142620 34246 142666 34298
rect 142666 34246 142676 34298
rect 142700 34246 142730 34298
rect 142730 34246 142756 34298
rect 142460 34244 142516 34246
rect 142540 34244 142596 34246
rect 142620 34244 142676 34246
rect 142700 34244 142756 34246
rect 142460 33210 142516 33212
rect 142540 33210 142596 33212
rect 142620 33210 142676 33212
rect 142700 33210 142756 33212
rect 142460 33158 142486 33210
rect 142486 33158 142516 33210
rect 142540 33158 142550 33210
rect 142550 33158 142596 33210
rect 142620 33158 142666 33210
rect 142666 33158 142676 33210
rect 142700 33158 142730 33210
rect 142730 33158 142756 33210
rect 142460 33156 142516 33158
rect 142540 33156 142596 33158
rect 142620 33156 142676 33158
rect 142700 33156 142756 33158
rect 142460 32122 142516 32124
rect 142540 32122 142596 32124
rect 142620 32122 142676 32124
rect 142700 32122 142756 32124
rect 142460 32070 142486 32122
rect 142486 32070 142516 32122
rect 142540 32070 142550 32122
rect 142550 32070 142596 32122
rect 142620 32070 142666 32122
rect 142666 32070 142676 32122
rect 142700 32070 142730 32122
rect 142730 32070 142756 32122
rect 142460 32068 142516 32070
rect 142540 32068 142596 32070
rect 142620 32068 142676 32070
rect 142700 32068 142756 32070
rect 142460 31034 142516 31036
rect 142540 31034 142596 31036
rect 142620 31034 142676 31036
rect 142700 31034 142756 31036
rect 142460 30982 142486 31034
rect 142486 30982 142516 31034
rect 142540 30982 142550 31034
rect 142550 30982 142596 31034
rect 142620 30982 142666 31034
rect 142666 30982 142676 31034
rect 142700 30982 142730 31034
rect 142730 30982 142756 31034
rect 142460 30980 142516 30982
rect 142540 30980 142596 30982
rect 142620 30980 142676 30982
rect 142700 30980 142756 30982
rect 142460 29946 142516 29948
rect 142540 29946 142596 29948
rect 142620 29946 142676 29948
rect 142700 29946 142756 29948
rect 142460 29894 142486 29946
rect 142486 29894 142516 29946
rect 142540 29894 142550 29946
rect 142550 29894 142596 29946
rect 142620 29894 142666 29946
rect 142666 29894 142676 29946
rect 142700 29894 142730 29946
rect 142730 29894 142756 29946
rect 142460 29892 142516 29894
rect 142540 29892 142596 29894
rect 142620 29892 142676 29894
rect 142700 29892 142756 29894
rect 142460 28858 142516 28860
rect 142540 28858 142596 28860
rect 142620 28858 142676 28860
rect 142700 28858 142756 28860
rect 142460 28806 142486 28858
rect 142486 28806 142516 28858
rect 142540 28806 142550 28858
rect 142550 28806 142596 28858
rect 142620 28806 142666 28858
rect 142666 28806 142676 28858
rect 142700 28806 142730 28858
rect 142730 28806 142756 28858
rect 142460 28804 142516 28806
rect 142540 28804 142596 28806
rect 142620 28804 142676 28806
rect 142700 28804 142756 28806
rect 142460 27770 142516 27772
rect 142540 27770 142596 27772
rect 142620 27770 142676 27772
rect 142700 27770 142756 27772
rect 142460 27718 142486 27770
rect 142486 27718 142516 27770
rect 142540 27718 142550 27770
rect 142550 27718 142596 27770
rect 142620 27718 142666 27770
rect 142666 27718 142676 27770
rect 142700 27718 142730 27770
rect 142730 27718 142756 27770
rect 142460 27716 142516 27718
rect 142540 27716 142596 27718
rect 142620 27716 142676 27718
rect 142700 27716 142756 27718
rect 142460 26682 142516 26684
rect 142540 26682 142596 26684
rect 142620 26682 142676 26684
rect 142700 26682 142756 26684
rect 142460 26630 142486 26682
rect 142486 26630 142516 26682
rect 142540 26630 142550 26682
rect 142550 26630 142596 26682
rect 142620 26630 142666 26682
rect 142666 26630 142676 26682
rect 142700 26630 142730 26682
rect 142730 26630 142756 26682
rect 142460 26628 142516 26630
rect 142540 26628 142596 26630
rect 142620 26628 142676 26630
rect 142700 26628 142756 26630
rect 142460 25594 142516 25596
rect 142540 25594 142596 25596
rect 142620 25594 142676 25596
rect 142700 25594 142756 25596
rect 142460 25542 142486 25594
rect 142486 25542 142516 25594
rect 142540 25542 142550 25594
rect 142550 25542 142596 25594
rect 142620 25542 142666 25594
rect 142666 25542 142676 25594
rect 142700 25542 142730 25594
rect 142730 25542 142756 25594
rect 142460 25540 142516 25542
rect 142540 25540 142596 25542
rect 142620 25540 142676 25542
rect 142700 25540 142756 25542
rect 142460 24506 142516 24508
rect 142540 24506 142596 24508
rect 142620 24506 142676 24508
rect 142700 24506 142756 24508
rect 142460 24454 142486 24506
rect 142486 24454 142516 24506
rect 142540 24454 142550 24506
rect 142550 24454 142596 24506
rect 142620 24454 142666 24506
rect 142666 24454 142676 24506
rect 142700 24454 142730 24506
rect 142730 24454 142756 24506
rect 142460 24452 142516 24454
rect 142540 24452 142596 24454
rect 142620 24452 142676 24454
rect 142700 24452 142756 24454
rect 142460 23418 142516 23420
rect 142540 23418 142596 23420
rect 142620 23418 142676 23420
rect 142700 23418 142756 23420
rect 142460 23366 142486 23418
rect 142486 23366 142516 23418
rect 142540 23366 142550 23418
rect 142550 23366 142596 23418
rect 142620 23366 142666 23418
rect 142666 23366 142676 23418
rect 142700 23366 142730 23418
rect 142730 23366 142756 23418
rect 142460 23364 142516 23366
rect 142540 23364 142596 23366
rect 142620 23364 142676 23366
rect 142700 23364 142756 23366
rect 142460 22330 142516 22332
rect 142540 22330 142596 22332
rect 142620 22330 142676 22332
rect 142700 22330 142756 22332
rect 142460 22278 142486 22330
rect 142486 22278 142516 22330
rect 142540 22278 142550 22330
rect 142550 22278 142596 22330
rect 142620 22278 142666 22330
rect 142666 22278 142676 22330
rect 142700 22278 142730 22330
rect 142730 22278 142756 22330
rect 142460 22276 142516 22278
rect 142540 22276 142596 22278
rect 142620 22276 142676 22278
rect 142700 22276 142756 22278
rect 142460 21242 142516 21244
rect 142540 21242 142596 21244
rect 142620 21242 142676 21244
rect 142700 21242 142756 21244
rect 142460 21190 142486 21242
rect 142486 21190 142516 21242
rect 142540 21190 142550 21242
rect 142550 21190 142596 21242
rect 142620 21190 142666 21242
rect 142666 21190 142676 21242
rect 142700 21190 142730 21242
rect 142730 21190 142756 21242
rect 142460 21188 142516 21190
rect 142540 21188 142596 21190
rect 142620 21188 142676 21190
rect 142700 21188 142756 21190
rect 142460 20154 142516 20156
rect 142540 20154 142596 20156
rect 142620 20154 142676 20156
rect 142700 20154 142756 20156
rect 142460 20102 142486 20154
rect 142486 20102 142516 20154
rect 142540 20102 142550 20154
rect 142550 20102 142596 20154
rect 142620 20102 142666 20154
rect 142666 20102 142676 20154
rect 142700 20102 142730 20154
rect 142730 20102 142756 20154
rect 142460 20100 142516 20102
rect 142540 20100 142596 20102
rect 142620 20100 142676 20102
rect 142700 20100 142756 20102
rect 81020 19066 81076 19068
rect 81100 19066 81156 19068
rect 81180 19066 81236 19068
rect 81260 19066 81316 19068
rect 81020 19014 81046 19066
rect 81046 19014 81076 19066
rect 81100 19014 81110 19066
rect 81110 19014 81156 19066
rect 81180 19014 81226 19066
rect 81226 19014 81236 19066
rect 81260 19014 81290 19066
rect 81290 19014 81316 19066
rect 81020 19012 81076 19014
rect 81100 19012 81156 19014
rect 81180 19012 81236 19014
rect 81260 19012 81316 19014
rect 111740 19066 111796 19068
rect 111820 19066 111876 19068
rect 111900 19066 111956 19068
rect 111980 19066 112036 19068
rect 111740 19014 111766 19066
rect 111766 19014 111796 19066
rect 111820 19014 111830 19066
rect 111830 19014 111876 19066
rect 111900 19014 111946 19066
rect 111946 19014 111956 19066
rect 111980 19014 112010 19066
rect 112010 19014 112036 19066
rect 111740 19012 111796 19014
rect 111820 19012 111876 19014
rect 111900 19012 111956 19014
rect 111980 19012 112036 19014
rect 142460 19066 142516 19068
rect 142540 19066 142596 19068
rect 142620 19066 142676 19068
rect 142700 19066 142756 19068
rect 142460 19014 142486 19066
rect 142486 19014 142516 19066
rect 142540 19014 142550 19066
rect 142550 19014 142596 19066
rect 142620 19014 142666 19066
rect 142666 19014 142676 19066
rect 142700 19014 142730 19066
rect 142730 19014 142756 19066
rect 142460 19012 142516 19014
rect 142540 19012 142596 19014
rect 142620 19012 142676 19014
rect 142700 19012 142756 19014
rect 157820 116442 157876 116444
rect 157900 116442 157956 116444
rect 157980 116442 158036 116444
rect 158060 116442 158116 116444
rect 157820 116390 157846 116442
rect 157846 116390 157876 116442
rect 157900 116390 157910 116442
rect 157910 116390 157956 116442
rect 157980 116390 158026 116442
rect 158026 116390 158036 116442
rect 158060 116390 158090 116442
rect 158090 116390 158116 116442
rect 157820 116388 157876 116390
rect 157900 116388 157956 116390
rect 157980 116388 158036 116390
rect 158060 116388 158116 116390
rect 173180 116986 173236 116988
rect 173260 116986 173316 116988
rect 173340 116986 173396 116988
rect 173420 116986 173476 116988
rect 173180 116934 173206 116986
rect 173206 116934 173236 116986
rect 173260 116934 173270 116986
rect 173270 116934 173316 116986
rect 173340 116934 173386 116986
rect 173386 116934 173396 116986
rect 173420 116934 173450 116986
rect 173450 116934 173476 116986
rect 173180 116932 173236 116934
rect 173260 116932 173316 116934
rect 173340 116932 173396 116934
rect 173420 116932 173476 116934
rect 173180 115898 173236 115900
rect 173260 115898 173316 115900
rect 173340 115898 173396 115900
rect 173420 115898 173476 115900
rect 173180 115846 173206 115898
rect 173206 115846 173236 115898
rect 173260 115846 173270 115898
rect 173270 115846 173316 115898
rect 173340 115846 173386 115898
rect 173386 115846 173396 115898
rect 173420 115846 173450 115898
rect 173450 115846 173476 115898
rect 173180 115844 173236 115846
rect 173260 115844 173316 115846
rect 173340 115844 173396 115846
rect 173420 115844 173476 115846
rect 157820 115354 157876 115356
rect 157900 115354 157956 115356
rect 157980 115354 158036 115356
rect 158060 115354 158116 115356
rect 157820 115302 157846 115354
rect 157846 115302 157876 115354
rect 157900 115302 157910 115354
rect 157910 115302 157956 115354
rect 157980 115302 158026 115354
rect 158026 115302 158036 115354
rect 158060 115302 158090 115354
rect 158090 115302 158116 115354
rect 157820 115300 157876 115302
rect 157900 115300 157956 115302
rect 157980 115300 158036 115302
rect 158060 115300 158116 115302
rect 173180 114810 173236 114812
rect 173260 114810 173316 114812
rect 173340 114810 173396 114812
rect 173420 114810 173476 114812
rect 173180 114758 173206 114810
rect 173206 114758 173236 114810
rect 173260 114758 173270 114810
rect 173270 114758 173316 114810
rect 173340 114758 173386 114810
rect 173386 114758 173396 114810
rect 173420 114758 173450 114810
rect 173450 114758 173476 114810
rect 173180 114756 173236 114758
rect 173260 114756 173316 114758
rect 173340 114756 173396 114758
rect 173420 114756 173476 114758
rect 157820 114266 157876 114268
rect 157900 114266 157956 114268
rect 157980 114266 158036 114268
rect 158060 114266 158116 114268
rect 157820 114214 157846 114266
rect 157846 114214 157876 114266
rect 157900 114214 157910 114266
rect 157910 114214 157956 114266
rect 157980 114214 158026 114266
rect 158026 114214 158036 114266
rect 158060 114214 158090 114266
rect 158090 114214 158116 114266
rect 157820 114212 157876 114214
rect 157900 114212 157956 114214
rect 157980 114212 158036 114214
rect 158060 114212 158116 114214
rect 173180 113722 173236 113724
rect 173260 113722 173316 113724
rect 173340 113722 173396 113724
rect 173420 113722 173476 113724
rect 173180 113670 173206 113722
rect 173206 113670 173236 113722
rect 173260 113670 173270 113722
rect 173270 113670 173316 113722
rect 173340 113670 173386 113722
rect 173386 113670 173396 113722
rect 173420 113670 173450 113722
rect 173450 113670 173476 113722
rect 173180 113668 173236 113670
rect 173260 113668 173316 113670
rect 173340 113668 173396 113670
rect 173420 113668 173476 113670
rect 157820 113178 157876 113180
rect 157900 113178 157956 113180
rect 157980 113178 158036 113180
rect 158060 113178 158116 113180
rect 157820 113126 157846 113178
rect 157846 113126 157876 113178
rect 157900 113126 157910 113178
rect 157910 113126 157956 113178
rect 157980 113126 158026 113178
rect 158026 113126 158036 113178
rect 158060 113126 158090 113178
rect 158090 113126 158116 113178
rect 157820 113124 157876 113126
rect 157900 113124 157956 113126
rect 157980 113124 158036 113126
rect 158060 113124 158116 113126
rect 173180 112634 173236 112636
rect 173260 112634 173316 112636
rect 173340 112634 173396 112636
rect 173420 112634 173476 112636
rect 173180 112582 173206 112634
rect 173206 112582 173236 112634
rect 173260 112582 173270 112634
rect 173270 112582 173316 112634
rect 173340 112582 173386 112634
rect 173386 112582 173396 112634
rect 173420 112582 173450 112634
rect 173450 112582 173476 112634
rect 173180 112580 173236 112582
rect 173260 112580 173316 112582
rect 173340 112580 173396 112582
rect 173420 112580 173476 112582
rect 157820 112090 157876 112092
rect 157900 112090 157956 112092
rect 157980 112090 158036 112092
rect 158060 112090 158116 112092
rect 157820 112038 157846 112090
rect 157846 112038 157876 112090
rect 157900 112038 157910 112090
rect 157910 112038 157956 112090
rect 157980 112038 158026 112090
rect 158026 112038 158036 112090
rect 158060 112038 158090 112090
rect 158090 112038 158116 112090
rect 157820 112036 157876 112038
rect 157900 112036 157956 112038
rect 157980 112036 158036 112038
rect 158060 112036 158116 112038
rect 173180 111546 173236 111548
rect 173260 111546 173316 111548
rect 173340 111546 173396 111548
rect 173420 111546 173476 111548
rect 173180 111494 173206 111546
rect 173206 111494 173236 111546
rect 173260 111494 173270 111546
rect 173270 111494 173316 111546
rect 173340 111494 173386 111546
rect 173386 111494 173396 111546
rect 173420 111494 173450 111546
rect 173450 111494 173476 111546
rect 173180 111492 173236 111494
rect 173260 111492 173316 111494
rect 173340 111492 173396 111494
rect 173420 111492 173476 111494
rect 157820 111002 157876 111004
rect 157900 111002 157956 111004
rect 157980 111002 158036 111004
rect 158060 111002 158116 111004
rect 157820 110950 157846 111002
rect 157846 110950 157876 111002
rect 157900 110950 157910 111002
rect 157910 110950 157956 111002
rect 157980 110950 158026 111002
rect 158026 110950 158036 111002
rect 158060 110950 158090 111002
rect 158090 110950 158116 111002
rect 157820 110948 157876 110950
rect 157900 110948 157956 110950
rect 157980 110948 158036 110950
rect 158060 110948 158116 110950
rect 173180 110458 173236 110460
rect 173260 110458 173316 110460
rect 173340 110458 173396 110460
rect 173420 110458 173476 110460
rect 173180 110406 173206 110458
rect 173206 110406 173236 110458
rect 173260 110406 173270 110458
rect 173270 110406 173316 110458
rect 173340 110406 173386 110458
rect 173386 110406 173396 110458
rect 173420 110406 173450 110458
rect 173450 110406 173476 110458
rect 173180 110404 173236 110406
rect 173260 110404 173316 110406
rect 173340 110404 173396 110406
rect 173420 110404 173476 110406
rect 157820 109914 157876 109916
rect 157900 109914 157956 109916
rect 157980 109914 158036 109916
rect 158060 109914 158116 109916
rect 157820 109862 157846 109914
rect 157846 109862 157876 109914
rect 157900 109862 157910 109914
rect 157910 109862 157956 109914
rect 157980 109862 158026 109914
rect 158026 109862 158036 109914
rect 158060 109862 158090 109914
rect 158090 109862 158116 109914
rect 157820 109860 157876 109862
rect 157900 109860 157956 109862
rect 157980 109860 158036 109862
rect 158060 109860 158116 109862
rect 173180 109370 173236 109372
rect 173260 109370 173316 109372
rect 173340 109370 173396 109372
rect 173420 109370 173476 109372
rect 173180 109318 173206 109370
rect 173206 109318 173236 109370
rect 173260 109318 173270 109370
rect 173270 109318 173316 109370
rect 173340 109318 173386 109370
rect 173386 109318 173396 109370
rect 173420 109318 173450 109370
rect 173450 109318 173476 109370
rect 173180 109316 173236 109318
rect 173260 109316 173316 109318
rect 173340 109316 173396 109318
rect 173420 109316 173476 109318
rect 157820 108826 157876 108828
rect 157900 108826 157956 108828
rect 157980 108826 158036 108828
rect 158060 108826 158116 108828
rect 157820 108774 157846 108826
rect 157846 108774 157876 108826
rect 157900 108774 157910 108826
rect 157910 108774 157956 108826
rect 157980 108774 158026 108826
rect 158026 108774 158036 108826
rect 158060 108774 158090 108826
rect 158090 108774 158116 108826
rect 157820 108772 157876 108774
rect 157900 108772 157956 108774
rect 157980 108772 158036 108774
rect 158060 108772 158116 108774
rect 173180 108282 173236 108284
rect 173260 108282 173316 108284
rect 173340 108282 173396 108284
rect 173420 108282 173476 108284
rect 173180 108230 173206 108282
rect 173206 108230 173236 108282
rect 173260 108230 173270 108282
rect 173270 108230 173316 108282
rect 173340 108230 173386 108282
rect 173386 108230 173396 108282
rect 173420 108230 173450 108282
rect 173450 108230 173476 108282
rect 173180 108228 173236 108230
rect 173260 108228 173316 108230
rect 173340 108228 173396 108230
rect 173420 108228 173476 108230
rect 157820 107738 157876 107740
rect 157900 107738 157956 107740
rect 157980 107738 158036 107740
rect 158060 107738 158116 107740
rect 157820 107686 157846 107738
rect 157846 107686 157876 107738
rect 157900 107686 157910 107738
rect 157910 107686 157956 107738
rect 157980 107686 158026 107738
rect 158026 107686 158036 107738
rect 158060 107686 158090 107738
rect 158090 107686 158116 107738
rect 157820 107684 157876 107686
rect 157900 107684 157956 107686
rect 157980 107684 158036 107686
rect 158060 107684 158116 107686
rect 173180 107194 173236 107196
rect 173260 107194 173316 107196
rect 173340 107194 173396 107196
rect 173420 107194 173476 107196
rect 173180 107142 173206 107194
rect 173206 107142 173236 107194
rect 173260 107142 173270 107194
rect 173270 107142 173316 107194
rect 173340 107142 173386 107194
rect 173386 107142 173396 107194
rect 173420 107142 173450 107194
rect 173450 107142 173476 107194
rect 173180 107140 173236 107142
rect 173260 107140 173316 107142
rect 173340 107140 173396 107142
rect 173420 107140 173476 107142
rect 157820 106650 157876 106652
rect 157900 106650 157956 106652
rect 157980 106650 158036 106652
rect 158060 106650 158116 106652
rect 157820 106598 157846 106650
rect 157846 106598 157876 106650
rect 157900 106598 157910 106650
rect 157910 106598 157956 106650
rect 157980 106598 158026 106650
rect 158026 106598 158036 106650
rect 158060 106598 158090 106650
rect 158090 106598 158116 106650
rect 157820 106596 157876 106598
rect 157900 106596 157956 106598
rect 157980 106596 158036 106598
rect 158060 106596 158116 106598
rect 173180 106106 173236 106108
rect 173260 106106 173316 106108
rect 173340 106106 173396 106108
rect 173420 106106 173476 106108
rect 173180 106054 173206 106106
rect 173206 106054 173236 106106
rect 173260 106054 173270 106106
rect 173270 106054 173316 106106
rect 173340 106054 173386 106106
rect 173386 106054 173396 106106
rect 173420 106054 173450 106106
rect 173450 106054 173476 106106
rect 173180 106052 173236 106054
rect 173260 106052 173316 106054
rect 173340 106052 173396 106054
rect 173420 106052 173476 106054
rect 157820 105562 157876 105564
rect 157900 105562 157956 105564
rect 157980 105562 158036 105564
rect 158060 105562 158116 105564
rect 157820 105510 157846 105562
rect 157846 105510 157876 105562
rect 157900 105510 157910 105562
rect 157910 105510 157956 105562
rect 157980 105510 158026 105562
rect 158026 105510 158036 105562
rect 158060 105510 158090 105562
rect 158090 105510 158116 105562
rect 157820 105508 157876 105510
rect 157900 105508 157956 105510
rect 157980 105508 158036 105510
rect 158060 105508 158116 105510
rect 173180 105018 173236 105020
rect 173260 105018 173316 105020
rect 173340 105018 173396 105020
rect 173420 105018 173476 105020
rect 173180 104966 173206 105018
rect 173206 104966 173236 105018
rect 173260 104966 173270 105018
rect 173270 104966 173316 105018
rect 173340 104966 173386 105018
rect 173386 104966 173396 105018
rect 173420 104966 173450 105018
rect 173450 104966 173476 105018
rect 173180 104964 173236 104966
rect 173260 104964 173316 104966
rect 173340 104964 173396 104966
rect 173420 104964 173476 104966
rect 157820 104474 157876 104476
rect 157900 104474 157956 104476
rect 157980 104474 158036 104476
rect 158060 104474 158116 104476
rect 157820 104422 157846 104474
rect 157846 104422 157876 104474
rect 157900 104422 157910 104474
rect 157910 104422 157956 104474
rect 157980 104422 158026 104474
rect 158026 104422 158036 104474
rect 158060 104422 158090 104474
rect 158090 104422 158116 104474
rect 157820 104420 157876 104422
rect 157900 104420 157956 104422
rect 157980 104420 158036 104422
rect 158060 104420 158116 104422
rect 173180 103930 173236 103932
rect 173260 103930 173316 103932
rect 173340 103930 173396 103932
rect 173420 103930 173476 103932
rect 173180 103878 173206 103930
rect 173206 103878 173236 103930
rect 173260 103878 173270 103930
rect 173270 103878 173316 103930
rect 173340 103878 173386 103930
rect 173386 103878 173396 103930
rect 173420 103878 173450 103930
rect 173450 103878 173476 103930
rect 173180 103876 173236 103878
rect 173260 103876 173316 103878
rect 173340 103876 173396 103878
rect 173420 103876 173476 103878
rect 157820 103386 157876 103388
rect 157900 103386 157956 103388
rect 157980 103386 158036 103388
rect 158060 103386 158116 103388
rect 157820 103334 157846 103386
rect 157846 103334 157876 103386
rect 157900 103334 157910 103386
rect 157910 103334 157956 103386
rect 157980 103334 158026 103386
rect 158026 103334 158036 103386
rect 158060 103334 158090 103386
rect 158090 103334 158116 103386
rect 157820 103332 157876 103334
rect 157900 103332 157956 103334
rect 157980 103332 158036 103334
rect 158060 103332 158116 103334
rect 173180 102842 173236 102844
rect 173260 102842 173316 102844
rect 173340 102842 173396 102844
rect 173420 102842 173476 102844
rect 173180 102790 173206 102842
rect 173206 102790 173236 102842
rect 173260 102790 173270 102842
rect 173270 102790 173316 102842
rect 173340 102790 173386 102842
rect 173386 102790 173396 102842
rect 173420 102790 173450 102842
rect 173450 102790 173476 102842
rect 173180 102788 173236 102790
rect 173260 102788 173316 102790
rect 173340 102788 173396 102790
rect 173420 102788 173476 102790
rect 157820 102298 157876 102300
rect 157900 102298 157956 102300
rect 157980 102298 158036 102300
rect 158060 102298 158116 102300
rect 157820 102246 157846 102298
rect 157846 102246 157876 102298
rect 157900 102246 157910 102298
rect 157910 102246 157956 102298
rect 157980 102246 158026 102298
rect 158026 102246 158036 102298
rect 158060 102246 158090 102298
rect 158090 102246 158116 102298
rect 157820 102244 157876 102246
rect 157900 102244 157956 102246
rect 157980 102244 158036 102246
rect 158060 102244 158116 102246
rect 173180 101754 173236 101756
rect 173260 101754 173316 101756
rect 173340 101754 173396 101756
rect 173420 101754 173476 101756
rect 173180 101702 173206 101754
rect 173206 101702 173236 101754
rect 173260 101702 173270 101754
rect 173270 101702 173316 101754
rect 173340 101702 173386 101754
rect 173386 101702 173396 101754
rect 173420 101702 173450 101754
rect 173450 101702 173476 101754
rect 173180 101700 173236 101702
rect 173260 101700 173316 101702
rect 173340 101700 173396 101702
rect 173420 101700 173476 101702
rect 157820 101210 157876 101212
rect 157900 101210 157956 101212
rect 157980 101210 158036 101212
rect 158060 101210 158116 101212
rect 157820 101158 157846 101210
rect 157846 101158 157876 101210
rect 157900 101158 157910 101210
rect 157910 101158 157956 101210
rect 157980 101158 158026 101210
rect 158026 101158 158036 101210
rect 158060 101158 158090 101210
rect 158090 101158 158116 101210
rect 157820 101156 157876 101158
rect 157900 101156 157956 101158
rect 157980 101156 158036 101158
rect 158060 101156 158116 101158
rect 173180 100666 173236 100668
rect 173260 100666 173316 100668
rect 173340 100666 173396 100668
rect 173420 100666 173476 100668
rect 173180 100614 173206 100666
rect 173206 100614 173236 100666
rect 173260 100614 173270 100666
rect 173270 100614 173316 100666
rect 173340 100614 173386 100666
rect 173386 100614 173396 100666
rect 173420 100614 173450 100666
rect 173450 100614 173476 100666
rect 173180 100612 173236 100614
rect 173260 100612 173316 100614
rect 173340 100612 173396 100614
rect 173420 100612 173476 100614
rect 157820 100122 157876 100124
rect 157900 100122 157956 100124
rect 157980 100122 158036 100124
rect 158060 100122 158116 100124
rect 157820 100070 157846 100122
rect 157846 100070 157876 100122
rect 157900 100070 157910 100122
rect 157910 100070 157956 100122
rect 157980 100070 158026 100122
rect 158026 100070 158036 100122
rect 158060 100070 158090 100122
rect 158090 100070 158116 100122
rect 157820 100068 157876 100070
rect 157900 100068 157956 100070
rect 157980 100068 158036 100070
rect 158060 100068 158116 100070
rect 173180 99578 173236 99580
rect 173260 99578 173316 99580
rect 173340 99578 173396 99580
rect 173420 99578 173476 99580
rect 173180 99526 173206 99578
rect 173206 99526 173236 99578
rect 173260 99526 173270 99578
rect 173270 99526 173316 99578
rect 173340 99526 173386 99578
rect 173386 99526 173396 99578
rect 173420 99526 173450 99578
rect 173450 99526 173476 99578
rect 173180 99524 173236 99526
rect 173260 99524 173316 99526
rect 173340 99524 173396 99526
rect 173420 99524 173476 99526
rect 157820 99034 157876 99036
rect 157900 99034 157956 99036
rect 157980 99034 158036 99036
rect 158060 99034 158116 99036
rect 157820 98982 157846 99034
rect 157846 98982 157876 99034
rect 157900 98982 157910 99034
rect 157910 98982 157956 99034
rect 157980 98982 158026 99034
rect 158026 98982 158036 99034
rect 158060 98982 158090 99034
rect 158090 98982 158116 99034
rect 157820 98980 157876 98982
rect 157900 98980 157956 98982
rect 157980 98980 158036 98982
rect 158060 98980 158116 98982
rect 173180 98490 173236 98492
rect 173260 98490 173316 98492
rect 173340 98490 173396 98492
rect 173420 98490 173476 98492
rect 173180 98438 173206 98490
rect 173206 98438 173236 98490
rect 173260 98438 173270 98490
rect 173270 98438 173316 98490
rect 173340 98438 173386 98490
rect 173386 98438 173396 98490
rect 173420 98438 173450 98490
rect 173450 98438 173476 98490
rect 173180 98436 173236 98438
rect 173260 98436 173316 98438
rect 173340 98436 173396 98438
rect 173420 98436 173476 98438
rect 157820 97946 157876 97948
rect 157900 97946 157956 97948
rect 157980 97946 158036 97948
rect 158060 97946 158116 97948
rect 157820 97894 157846 97946
rect 157846 97894 157876 97946
rect 157900 97894 157910 97946
rect 157910 97894 157956 97946
rect 157980 97894 158026 97946
rect 158026 97894 158036 97946
rect 158060 97894 158090 97946
rect 158090 97894 158116 97946
rect 157820 97892 157876 97894
rect 157900 97892 157956 97894
rect 157980 97892 158036 97894
rect 158060 97892 158116 97894
rect 173180 97402 173236 97404
rect 173260 97402 173316 97404
rect 173340 97402 173396 97404
rect 173420 97402 173476 97404
rect 173180 97350 173206 97402
rect 173206 97350 173236 97402
rect 173260 97350 173270 97402
rect 173270 97350 173316 97402
rect 173340 97350 173386 97402
rect 173386 97350 173396 97402
rect 173420 97350 173450 97402
rect 173450 97350 173476 97402
rect 173180 97348 173236 97350
rect 173260 97348 173316 97350
rect 173340 97348 173396 97350
rect 173420 97348 173476 97350
rect 157820 96858 157876 96860
rect 157900 96858 157956 96860
rect 157980 96858 158036 96860
rect 158060 96858 158116 96860
rect 157820 96806 157846 96858
rect 157846 96806 157876 96858
rect 157900 96806 157910 96858
rect 157910 96806 157956 96858
rect 157980 96806 158026 96858
rect 158026 96806 158036 96858
rect 158060 96806 158090 96858
rect 158090 96806 158116 96858
rect 157820 96804 157876 96806
rect 157900 96804 157956 96806
rect 157980 96804 158036 96806
rect 158060 96804 158116 96806
rect 173180 96314 173236 96316
rect 173260 96314 173316 96316
rect 173340 96314 173396 96316
rect 173420 96314 173476 96316
rect 173180 96262 173206 96314
rect 173206 96262 173236 96314
rect 173260 96262 173270 96314
rect 173270 96262 173316 96314
rect 173340 96262 173386 96314
rect 173386 96262 173396 96314
rect 173420 96262 173450 96314
rect 173450 96262 173476 96314
rect 173180 96260 173236 96262
rect 173260 96260 173316 96262
rect 173340 96260 173396 96262
rect 173420 96260 173476 96262
rect 157820 95770 157876 95772
rect 157900 95770 157956 95772
rect 157980 95770 158036 95772
rect 158060 95770 158116 95772
rect 157820 95718 157846 95770
rect 157846 95718 157876 95770
rect 157900 95718 157910 95770
rect 157910 95718 157956 95770
rect 157980 95718 158026 95770
rect 158026 95718 158036 95770
rect 158060 95718 158090 95770
rect 158090 95718 158116 95770
rect 157820 95716 157876 95718
rect 157900 95716 157956 95718
rect 157980 95716 158036 95718
rect 158060 95716 158116 95718
rect 173180 95226 173236 95228
rect 173260 95226 173316 95228
rect 173340 95226 173396 95228
rect 173420 95226 173476 95228
rect 173180 95174 173206 95226
rect 173206 95174 173236 95226
rect 173260 95174 173270 95226
rect 173270 95174 173316 95226
rect 173340 95174 173386 95226
rect 173386 95174 173396 95226
rect 173420 95174 173450 95226
rect 173450 95174 173476 95226
rect 173180 95172 173236 95174
rect 173260 95172 173316 95174
rect 173340 95172 173396 95174
rect 173420 95172 173476 95174
rect 157820 94682 157876 94684
rect 157900 94682 157956 94684
rect 157980 94682 158036 94684
rect 158060 94682 158116 94684
rect 157820 94630 157846 94682
rect 157846 94630 157876 94682
rect 157900 94630 157910 94682
rect 157910 94630 157956 94682
rect 157980 94630 158026 94682
rect 158026 94630 158036 94682
rect 158060 94630 158090 94682
rect 158090 94630 158116 94682
rect 157820 94628 157876 94630
rect 157900 94628 157956 94630
rect 157980 94628 158036 94630
rect 158060 94628 158116 94630
rect 173180 94138 173236 94140
rect 173260 94138 173316 94140
rect 173340 94138 173396 94140
rect 173420 94138 173476 94140
rect 173180 94086 173206 94138
rect 173206 94086 173236 94138
rect 173260 94086 173270 94138
rect 173270 94086 173316 94138
rect 173340 94086 173386 94138
rect 173386 94086 173396 94138
rect 173420 94086 173450 94138
rect 173450 94086 173476 94138
rect 173180 94084 173236 94086
rect 173260 94084 173316 94086
rect 173340 94084 173396 94086
rect 173420 94084 173476 94086
rect 157820 93594 157876 93596
rect 157900 93594 157956 93596
rect 157980 93594 158036 93596
rect 158060 93594 158116 93596
rect 157820 93542 157846 93594
rect 157846 93542 157876 93594
rect 157900 93542 157910 93594
rect 157910 93542 157956 93594
rect 157980 93542 158026 93594
rect 158026 93542 158036 93594
rect 158060 93542 158090 93594
rect 158090 93542 158116 93594
rect 157820 93540 157876 93542
rect 157900 93540 157956 93542
rect 157980 93540 158036 93542
rect 158060 93540 158116 93542
rect 173180 93050 173236 93052
rect 173260 93050 173316 93052
rect 173340 93050 173396 93052
rect 173420 93050 173476 93052
rect 173180 92998 173206 93050
rect 173206 92998 173236 93050
rect 173260 92998 173270 93050
rect 173270 92998 173316 93050
rect 173340 92998 173386 93050
rect 173386 92998 173396 93050
rect 173420 92998 173450 93050
rect 173450 92998 173476 93050
rect 173180 92996 173236 92998
rect 173260 92996 173316 92998
rect 173340 92996 173396 92998
rect 173420 92996 173476 92998
rect 157820 92506 157876 92508
rect 157900 92506 157956 92508
rect 157980 92506 158036 92508
rect 158060 92506 158116 92508
rect 157820 92454 157846 92506
rect 157846 92454 157876 92506
rect 157900 92454 157910 92506
rect 157910 92454 157956 92506
rect 157980 92454 158026 92506
rect 158026 92454 158036 92506
rect 158060 92454 158090 92506
rect 158090 92454 158116 92506
rect 157820 92452 157876 92454
rect 157900 92452 157956 92454
rect 157980 92452 158036 92454
rect 158060 92452 158116 92454
rect 173180 91962 173236 91964
rect 173260 91962 173316 91964
rect 173340 91962 173396 91964
rect 173420 91962 173476 91964
rect 173180 91910 173206 91962
rect 173206 91910 173236 91962
rect 173260 91910 173270 91962
rect 173270 91910 173316 91962
rect 173340 91910 173386 91962
rect 173386 91910 173396 91962
rect 173420 91910 173450 91962
rect 173450 91910 173476 91962
rect 173180 91908 173236 91910
rect 173260 91908 173316 91910
rect 173340 91908 173396 91910
rect 173420 91908 173476 91910
rect 157820 91418 157876 91420
rect 157900 91418 157956 91420
rect 157980 91418 158036 91420
rect 158060 91418 158116 91420
rect 157820 91366 157846 91418
rect 157846 91366 157876 91418
rect 157900 91366 157910 91418
rect 157910 91366 157956 91418
rect 157980 91366 158026 91418
rect 158026 91366 158036 91418
rect 158060 91366 158090 91418
rect 158090 91366 158116 91418
rect 157820 91364 157876 91366
rect 157900 91364 157956 91366
rect 157980 91364 158036 91366
rect 158060 91364 158116 91366
rect 173180 90874 173236 90876
rect 173260 90874 173316 90876
rect 173340 90874 173396 90876
rect 173420 90874 173476 90876
rect 173180 90822 173206 90874
rect 173206 90822 173236 90874
rect 173260 90822 173270 90874
rect 173270 90822 173316 90874
rect 173340 90822 173386 90874
rect 173386 90822 173396 90874
rect 173420 90822 173450 90874
rect 173450 90822 173476 90874
rect 173180 90820 173236 90822
rect 173260 90820 173316 90822
rect 173340 90820 173396 90822
rect 173420 90820 173476 90822
rect 157820 90330 157876 90332
rect 157900 90330 157956 90332
rect 157980 90330 158036 90332
rect 158060 90330 158116 90332
rect 157820 90278 157846 90330
rect 157846 90278 157876 90330
rect 157900 90278 157910 90330
rect 157910 90278 157956 90330
rect 157980 90278 158026 90330
rect 158026 90278 158036 90330
rect 158060 90278 158090 90330
rect 158090 90278 158116 90330
rect 157820 90276 157876 90278
rect 157900 90276 157956 90278
rect 157980 90276 158036 90278
rect 158060 90276 158116 90278
rect 173180 89786 173236 89788
rect 173260 89786 173316 89788
rect 173340 89786 173396 89788
rect 173420 89786 173476 89788
rect 173180 89734 173206 89786
rect 173206 89734 173236 89786
rect 173260 89734 173270 89786
rect 173270 89734 173316 89786
rect 173340 89734 173386 89786
rect 173386 89734 173396 89786
rect 173420 89734 173450 89786
rect 173450 89734 173476 89786
rect 173180 89732 173236 89734
rect 173260 89732 173316 89734
rect 173340 89732 173396 89734
rect 173420 89732 173476 89734
rect 157820 89242 157876 89244
rect 157900 89242 157956 89244
rect 157980 89242 158036 89244
rect 158060 89242 158116 89244
rect 157820 89190 157846 89242
rect 157846 89190 157876 89242
rect 157900 89190 157910 89242
rect 157910 89190 157956 89242
rect 157980 89190 158026 89242
rect 158026 89190 158036 89242
rect 158060 89190 158090 89242
rect 158090 89190 158116 89242
rect 157820 89188 157876 89190
rect 157900 89188 157956 89190
rect 157980 89188 158036 89190
rect 158060 89188 158116 89190
rect 173180 88698 173236 88700
rect 173260 88698 173316 88700
rect 173340 88698 173396 88700
rect 173420 88698 173476 88700
rect 173180 88646 173206 88698
rect 173206 88646 173236 88698
rect 173260 88646 173270 88698
rect 173270 88646 173316 88698
rect 173340 88646 173386 88698
rect 173386 88646 173396 88698
rect 173420 88646 173450 88698
rect 173450 88646 173476 88698
rect 173180 88644 173236 88646
rect 173260 88644 173316 88646
rect 173340 88644 173396 88646
rect 173420 88644 173476 88646
rect 157820 88154 157876 88156
rect 157900 88154 157956 88156
rect 157980 88154 158036 88156
rect 158060 88154 158116 88156
rect 157820 88102 157846 88154
rect 157846 88102 157876 88154
rect 157900 88102 157910 88154
rect 157910 88102 157956 88154
rect 157980 88102 158026 88154
rect 158026 88102 158036 88154
rect 158060 88102 158090 88154
rect 158090 88102 158116 88154
rect 157820 88100 157876 88102
rect 157900 88100 157956 88102
rect 157980 88100 158036 88102
rect 158060 88100 158116 88102
rect 173180 87610 173236 87612
rect 173260 87610 173316 87612
rect 173340 87610 173396 87612
rect 173420 87610 173476 87612
rect 173180 87558 173206 87610
rect 173206 87558 173236 87610
rect 173260 87558 173270 87610
rect 173270 87558 173316 87610
rect 173340 87558 173386 87610
rect 173386 87558 173396 87610
rect 173420 87558 173450 87610
rect 173450 87558 173476 87610
rect 173180 87556 173236 87558
rect 173260 87556 173316 87558
rect 173340 87556 173396 87558
rect 173420 87556 173476 87558
rect 157820 87066 157876 87068
rect 157900 87066 157956 87068
rect 157980 87066 158036 87068
rect 158060 87066 158116 87068
rect 157820 87014 157846 87066
rect 157846 87014 157876 87066
rect 157900 87014 157910 87066
rect 157910 87014 157956 87066
rect 157980 87014 158026 87066
rect 158026 87014 158036 87066
rect 158060 87014 158090 87066
rect 158090 87014 158116 87066
rect 157820 87012 157876 87014
rect 157900 87012 157956 87014
rect 157980 87012 158036 87014
rect 158060 87012 158116 87014
rect 173180 86522 173236 86524
rect 173260 86522 173316 86524
rect 173340 86522 173396 86524
rect 173420 86522 173476 86524
rect 173180 86470 173206 86522
rect 173206 86470 173236 86522
rect 173260 86470 173270 86522
rect 173270 86470 173316 86522
rect 173340 86470 173386 86522
rect 173386 86470 173396 86522
rect 173420 86470 173450 86522
rect 173450 86470 173476 86522
rect 173180 86468 173236 86470
rect 173260 86468 173316 86470
rect 173340 86468 173396 86470
rect 173420 86468 173476 86470
rect 157820 85978 157876 85980
rect 157900 85978 157956 85980
rect 157980 85978 158036 85980
rect 158060 85978 158116 85980
rect 157820 85926 157846 85978
rect 157846 85926 157876 85978
rect 157900 85926 157910 85978
rect 157910 85926 157956 85978
rect 157980 85926 158026 85978
rect 158026 85926 158036 85978
rect 158060 85926 158090 85978
rect 158090 85926 158116 85978
rect 157820 85924 157876 85926
rect 157900 85924 157956 85926
rect 157980 85924 158036 85926
rect 158060 85924 158116 85926
rect 173180 85434 173236 85436
rect 173260 85434 173316 85436
rect 173340 85434 173396 85436
rect 173420 85434 173476 85436
rect 173180 85382 173206 85434
rect 173206 85382 173236 85434
rect 173260 85382 173270 85434
rect 173270 85382 173316 85434
rect 173340 85382 173386 85434
rect 173386 85382 173396 85434
rect 173420 85382 173450 85434
rect 173450 85382 173476 85434
rect 173180 85380 173236 85382
rect 173260 85380 173316 85382
rect 173340 85380 173396 85382
rect 173420 85380 173476 85382
rect 157820 84890 157876 84892
rect 157900 84890 157956 84892
rect 157980 84890 158036 84892
rect 158060 84890 158116 84892
rect 157820 84838 157846 84890
rect 157846 84838 157876 84890
rect 157900 84838 157910 84890
rect 157910 84838 157956 84890
rect 157980 84838 158026 84890
rect 158026 84838 158036 84890
rect 158060 84838 158090 84890
rect 158090 84838 158116 84890
rect 157820 84836 157876 84838
rect 157900 84836 157956 84838
rect 157980 84836 158036 84838
rect 158060 84836 158116 84838
rect 173180 84346 173236 84348
rect 173260 84346 173316 84348
rect 173340 84346 173396 84348
rect 173420 84346 173476 84348
rect 173180 84294 173206 84346
rect 173206 84294 173236 84346
rect 173260 84294 173270 84346
rect 173270 84294 173316 84346
rect 173340 84294 173386 84346
rect 173386 84294 173396 84346
rect 173420 84294 173450 84346
rect 173450 84294 173476 84346
rect 173180 84292 173236 84294
rect 173260 84292 173316 84294
rect 173340 84292 173396 84294
rect 173420 84292 173476 84294
rect 157820 83802 157876 83804
rect 157900 83802 157956 83804
rect 157980 83802 158036 83804
rect 158060 83802 158116 83804
rect 157820 83750 157846 83802
rect 157846 83750 157876 83802
rect 157900 83750 157910 83802
rect 157910 83750 157956 83802
rect 157980 83750 158026 83802
rect 158026 83750 158036 83802
rect 158060 83750 158090 83802
rect 158090 83750 158116 83802
rect 157820 83748 157876 83750
rect 157900 83748 157956 83750
rect 157980 83748 158036 83750
rect 158060 83748 158116 83750
rect 173180 83258 173236 83260
rect 173260 83258 173316 83260
rect 173340 83258 173396 83260
rect 173420 83258 173476 83260
rect 173180 83206 173206 83258
rect 173206 83206 173236 83258
rect 173260 83206 173270 83258
rect 173270 83206 173316 83258
rect 173340 83206 173386 83258
rect 173386 83206 173396 83258
rect 173420 83206 173450 83258
rect 173450 83206 173476 83258
rect 173180 83204 173236 83206
rect 173260 83204 173316 83206
rect 173340 83204 173396 83206
rect 173420 83204 173476 83206
rect 157820 82714 157876 82716
rect 157900 82714 157956 82716
rect 157980 82714 158036 82716
rect 158060 82714 158116 82716
rect 157820 82662 157846 82714
rect 157846 82662 157876 82714
rect 157900 82662 157910 82714
rect 157910 82662 157956 82714
rect 157980 82662 158026 82714
rect 158026 82662 158036 82714
rect 158060 82662 158090 82714
rect 158090 82662 158116 82714
rect 157820 82660 157876 82662
rect 157900 82660 157956 82662
rect 157980 82660 158036 82662
rect 158060 82660 158116 82662
rect 173180 82170 173236 82172
rect 173260 82170 173316 82172
rect 173340 82170 173396 82172
rect 173420 82170 173476 82172
rect 173180 82118 173206 82170
rect 173206 82118 173236 82170
rect 173260 82118 173270 82170
rect 173270 82118 173316 82170
rect 173340 82118 173386 82170
rect 173386 82118 173396 82170
rect 173420 82118 173450 82170
rect 173450 82118 173476 82170
rect 173180 82116 173236 82118
rect 173260 82116 173316 82118
rect 173340 82116 173396 82118
rect 173420 82116 173476 82118
rect 157820 81626 157876 81628
rect 157900 81626 157956 81628
rect 157980 81626 158036 81628
rect 158060 81626 158116 81628
rect 157820 81574 157846 81626
rect 157846 81574 157876 81626
rect 157900 81574 157910 81626
rect 157910 81574 157956 81626
rect 157980 81574 158026 81626
rect 158026 81574 158036 81626
rect 158060 81574 158090 81626
rect 158090 81574 158116 81626
rect 157820 81572 157876 81574
rect 157900 81572 157956 81574
rect 157980 81572 158036 81574
rect 158060 81572 158116 81574
rect 173180 81082 173236 81084
rect 173260 81082 173316 81084
rect 173340 81082 173396 81084
rect 173420 81082 173476 81084
rect 173180 81030 173206 81082
rect 173206 81030 173236 81082
rect 173260 81030 173270 81082
rect 173270 81030 173316 81082
rect 173340 81030 173386 81082
rect 173386 81030 173396 81082
rect 173420 81030 173450 81082
rect 173450 81030 173476 81082
rect 173180 81028 173236 81030
rect 173260 81028 173316 81030
rect 173340 81028 173396 81030
rect 173420 81028 173476 81030
rect 157820 80538 157876 80540
rect 157900 80538 157956 80540
rect 157980 80538 158036 80540
rect 158060 80538 158116 80540
rect 157820 80486 157846 80538
rect 157846 80486 157876 80538
rect 157900 80486 157910 80538
rect 157910 80486 157956 80538
rect 157980 80486 158026 80538
rect 158026 80486 158036 80538
rect 158060 80486 158090 80538
rect 158090 80486 158116 80538
rect 157820 80484 157876 80486
rect 157900 80484 157956 80486
rect 157980 80484 158036 80486
rect 158060 80484 158116 80486
rect 173180 79994 173236 79996
rect 173260 79994 173316 79996
rect 173340 79994 173396 79996
rect 173420 79994 173476 79996
rect 173180 79942 173206 79994
rect 173206 79942 173236 79994
rect 173260 79942 173270 79994
rect 173270 79942 173316 79994
rect 173340 79942 173386 79994
rect 173386 79942 173396 79994
rect 173420 79942 173450 79994
rect 173450 79942 173476 79994
rect 173180 79940 173236 79942
rect 173260 79940 173316 79942
rect 173340 79940 173396 79942
rect 173420 79940 173476 79942
rect 157820 79450 157876 79452
rect 157900 79450 157956 79452
rect 157980 79450 158036 79452
rect 158060 79450 158116 79452
rect 157820 79398 157846 79450
rect 157846 79398 157876 79450
rect 157900 79398 157910 79450
rect 157910 79398 157956 79450
rect 157980 79398 158026 79450
rect 158026 79398 158036 79450
rect 158060 79398 158090 79450
rect 158090 79398 158116 79450
rect 157820 79396 157876 79398
rect 157900 79396 157956 79398
rect 157980 79396 158036 79398
rect 158060 79396 158116 79398
rect 173180 78906 173236 78908
rect 173260 78906 173316 78908
rect 173340 78906 173396 78908
rect 173420 78906 173476 78908
rect 173180 78854 173206 78906
rect 173206 78854 173236 78906
rect 173260 78854 173270 78906
rect 173270 78854 173316 78906
rect 173340 78854 173386 78906
rect 173386 78854 173396 78906
rect 173420 78854 173450 78906
rect 173450 78854 173476 78906
rect 173180 78852 173236 78854
rect 173260 78852 173316 78854
rect 173340 78852 173396 78854
rect 173420 78852 173476 78854
rect 157820 78362 157876 78364
rect 157900 78362 157956 78364
rect 157980 78362 158036 78364
rect 158060 78362 158116 78364
rect 157820 78310 157846 78362
rect 157846 78310 157876 78362
rect 157900 78310 157910 78362
rect 157910 78310 157956 78362
rect 157980 78310 158026 78362
rect 158026 78310 158036 78362
rect 158060 78310 158090 78362
rect 158090 78310 158116 78362
rect 157820 78308 157876 78310
rect 157900 78308 157956 78310
rect 157980 78308 158036 78310
rect 158060 78308 158116 78310
rect 173180 77818 173236 77820
rect 173260 77818 173316 77820
rect 173340 77818 173396 77820
rect 173420 77818 173476 77820
rect 173180 77766 173206 77818
rect 173206 77766 173236 77818
rect 173260 77766 173270 77818
rect 173270 77766 173316 77818
rect 173340 77766 173386 77818
rect 173386 77766 173396 77818
rect 173420 77766 173450 77818
rect 173450 77766 173476 77818
rect 173180 77764 173236 77766
rect 173260 77764 173316 77766
rect 173340 77764 173396 77766
rect 173420 77764 173476 77766
rect 157820 77274 157876 77276
rect 157900 77274 157956 77276
rect 157980 77274 158036 77276
rect 158060 77274 158116 77276
rect 157820 77222 157846 77274
rect 157846 77222 157876 77274
rect 157900 77222 157910 77274
rect 157910 77222 157956 77274
rect 157980 77222 158026 77274
rect 158026 77222 158036 77274
rect 158060 77222 158090 77274
rect 158090 77222 158116 77274
rect 157820 77220 157876 77222
rect 157900 77220 157956 77222
rect 157980 77220 158036 77222
rect 158060 77220 158116 77222
rect 173180 76730 173236 76732
rect 173260 76730 173316 76732
rect 173340 76730 173396 76732
rect 173420 76730 173476 76732
rect 173180 76678 173206 76730
rect 173206 76678 173236 76730
rect 173260 76678 173270 76730
rect 173270 76678 173316 76730
rect 173340 76678 173386 76730
rect 173386 76678 173396 76730
rect 173420 76678 173450 76730
rect 173450 76678 173476 76730
rect 173180 76676 173236 76678
rect 173260 76676 173316 76678
rect 173340 76676 173396 76678
rect 173420 76676 173476 76678
rect 157820 76186 157876 76188
rect 157900 76186 157956 76188
rect 157980 76186 158036 76188
rect 158060 76186 158116 76188
rect 157820 76134 157846 76186
rect 157846 76134 157876 76186
rect 157900 76134 157910 76186
rect 157910 76134 157956 76186
rect 157980 76134 158026 76186
rect 158026 76134 158036 76186
rect 158060 76134 158090 76186
rect 158090 76134 158116 76186
rect 157820 76132 157876 76134
rect 157900 76132 157956 76134
rect 157980 76132 158036 76134
rect 158060 76132 158116 76134
rect 173180 75642 173236 75644
rect 173260 75642 173316 75644
rect 173340 75642 173396 75644
rect 173420 75642 173476 75644
rect 173180 75590 173206 75642
rect 173206 75590 173236 75642
rect 173260 75590 173270 75642
rect 173270 75590 173316 75642
rect 173340 75590 173386 75642
rect 173386 75590 173396 75642
rect 173420 75590 173450 75642
rect 173450 75590 173476 75642
rect 173180 75588 173236 75590
rect 173260 75588 173316 75590
rect 173340 75588 173396 75590
rect 173420 75588 173476 75590
rect 157820 75098 157876 75100
rect 157900 75098 157956 75100
rect 157980 75098 158036 75100
rect 158060 75098 158116 75100
rect 157820 75046 157846 75098
rect 157846 75046 157876 75098
rect 157900 75046 157910 75098
rect 157910 75046 157956 75098
rect 157980 75046 158026 75098
rect 158026 75046 158036 75098
rect 158060 75046 158090 75098
rect 158090 75046 158116 75098
rect 157820 75044 157876 75046
rect 157900 75044 157956 75046
rect 157980 75044 158036 75046
rect 158060 75044 158116 75046
rect 173180 74554 173236 74556
rect 173260 74554 173316 74556
rect 173340 74554 173396 74556
rect 173420 74554 173476 74556
rect 173180 74502 173206 74554
rect 173206 74502 173236 74554
rect 173260 74502 173270 74554
rect 173270 74502 173316 74554
rect 173340 74502 173386 74554
rect 173386 74502 173396 74554
rect 173420 74502 173450 74554
rect 173450 74502 173476 74554
rect 173180 74500 173236 74502
rect 173260 74500 173316 74502
rect 173340 74500 173396 74502
rect 173420 74500 173476 74502
rect 157820 74010 157876 74012
rect 157900 74010 157956 74012
rect 157980 74010 158036 74012
rect 158060 74010 158116 74012
rect 157820 73958 157846 74010
rect 157846 73958 157876 74010
rect 157900 73958 157910 74010
rect 157910 73958 157956 74010
rect 157980 73958 158026 74010
rect 158026 73958 158036 74010
rect 158060 73958 158090 74010
rect 158090 73958 158116 74010
rect 157820 73956 157876 73958
rect 157900 73956 157956 73958
rect 157980 73956 158036 73958
rect 158060 73956 158116 73958
rect 173180 73466 173236 73468
rect 173260 73466 173316 73468
rect 173340 73466 173396 73468
rect 173420 73466 173476 73468
rect 173180 73414 173206 73466
rect 173206 73414 173236 73466
rect 173260 73414 173270 73466
rect 173270 73414 173316 73466
rect 173340 73414 173386 73466
rect 173386 73414 173396 73466
rect 173420 73414 173450 73466
rect 173450 73414 173476 73466
rect 173180 73412 173236 73414
rect 173260 73412 173316 73414
rect 173340 73412 173396 73414
rect 173420 73412 173476 73414
rect 157820 72922 157876 72924
rect 157900 72922 157956 72924
rect 157980 72922 158036 72924
rect 158060 72922 158116 72924
rect 157820 72870 157846 72922
rect 157846 72870 157876 72922
rect 157900 72870 157910 72922
rect 157910 72870 157956 72922
rect 157980 72870 158026 72922
rect 158026 72870 158036 72922
rect 158060 72870 158090 72922
rect 158090 72870 158116 72922
rect 157820 72868 157876 72870
rect 157900 72868 157956 72870
rect 157980 72868 158036 72870
rect 158060 72868 158116 72870
rect 173180 72378 173236 72380
rect 173260 72378 173316 72380
rect 173340 72378 173396 72380
rect 173420 72378 173476 72380
rect 173180 72326 173206 72378
rect 173206 72326 173236 72378
rect 173260 72326 173270 72378
rect 173270 72326 173316 72378
rect 173340 72326 173386 72378
rect 173386 72326 173396 72378
rect 173420 72326 173450 72378
rect 173450 72326 173476 72378
rect 173180 72324 173236 72326
rect 173260 72324 173316 72326
rect 173340 72324 173396 72326
rect 173420 72324 173476 72326
rect 157820 71834 157876 71836
rect 157900 71834 157956 71836
rect 157980 71834 158036 71836
rect 158060 71834 158116 71836
rect 157820 71782 157846 71834
rect 157846 71782 157876 71834
rect 157900 71782 157910 71834
rect 157910 71782 157956 71834
rect 157980 71782 158026 71834
rect 158026 71782 158036 71834
rect 158060 71782 158090 71834
rect 158090 71782 158116 71834
rect 157820 71780 157876 71782
rect 157900 71780 157956 71782
rect 157980 71780 158036 71782
rect 158060 71780 158116 71782
rect 173180 71290 173236 71292
rect 173260 71290 173316 71292
rect 173340 71290 173396 71292
rect 173420 71290 173476 71292
rect 173180 71238 173206 71290
rect 173206 71238 173236 71290
rect 173260 71238 173270 71290
rect 173270 71238 173316 71290
rect 173340 71238 173386 71290
rect 173386 71238 173396 71290
rect 173420 71238 173450 71290
rect 173450 71238 173476 71290
rect 173180 71236 173236 71238
rect 173260 71236 173316 71238
rect 173340 71236 173396 71238
rect 173420 71236 173476 71238
rect 157820 70746 157876 70748
rect 157900 70746 157956 70748
rect 157980 70746 158036 70748
rect 158060 70746 158116 70748
rect 157820 70694 157846 70746
rect 157846 70694 157876 70746
rect 157900 70694 157910 70746
rect 157910 70694 157956 70746
rect 157980 70694 158026 70746
rect 158026 70694 158036 70746
rect 158060 70694 158090 70746
rect 158090 70694 158116 70746
rect 157820 70692 157876 70694
rect 157900 70692 157956 70694
rect 157980 70692 158036 70694
rect 158060 70692 158116 70694
rect 173180 70202 173236 70204
rect 173260 70202 173316 70204
rect 173340 70202 173396 70204
rect 173420 70202 173476 70204
rect 173180 70150 173206 70202
rect 173206 70150 173236 70202
rect 173260 70150 173270 70202
rect 173270 70150 173316 70202
rect 173340 70150 173386 70202
rect 173386 70150 173396 70202
rect 173420 70150 173450 70202
rect 173450 70150 173476 70202
rect 173180 70148 173236 70150
rect 173260 70148 173316 70150
rect 173340 70148 173396 70150
rect 173420 70148 173476 70150
rect 157820 69658 157876 69660
rect 157900 69658 157956 69660
rect 157980 69658 158036 69660
rect 158060 69658 158116 69660
rect 157820 69606 157846 69658
rect 157846 69606 157876 69658
rect 157900 69606 157910 69658
rect 157910 69606 157956 69658
rect 157980 69606 158026 69658
rect 158026 69606 158036 69658
rect 158060 69606 158090 69658
rect 158090 69606 158116 69658
rect 157820 69604 157876 69606
rect 157900 69604 157956 69606
rect 157980 69604 158036 69606
rect 158060 69604 158116 69606
rect 173180 69114 173236 69116
rect 173260 69114 173316 69116
rect 173340 69114 173396 69116
rect 173420 69114 173476 69116
rect 173180 69062 173206 69114
rect 173206 69062 173236 69114
rect 173260 69062 173270 69114
rect 173270 69062 173316 69114
rect 173340 69062 173386 69114
rect 173386 69062 173396 69114
rect 173420 69062 173450 69114
rect 173450 69062 173476 69114
rect 173180 69060 173236 69062
rect 173260 69060 173316 69062
rect 173340 69060 173396 69062
rect 173420 69060 173476 69062
rect 157820 68570 157876 68572
rect 157900 68570 157956 68572
rect 157980 68570 158036 68572
rect 158060 68570 158116 68572
rect 157820 68518 157846 68570
rect 157846 68518 157876 68570
rect 157900 68518 157910 68570
rect 157910 68518 157956 68570
rect 157980 68518 158026 68570
rect 158026 68518 158036 68570
rect 158060 68518 158090 68570
rect 158090 68518 158116 68570
rect 157820 68516 157876 68518
rect 157900 68516 157956 68518
rect 157980 68516 158036 68518
rect 158060 68516 158116 68518
rect 173180 68026 173236 68028
rect 173260 68026 173316 68028
rect 173340 68026 173396 68028
rect 173420 68026 173476 68028
rect 173180 67974 173206 68026
rect 173206 67974 173236 68026
rect 173260 67974 173270 68026
rect 173270 67974 173316 68026
rect 173340 67974 173386 68026
rect 173386 67974 173396 68026
rect 173420 67974 173450 68026
rect 173450 67974 173476 68026
rect 173180 67972 173236 67974
rect 173260 67972 173316 67974
rect 173340 67972 173396 67974
rect 173420 67972 173476 67974
rect 157820 67482 157876 67484
rect 157900 67482 157956 67484
rect 157980 67482 158036 67484
rect 158060 67482 158116 67484
rect 157820 67430 157846 67482
rect 157846 67430 157876 67482
rect 157900 67430 157910 67482
rect 157910 67430 157956 67482
rect 157980 67430 158026 67482
rect 158026 67430 158036 67482
rect 158060 67430 158090 67482
rect 158090 67430 158116 67482
rect 157820 67428 157876 67430
rect 157900 67428 157956 67430
rect 157980 67428 158036 67430
rect 158060 67428 158116 67430
rect 173180 66938 173236 66940
rect 173260 66938 173316 66940
rect 173340 66938 173396 66940
rect 173420 66938 173476 66940
rect 173180 66886 173206 66938
rect 173206 66886 173236 66938
rect 173260 66886 173270 66938
rect 173270 66886 173316 66938
rect 173340 66886 173386 66938
rect 173386 66886 173396 66938
rect 173420 66886 173450 66938
rect 173450 66886 173476 66938
rect 173180 66884 173236 66886
rect 173260 66884 173316 66886
rect 173340 66884 173396 66886
rect 173420 66884 173476 66886
rect 157820 66394 157876 66396
rect 157900 66394 157956 66396
rect 157980 66394 158036 66396
rect 158060 66394 158116 66396
rect 157820 66342 157846 66394
rect 157846 66342 157876 66394
rect 157900 66342 157910 66394
rect 157910 66342 157956 66394
rect 157980 66342 158026 66394
rect 158026 66342 158036 66394
rect 158060 66342 158090 66394
rect 158090 66342 158116 66394
rect 157820 66340 157876 66342
rect 157900 66340 157956 66342
rect 157980 66340 158036 66342
rect 158060 66340 158116 66342
rect 173180 65850 173236 65852
rect 173260 65850 173316 65852
rect 173340 65850 173396 65852
rect 173420 65850 173476 65852
rect 173180 65798 173206 65850
rect 173206 65798 173236 65850
rect 173260 65798 173270 65850
rect 173270 65798 173316 65850
rect 173340 65798 173386 65850
rect 173386 65798 173396 65850
rect 173420 65798 173450 65850
rect 173450 65798 173476 65850
rect 173180 65796 173236 65798
rect 173260 65796 173316 65798
rect 173340 65796 173396 65798
rect 173420 65796 173476 65798
rect 157820 65306 157876 65308
rect 157900 65306 157956 65308
rect 157980 65306 158036 65308
rect 158060 65306 158116 65308
rect 157820 65254 157846 65306
rect 157846 65254 157876 65306
rect 157900 65254 157910 65306
rect 157910 65254 157956 65306
rect 157980 65254 158026 65306
rect 158026 65254 158036 65306
rect 158060 65254 158090 65306
rect 158090 65254 158116 65306
rect 157820 65252 157876 65254
rect 157900 65252 157956 65254
rect 157980 65252 158036 65254
rect 158060 65252 158116 65254
rect 173180 64762 173236 64764
rect 173260 64762 173316 64764
rect 173340 64762 173396 64764
rect 173420 64762 173476 64764
rect 173180 64710 173206 64762
rect 173206 64710 173236 64762
rect 173260 64710 173270 64762
rect 173270 64710 173316 64762
rect 173340 64710 173386 64762
rect 173386 64710 173396 64762
rect 173420 64710 173450 64762
rect 173450 64710 173476 64762
rect 173180 64708 173236 64710
rect 173260 64708 173316 64710
rect 173340 64708 173396 64710
rect 173420 64708 173476 64710
rect 157820 64218 157876 64220
rect 157900 64218 157956 64220
rect 157980 64218 158036 64220
rect 158060 64218 158116 64220
rect 157820 64166 157846 64218
rect 157846 64166 157876 64218
rect 157900 64166 157910 64218
rect 157910 64166 157956 64218
rect 157980 64166 158026 64218
rect 158026 64166 158036 64218
rect 158060 64166 158090 64218
rect 158090 64166 158116 64218
rect 157820 64164 157876 64166
rect 157900 64164 157956 64166
rect 157980 64164 158036 64166
rect 158060 64164 158116 64166
rect 173180 63674 173236 63676
rect 173260 63674 173316 63676
rect 173340 63674 173396 63676
rect 173420 63674 173476 63676
rect 173180 63622 173206 63674
rect 173206 63622 173236 63674
rect 173260 63622 173270 63674
rect 173270 63622 173316 63674
rect 173340 63622 173386 63674
rect 173386 63622 173396 63674
rect 173420 63622 173450 63674
rect 173450 63622 173476 63674
rect 173180 63620 173236 63622
rect 173260 63620 173316 63622
rect 173340 63620 173396 63622
rect 173420 63620 173476 63622
rect 157820 63130 157876 63132
rect 157900 63130 157956 63132
rect 157980 63130 158036 63132
rect 158060 63130 158116 63132
rect 157820 63078 157846 63130
rect 157846 63078 157876 63130
rect 157900 63078 157910 63130
rect 157910 63078 157956 63130
rect 157980 63078 158026 63130
rect 158026 63078 158036 63130
rect 158060 63078 158090 63130
rect 158090 63078 158116 63130
rect 157820 63076 157876 63078
rect 157900 63076 157956 63078
rect 157980 63076 158036 63078
rect 158060 63076 158116 63078
rect 173180 62586 173236 62588
rect 173260 62586 173316 62588
rect 173340 62586 173396 62588
rect 173420 62586 173476 62588
rect 173180 62534 173206 62586
rect 173206 62534 173236 62586
rect 173260 62534 173270 62586
rect 173270 62534 173316 62586
rect 173340 62534 173386 62586
rect 173386 62534 173396 62586
rect 173420 62534 173450 62586
rect 173450 62534 173476 62586
rect 173180 62532 173236 62534
rect 173260 62532 173316 62534
rect 173340 62532 173396 62534
rect 173420 62532 173476 62534
rect 157820 62042 157876 62044
rect 157900 62042 157956 62044
rect 157980 62042 158036 62044
rect 158060 62042 158116 62044
rect 157820 61990 157846 62042
rect 157846 61990 157876 62042
rect 157900 61990 157910 62042
rect 157910 61990 157956 62042
rect 157980 61990 158026 62042
rect 158026 61990 158036 62042
rect 158060 61990 158090 62042
rect 158090 61990 158116 62042
rect 157820 61988 157876 61990
rect 157900 61988 157956 61990
rect 157980 61988 158036 61990
rect 158060 61988 158116 61990
rect 173180 61498 173236 61500
rect 173260 61498 173316 61500
rect 173340 61498 173396 61500
rect 173420 61498 173476 61500
rect 173180 61446 173206 61498
rect 173206 61446 173236 61498
rect 173260 61446 173270 61498
rect 173270 61446 173316 61498
rect 173340 61446 173386 61498
rect 173386 61446 173396 61498
rect 173420 61446 173450 61498
rect 173450 61446 173476 61498
rect 173180 61444 173236 61446
rect 173260 61444 173316 61446
rect 173340 61444 173396 61446
rect 173420 61444 173476 61446
rect 157820 60954 157876 60956
rect 157900 60954 157956 60956
rect 157980 60954 158036 60956
rect 158060 60954 158116 60956
rect 157820 60902 157846 60954
rect 157846 60902 157876 60954
rect 157900 60902 157910 60954
rect 157910 60902 157956 60954
rect 157980 60902 158026 60954
rect 158026 60902 158036 60954
rect 158060 60902 158090 60954
rect 158090 60902 158116 60954
rect 157820 60900 157876 60902
rect 157900 60900 157956 60902
rect 157980 60900 158036 60902
rect 158060 60900 158116 60902
rect 173180 60410 173236 60412
rect 173260 60410 173316 60412
rect 173340 60410 173396 60412
rect 173420 60410 173476 60412
rect 173180 60358 173206 60410
rect 173206 60358 173236 60410
rect 173260 60358 173270 60410
rect 173270 60358 173316 60410
rect 173340 60358 173386 60410
rect 173386 60358 173396 60410
rect 173420 60358 173450 60410
rect 173450 60358 173476 60410
rect 173180 60356 173236 60358
rect 173260 60356 173316 60358
rect 173340 60356 173396 60358
rect 173420 60356 173476 60358
rect 157820 59866 157876 59868
rect 157900 59866 157956 59868
rect 157980 59866 158036 59868
rect 158060 59866 158116 59868
rect 157820 59814 157846 59866
rect 157846 59814 157876 59866
rect 157900 59814 157910 59866
rect 157910 59814 157956 59866
rect 157980 59814 158026 59866
rect 158026 59814 158036 59866
rect 158060 59814 158090 59866
rect 158090 59814 158116 59866
rect 157820 59812 157876 59814
rect 157900 59812 157956 59814
rect 157980 59812 158036 59814
rect 158060 59812 158116 59814
rect 178130 60036 178186 60072
rect 178130 60016 178132 60036
rect 178132 60016 178184 60036
rect 178184 60016 178186 60036
rect 173180 59322 173236 59324
rect 173260 59322 173316 59324
rect 173340 59322 173396 59324
rect 173420 59322 173476 59324
rect 173180 59270 173206 59322
rect 173206 59270 173236 59322
rect 173260 59270 173270 59322
rect 173270 59270 173316 59322
rect 173340 59270 173386 59322
rect 173386 59270 173396 59322
rect 173420 59270 173450 59322
rect 173450 59270 173476 59322
rect 173180 59268 173236 59270
rect 173260 59268 173316 59270
rect 173340 59268 173396 59270
rect 173420 59268 173476 59270
rect 157820 58778 157876 58780
rect 157900 58778 157956 58780
rect 157980 58778 158036 58780
rect 158060 58778 158116 58780
rect 157820 58726 157846 58778
rect 157846 58726 157876 58778
rect 157900 58726 157910 58778
rect 157910 58726 157956 58778
rect 157980 58726 158026 58778
rect 158026 58726 158036 58778
rect 158060 58726 158090 58778
rect 158090 58726 158116 58778
rect 157820 58724 157876 58726
rect 157900 58724 157956 58726
rect 157980 58724 158036 58726
rect 158060 58724 158116 58726
rect 173180 58234 173236 58236
rect 173260 58234 173316 58236
rect 173340 58234 173396 58236
rect 173420 58234 173476 58236
rect 173180 58182 173206 58234
rect 173206 58182 173236 58234
rect 173260 58182 173270 58234
rect 173270 58182 173316 58234
rect 173340 58182 173386 58234
rect 173386 58182 173396 58234
rect 173420 58182 173450 58234
rect 173450 58182 173476 58234
rect 173180 58180 173236 58182
rect 173260 58180 173316 58182
rect 173340 58180 173396 58182
rect 173420 58180 173476 58182
rect 157820 57690 157876 57692
rect 157900 57690 157956 57692
rect 157980 57690 158036 57692
rect 158060 57690 158116 57692
rect 157820 57638 157846 57690
rect 157846 57638 157876 57690
rect 157900 57638 157910 57690
rect 157910 57638 157956 57690
rect 157980 57638 158026 57690
rect 158026 57638 158036 57690
rect 158060 57638 158090 57690
rect 158090 57638 158116 57690
rect 157820 57636 157876 57638
rect 157900 57636 157956 57638
rect 157980 57636 158036 57638
rect 158060 57636 158116 57638
rect 173180 57146 173236 57148
rect 173260 57146 173316 57148
rect 173340 57146 173396 57148
rect 173420 57146 173476 57148
rect 173180 57094 173206 57146
rect 173206 57094 173236 57146
rect 173260 57094 173270 57146
rect 173270 57094 173316 57146
rect 173340 57094 173386 57146
rect 173386 57094 173396 57146
rect 173420 57094 173450 57146
rect 173450 57094 173476 57146
rect 173180 57092 173236 57094
rect 173260 57092 173316 57094
rect 173340 57092 173396 57094
rect 173420 57092 173476 57094
rect 157820 56602 157876 56604
rect 157900 56602 157956 56604
rect 157980 56602 158036 56604
rect 158060 56602 158116 56604
rect 157820 56550 157846 56602
rect 157846 56550 157876 56602
rect 157900 56550 157910 56602
rect 157910 56550 157956 56602
rect 157980 56550 158026 56602
rect 158026 56550 158036 56602
rect 158060 56550 158090 56602
rect 158090 56550 158116 56602
rect 157820 56548 157876 56550
rect 157900 56548 157956 56550
rect 157980 56548 158036 56550
rect 158060 56548 158116 56550
rect 173180 56058 173236 56060
rect 173260 56058 173316 56060
rect 173340 56058 173396 56060
rect 173420 56058 173476 56060
rect 173180 56006 173206 56058
rect 173206 56006 173236 56058
rect 173260 56006 173270 56058
rect 173270 56006 173316 56058
rect 173340 56006 173386 56058
rect 173386 56006 173396 56058
rect 173420 56006 173450 56058
rect 173450 56006 173476 56058
rect 173180 56004 173236 56006
rect 173260 56004 173316 56006
rect 173340 56004 173396 56006
rect 173420 56004 173476 56006
rect 157820 55514 157876 55516
rect 157900 55514 157956 55516
rect 157980 55514 158036 55516
rect 158060 55514 158116 55516
rect 157820 55462 157846 55514
rect 157846 55462 157876 55514
rect 157900 55462 157910 55514
rect 157910 55462 157956 55514
rect 157980 55462 158026 55514
rect 158026 55462 158036 55514
rect 158060 55462 158090 55514
rect 158090 55462 158116 55514
rect 157820 55460 157876 55462
rect 157900 55460 157956 55462
rect 157980 55460 158036 55462
rect 158060 55460 158116 55462
rect 173180 54970 173236 54972
rect 173260 54970 173316 54972
rect 173340 54970 173396 54972
rect 173420 54970 173476 54972
rect 173180 54918 173206 54970
rect 173206 54918 173236 54970
rect 173260 54918 173270 54970
rect 173270 54918 173316 54970
rect 173340 54918 173386 54970
rect 173386 54918 173396 54970
rect 173420 54918 173450 54970
rect 173450 54918 173476 54970
rect 173180 54916 173236 54918
rect 173260 54916 173316 54918
rect 173340 54916 173396 54918
rect 173420 54916 173476 54918
rect 157820 54426 157876 54428
rect 157900 54426 157956 54428
rect 157980 54426 158036 54428
rect 158060 54426 158116 54428
rect 157820 54374 157846 54426
rect 157846 54374 157876 54426
rect 157900 54374 157910 54426
rect 157910 54374 157956 54426
rect 157980 54374 158026 54426
rect 158026 54374 158036 54426
rect 158060 54374 158090 54426
rect 158090 54374 158116 54426
rect 157820 54372 157876 54374
rect 157900 54372 157956 54374
rect 157980 54372 158036 54374
rect 158060 54372 158116 54374
rect 173180 53882 173236 53884
rect 173260 53882 173316 53884
rect 173340 53882 173396 53884
rect 173420 53882 173476 53884
rect 173180 53830 173206 53882
rect 173206 53830 173236 53882
rect 173260 53830 173270 53882
rect 173270 53830 173316 53882
rect 173340 53830 173386 53882
rect 173386 53830 173396 53882
rect 173420 53830 173450 53882
rect 173450 53830 173476 53882
rect 173180 53828 173236 53830
rect 173260 53828 173316 53830
rect 173340 53828 173396 53830
rect 173420 53828 173476 53830
rect 157820 53338 157876 53340
rect 157900 53338 157956 53340
rect 157980 53338 158036 53340
rect 158060 53338 158116 53340
rect 157820 53286 157846 53338
rect 157846 53286 157876 53338
rect 157900 53286 157910 53338
rect 157910 53286 157956 53338
rect 157980 53286 158026 53338
rect 158026 53286 158036 53338
rect 158060 53286 158090 53338
rect 158090 53286 158116 53338
rect 157820 53284 157876 53286
rect 157900 53284 157956 53286
rect 157980 53284 158036 53286
rect 158060 53284 158116 53286
rect 173180 52794 173236 52796
rect 173260 52794 173316 52796
rect 173340 52794 173396 52796
rect 173420 52794 173476 52796
rect 173180 52742 173206 52794
rect 173206 52742 173236 52794
rect 173260 52742 173270 52794
rect 173270 52742 173316 52794
rect 173340 52742 173386 52794
rect 173386 52742 173396 52794
rect 173420 52742 173450 52794
rect 173450 52742 173476 52794
rect 173180 52740 173236 52742
rect 173260 52740 173316 52742
rect 173340 52740 173396 52742
rect 173420 52740 173476 52742
rect 157820 52250 157876 52252
rect 157900 52250 157956 52252
rect 157980 52250 158036 52252
rect 158060 52250 158116 52252
rect 157820 52198 157846 52250
rect 157846 52198 157876 52250
rect 157900 52198 157910 52250
rect 157910 52198 157956 52250
rect 157980 52198 158026 52250
rect 158026 52198 158036 52250
rect 158060 52198 158090 52250
rect 158090 52198 158116 52250
rect 157820 52196 157876 52198
rect 157900 52196 157956 52198
rect 157980 52196 158036 52198
rect 158060 52196 158116 52198
rect 173180 51706 173236 51708
rect 173260 51706 173316 51708
rect 173340 51706 173396 51708
rect 173420 51706 173476 51708
rect 173180 51654 173206 51706
rect 173206 51654 173236 51706
rect 173260 51654 173270 51706
rect 173270 51654 173316 51706
rect 173340 51654 173386 51706
rect 173386 51654 173396 51706
rect 173420 51654 173450 51706
rect 173450 51654 173476 51706
rect 173180 51652 173236 51654
rect 173260 51652 173316 51654
rect 173340 51652 173396 51654
rect 173420 51652 173476 51654
rect 157820 51162 157876 51164
rect 157900 51162 157956 51164
rect 157980 51162 158036 51164
rect 158060 51162 158116 51164
rect 157820 51110 157846 51162
rect 157846 51110 157876 51162
rect 157900 51110 157910 51162
rect 157910 51110 157956 51162
rect 157980 51110 158026 51162
rect 158026 51110 158036 51162
rect 158060 51110 158090 51162
rect 158090 51110 158116 51162
rect 157820 51108 157876 51110
rect 157900 51108 157956 51110
rect 157980 51108 158036 51110
rect 158060 51108 158116 51110
rect 173180 50618 173236 50620
rect 173260 50618 173316 50620
rect 173340 50618 173396 50620
rect 173420 50618 173476 50620
rect 173180 50566 173206 50618
rect 173206 50566 173236 50618
rect 173260 50566 173270 50618
rect 173270 50566 173316 50618
rect 173340 50566 173386 50618
rect 173386 50566 173396 50618
rect 173420 50566 173450 50618
rect 173450 50566 173476 50618
rect 173180 50564 173236 50566
rect 173260 50564 173316 50566
rect 173340 50564 173396 50566
rect 173420 50564 173476 50566
rect 157820 50074 157876 50076
rect 157900 50074 157956 50076
rect 157980 50074 158036 50076
rect 158060 50074 158116 50076
rect 157820 50022 157846 50074
rect 157846 50022 157876 50074
rect 157900 50022 157910 50074
rect 157910 50022 157956 50074
rect 157980 50022 158026 50074
rect 158026 50022 158036 50074
rect 158060 50022 158090 50074
rect 158090 50022 158116 50074
rect 157820 50020 157876 50022
rect 157900 50020 157956 50022
rect 157980 50020 158036 50022
rect 158060 50020 158116 50022
rect 173180 49530 173236 49532
rect 173260 49530 173316 49532
rect 173340 49530 173396 49532
rect 173420 49530 173476 49532
rect 173180 49478 173206 49530
rect 173206 49478 173236 49530
rect 173260 49478 173270 49530
rect 173270 49478 173316 49530
rect 173340 49478 173386 49530
rect 173386 49478 173396 49530
rect 173420 49478 173450 49530
rect 173450 49478 173476 49530
rect 173180 49476 173236 49478
rect 173260 49476 173316 49478
rect 173340 49476 173396 49478
rect 173420 49476 173476 49478
rect 157820 48986 157876 48988
rect 157900 48986 157956 48988
rect 157980 48986 158036 48988
rect 158060 48986 158116 48988
rect 157820 48934 157846 48986
rect 157846 48934 157876 48986
rect 157900 48934 157910 48986
rect 157910 48934 157956 48986
rect 157980 48934 158026 48986
rect 158026 48934 158036 48986
rect 158060 48934 158090 48986
rect 158090 48934 158116 48986
rect 157820 48932 157876 48934
rect 157900 48932 157956 48934
rect 157980 48932 158036 48934
rect 158060 48932 158116 48934
rect 173180 48442 173236 48444
rect 173260 48442 173316 48444
rect 173340 48442 173396 48444
rect 173420 48442 173476 48444
rect 173180 48390 173206 48442
rect 173206 48390 173236 48442
rect 173260 48390 173270 48442
rect 173270 48390 173316 48442
rect 173340 48390 173386 48442
rect 173386 48390 173396 48442
rect 173420 48390 173450 48442
rect 173450 48390 173476 48442
rect 173180 48388 173236 48390
rect 173260 48388 173316 48390
rect 173340 48388 173396 48390
rect 173420 48388 173476 48390
rect 157820 47898 157876 47900
rect 157900 47898 157956 47900
rect 157980 47898 158036 47900
rect 158060 47898 158116 47900
rect 157820 47846 157846 47898
rect 157846 47846 157876 47898
rect 157900 47846 157910 47898
rect 157910 47846 157956 47898
rect 157980 47846 158026 47898
rect 158026 47846 158036 47898
rect 158060 47846 158090 47898
rect 158090 47846 158116 47898
rect 157820 47844 157876 47846
rect 157900 47844 157956 47846
rect 157980 47844 158036 47846
rect 158060 47844 158116 47846
rect 173180 47354 173236 47356
rect 173260 47354 173316 47356
rect 173340 47354 173396 47356
rect 173420 47354 173476 47356
rect 173180 47302 173206 47354
rect 173206 47302 173236 47354
rect 173260 47302 173270 47354
rect 173270 47302 173316 47354
rect 173340 47302 173386 47354
rect 173386 47302 173396 47354
rect 173420 47302 173450 47354
rect 173450 47302 173476 47354
rect 173180 47300 173236 47302
rect 173260 47300 173316 47302
rect 173340 47300 173396 47302
rect 173420 47300 173476 47302
rect 157820 46810 157876 46812
rect 157900 46810 157956 46812
rect 157980 46810 158036 46812
rect 158060 46810 158116 46812
rect 157820 46758 157846 46810
rect 157846 46758 157876 46810
rect 157900 46758 157910 46810
rect 157910 46758 157956 46810
rect 157980 46758 158026 46810
rect 158026 46758 158036 46810
rect 158060 46758 158090 46810
rect 158090 46758 158116 46810
rect 157820 46756 157876 46758
rect 157900 46756 157956 46758
rect 157980 46756 158036 46758
rect 158060 46756 158116 46758
rect 173180 46266 173236 46268
rect 173260 46266 173316 46268
rect 173340 46266 173396 46268
rect 173420 46266 173476 46268
rect 173180 46214 173206 46266
rect 173206 46214 173236 46266
rect 173260 46214 173270 46266
rect 173270 46214 173316 46266
rect 173340 46214 173386 46266
rect 173386 46214 173396 46266
rect 173420 46214 173450 46266
rect 173450 46214 173476 46266
rect 173180 46212 173236 46214
rect 173260 46212 173316 46214
rect 173340 46212 173396 46214
rect 173420 46212 173476 46214
rect 157820 45722 157876 45724
rect 157900 45722 157956 45724
rect 157980 45722 158036 45724
rect 158060 45722 158116 45724
rect 157820 45670 157846 45722
rect 157846 45670 157876 45722
rect 157900 45670 157910 45722
rect 157910 45670 157956 45722
rect 157980 45670 158026 45722
rect 158026 45670 158036 45722
rect 158060 45670 158090 45722
rect 158090 45670 158116 45722
rect 157820 45668 157876 45670
rect 157900 45668 157956 45670
rect 157980 45668 158036 45670
rect 158060 45668 158116 45670
rect 173180 45178 173236 45180
rect 173260 45178 173316 45180
rect 173340 45178 173396 45180
rect 173420 45178 173476 45180
rect 173180 45126 173206 45178
rect 173206 45126 173236 45178
rect 173260 45126 173270 45178
rect 173270 45126 173316 45178
rect 173340 45126 173386 45178
rect 173386 45126 173396 45178
rect 173420 45126 173450 45178
rect 173450 45126 173476 45178
rect 173180 45124 173236 45126
rect 173260 45124 173316 45126
rect 173340 45124 173396 45126
rect 173420 45124 173476 45126
rect 157820 44634 157876 44636
rect 157900 44634 157956 44636
rect 157980 44634 158036 44636
rect 158060 44634 158116 44636
rect 157820 44582 157846 44634
rect 157846 44582 157876 44634
rect 157900 44582 157910 44634
rect 157910 44582 157956 44634
rect 157980 44582 158026 44634
rect 158026 44582 158036 44634
rect 158060 44582 158090 44634
rect 158090 44582 158116 44634
rect 157820 44580 157876 44582
rect 157900 44580 157956 44582
rect 157980 44580 158036 44582
rect 158060 44580 158116 44582
rect 173180 44090 173236 44092
rect 173260 44090 173316 44092
rect 173340 44090 173396 44092
rect 173420 44090 173476 44092
rect 173180 44038 173206 44090
rect 173206 44038 173236 44090
rect 173260 44038 173270 44090
rect 173270 44038 173316 44090
rect 173340 44038 173386 44090
rect 173386 44038 173396 44090
rect 173420 44038 173450 44090
rect 173450 44038 173476 44090
rect 173180 44036 173236 44038
rect 173260 44036 173316 44038
rect 173340 44036 173396 44038
rect 173420 44036 173476 44038
rect 157820 43546 157876 43548
rect 157900 43546 157956 43548
rect 157980 43546 158036 43548
rect 158060 43546 158116 43548
rect 157820 43494 157846 43546
rect 157846 43494 157876 43546
rect 157900 43494 157910 43546
rect 157910 43494 157956 43546
rect 157980 43494 158026 43546
rect 158026 43494 158036 43546
rect 158060 43494 158090 43546
rect 158090 43494 158116 43546
rect 157820 43492 157876 43494
rect 157900 43492 157956 43494
rect 157980 43492 158036 43494
rect 158060 43492 158116 43494
rect 173180 43002 173236 43004
rect 173260 43002 173316 43004
rect 173340 43002 173396 43004
rect 173420 43002 173476 43004
rect 173180 42950 173206 43002
rect 173206 42950 173236 43002
rect 173260 42950 173270 43002
rect 173270 42950 173316 43002
rect 173340 42950 173386 43002
rect 173386 42950 173396 43002
rect 173420 42950 173450 43002
rect 173450 42950 173476 43002
rect 173180 42948 173236 42950
rect 173260 42948 173316 42950
rect 173340 42948 173396 42950
rect 173420 42948 173476 42950
rect 157820 42458 157876 42460
rect 157900 42458 157956 42460
rect 157980 42458 158036 42460
rect 158060 42458 158116 42460
rect 157820 42406 157846 42458
rect 157846 42406 157876 42458
rect 157900 42406 157910 42458
rect 157910 42406 157956 42458
rect 157980 42406 158026 42458
rect 158026 42406 158036 42458
rect 158060 42406 158090 42458
rect 158090 42406 158116 42458
rect 157820 42404 157876 42406
rect 157900 42404 157956 42406
rect 157980 42404 158036 42406
rect 158060 42404 158116 42406
rect 173180 41914 173236 41916
rect 173260 41914 173316 41916
rect 173340 41914 173396 41916
rect 173420 41914 173476 41916
rect 173180 41862 173206 41914
rect 173206 41862 173236 41914
rect 173260 41862 173270 41914
rect 173270 41862 173316 41914
rect 173340 41862 173386 41914
rect 173386 41862 173396 41914
rect 173420 41862 173450 41914
rect 173450 41862 173476 41914
rect 173180 41860 173236 41862
rect 173260 41860 173316 41862
rect 173340 41860 173396 41862
rect 173420 41860 173476 41862
rect 157820 41370 157876 41372
rect 157900 41370 157956 41372
rect 157980 41370 158036 41372
rect 158060 41370 158116 41372
rect 157820 41318 157846 41370
rect 157846 41318 157876 41370
rect 157900 41318 157910 41370
rect 157910 41318 157956 41370
rect 157980 41318 158026 41370
rect 158026 41318 158036 41370
rect 158060 41318 158090 41370
rect 158090 41318 158116 41370
rect 157820 41316 157876 41318
rect 157900 41316 157956 41318
rect 157980 41316 158036 41318
rect 158060 41316 158116 41318
rect 173180 40826 173236 40828
rect 173260 40826 173316 40828
rect 173340 40826 173396 40828
rect 173420 40826 173476 40828
rect 173180 40774 173206 40826
rect 173206 40774 173236 40826
rect 173260 40774 173270 40826
rect 173270 40774 173316 40826
rect 173340 40774 173386 40826
rect 173386 40774 173396 40826
rect 173420 40774 173450 40826
rect 173450 40774 173476 40826
rect 173180 40772 173236 40774
rect 173260 40772 173316 40774
rect 173340 40772 173396 40774
rect 173420 40772 173476 40774
rect 157820 40282 157876 40284
rect 157900 40282 157956 40284
rect 157980 40282 158036 40284
rect 158060 40282 158116 40284
rect 157820 40230 157846 40282
rect 157846 40230 157876 40282
rect 157900 40230 157910 40282
rect 157910 40230 157956 40282
rect 157980 40230 158026 40282
rect 158026 40230 158036 40282
rect 158060 40230 158090 40282
rect 158090 40230 158116 40282
rect 157820 40228 157876 40230
rect 157900 40228 157956 40230
rect 157980 40228 158036 40230
rect 158060 40228 158116 40230
rect 173180 39738 173236 39740
rect 173260 39738 173316 39740
rect 173340 39738 173396 39740
rect 173420 39738 173476 39740
rect 173180 39686 173206 39738
rect 173206 39686 173236 39738
rect 173260 39686 173270 39738
rect 173270 39686 173316 39738
rect 173340 39686 173386 39738
rect 173386 39686 173396 39738
rect 173420 39686 173450 39738
rect 173450 39686 173476 39738
rect 173180 39684 173236 39686
rect 173260 39684 173316 39686
rect 173340 39684 173396 39686
rect 173420 39684 173476 39686
rect 157820 39194 157876 39196
rect 157900 39194 157956 39196
rect 157980 39194 158036 39196
rect 158060 39194 158116 39196
rect 157820 39142 157846 39194
rect 157846 39142 157876 39194
rect 157900 39142 157910 39194
rect 157910 39142 157956 39194
rect 157980 39142 158026 39194
rect 158026 39142 158036 39194
rect 158060 39142 158090 39194
rect 158090 39142 158116 39194
rect 157820 39140 157876 39142
rect 157900 39140 157956 39142
rect 157980 39140 158036 39142
rect 158060 39140 158116 39142
rect 173180 38650 173236 38652
rect 173260 38650 173316 38652
rect 173340 38650 173396 38652
rect 173420 38650 173476 38652
rect 173180 38598 173206 38650
rect 173206 38598 173236 38650
rect 173260 38598 173270 38650
rect 173270 38598 173316 38650
rect 173340 38598 173386 38650
rect 173386 38598 173396 38650
rect 173420 38598 173450 38650
rect 173450 38598 173476 38650
rect 173180 38596 173236 38598
rect 173260 38596 173316 38598
rect 173340 38596 173396 38598
rect 173420 38596 173476 38598
rect 157820 38106 157876 38108
rect 157900 38106 157956 38108
rect 157980 38106 158036 38108
rect 158060 38106 158116 38108
rect 157820 38054 157846 38106
rect 157846 38054 157876 38106
rect 157900 38054 157910 38106
rect 157910 38054 157956 38106
rect 157980 38054 158026 38106
rect 158026 38054 158036 38106
rect 158060 38054 158090 38106
rect 158090 38054 158116 38106
rect 157820 38052 157876 38054
rect 157900 38052 157956 38054
rect 157980 38052 158036 38054
rect 158060 38052 158116 38054
rect 173180 37562 173236 37564
rect 173260 37562 173316 37564
rect 173340 37562 173396 37564
rect 173420 37562 173476 37564
rect 173180 37510 173206 37562
rect 173206 37510 173236 37562
rect 173260 37510 173270 37562
rect 173270 37510 173316 37562
rect 173340 37510 173386 37562
rect 173386 37510 173396 37562
rect 173420 37510 173450 37562
rect 173450 37510 173476 37562
rect 173180 37508 173236 37510
rect 173260 37508 173316 37510
rect 173340 37508 173396 37510
rect 173420 37508 173476 37510
rect 157820 37018 157876 37020
rect 157900 37018 157956 37020
rect 157980 37018 158036 37020
rect 158060 37018 158116 37020
rect 157820 36966 157846 37018
rect 157846 36966 157876 37018
rect 157900 36966 157910 37018
rect 157910 36966 157956 37018
rect 157980 36966 158026 37018
rect 158026 36966 158036 37018
rect 158060 36966 158090 37018
rect 158090 36966 158116 37018
rect 157820 36964 157876 36966
rect 157900 36964 157956 36966
rect 157980 36964 158036 36966
rect 158060 36964 158116 36966
rect 173180 36474 173236 36476
rect 173260 36474 173316 36476
rect 173340 36474 173396 36476
rect 173420 36474 173476 36476
rect 173180 36422 173206 36474
rect 173206 36422 173236 36474
rect 173260 36422 173270 36474
rect 173270 36422 173316 36474
rect 173340 36422 173386 36474
rect 173386 36422 173396 36474
rect 173420 36422 173450 36474
rect 173450 36422 173476 36474
rect 173180 36420 173236 36422
rect 173260 36420 173316 36422
rect 173340 36420 173396 36422
rect 173420 36420 173476 36422
rect 157820 35930 157876 35932
rect 157900 35930 157956 35932
rect 157980 35930 158036 35932
rect 158060 35930 158116 35932
rect 157820 35878 157846 35930
rect 157846 35878 157876 35930
rect 157900 35878 157910 35930
rect 157910 35878 157956 35930
rect 157980 35878 158026 35930
rect 158026 35878 158036 35930
rect 158060 35878 158090 35930
rect 158090 35878 158116 35930
rect 157820 35876 157876 35878
rect 157900 35876 157956 35878
rect 157980 35876 158036 35878
rect 158060 35876 158116 35878
rect 173180 35386 173236 35388
rect 173260 35386 173316 35388
rect 173340 35386 173396 35388
rect 173420 35386 173476 35388
rect 173180 35334 173206 35386
rect 173206 35334 173236 35386
rect 173260 35334 173270 35386
rect 173270 35334 173316 35386
rect 173340 35334 173386 35386
rect 173386 35334 173396 35386
rect 173420 35334 173450 35386
rect 173450 35334 173476 35386
rect 173180 35332 173236 35334
rect 173260 35332 173316 35334
rect 173340 35332 173396 35334
rect 173420 35332 173476 35334
rect 157820 34842 157876 34844
rect 157900 34842 157956 34844
rect 157980 34842 158036 34844
rect 158060 34842 158116 34844
rect 157820 34790 157846 34842
rect 157846 34790 157876 34842
rect 157900 34790 157910 34842
rect 157910 34790 157956 34842
rect 157980 34790 158026 34842
rect 158026 34790 158036 34842
rect 158060 34790 158090 34842
rect 158090 34790 158116 34842
rect 157820 34788 157876 34790
rect 157900 34788 157956 34790
rect 157980 34788 158036 34790
rect 158060 34788 158116 34790
rect 173180 34298 173236 34300
rect 173260 34298 173316 34300
rect 173340 34298 173396 34300
rect 173420 34298 173476 34300
rect 173180 34246 173206 34298
rect 173206 34246 173236 34298
rect 173260 34246 173270 34298
rect 173270 34246 173316 34298
rect 173340 34246 173386 34298
rect 173386 34246 173396 34298
rect 173420 34246 173450 34298
rect 173450 34246 173476 34298
rect 173180 34244 173236 34246
rect 173260 34244 173316 34246
rect 173340 34244 173396 34246
rect 173420 34244 173476 34246
rect 157820 33754 157876 33756
rect 157900 33754 157956 33756
rect 157980 33754 158036 33756
rect 158060 33754 158116 33756
rect 157820 33702 157846 33754
rect 157846 33702 157876 33754
rect 157900 33702 157910 33754
rect 157910 33702 157956 33754
rect 157980 33702 158026 33754
rect 158026 33702 158036 33754
rect 158060 33702 158090 33754
rect 158090 33702 158116 33754
rect 157820 33700 157876 33702
rect 157900 33700 157956 33702
rect 157980 33700 158036 33702
rect 158060 33700 158116 33702
rect 173180 33210 173236 33212
rect 173260 33210 173316 33212
rect 173340 33210 173396 33212
rect 173420 33210 173476 33212
rect 173180 33158 173206 33210
rect 173206 33158 173236 33210
rect 173260 33158 173270 33210
rect 173270 33158 173316 33210
rect 173340 33158 173386 33210
rect 173386 33158 173396 33210
rect 173420 33158 173450 33210
rect 173450 33158 173476 33210
rect 173180 33156 173236 33158
rect 173260 33156 173316 33158
rect 173340 33156 173396 33158
rect 173420 33156 173476 33158
rect 157820 32666 157876 32668
rect 157900 32666 157956 32668
rect 157980 32666 158036 32668
rect 158060 32666 158116 32668
rect 157820 32614 157846 32666
rect 157846 32614 157876 32666
rect 157900 32614 157910 32666
rect 157910 32614 157956 32666
rect 157980 32614 158026 32666
rect 158026 32614 158036 32666
rect 158060 32614 158090 32666
rect 158090 32614 158116 32666
rect 157820 32612 157876 32614
rect 157900 32612 157956 32614
rect 157980 32612 158036 32614
rect 158060 32612 158116 32614
rect 173180 32122 173236 32124
rect 173260 32122 173316 32124
rect 173340 32122 173396 32124
rect 173420 32122 173476 32124
rect 173180 32070 173206 32122
rect 173206 32070 173236 32122
rect 173260 32070 173270 32122
rect 173270 32070 173316 32122
rect 173340 32070 173386 32122
rect 173386 32070 173396 32122
rect 173420 32070 173450 32122
rect 173450 32070 173476 32122
rect 173180 32068 173236 32070
rect 173260 32068 173316 32070
rect 173340 32068 173396 32070
rect 173420 32068 173476 32070
rect 157820 31578 157876 31580
rect 157900 31578 157956 31580
rect 157980 31578 158036 31580
rect 158060 31578 158116 31580
rect 157820 31526 157846 31578
rect 157846 31526 157876 31578
rect 157900 31526 157910 31578
rect 157910 31526 157956 31578
rect 157980 31526 158026 31578
rect 158026 31526 158036 31578
rect 158060 31526 158090 31578
rect 158090 31526 158116 31578
rect 157820 31524 157876 31526
rect 157900 31524 157956 31526
rect 157980 31524 158036 31526
rect 158060 31524 158116 31526
rect 173180 31034 173236 31036
rect 173260 31034 173316 31036
rect 173340 31034 173396 31036
rect 173420 31034 173476 31036
rect 173180 30982 173206 31034
rect 173206 30982 173236 31034
rect 173260 30982 173270 31034
rect 173270 30982 173316 31034
rect 173340 30982 173386 31034
rect 173386 30982 173396 31034
rect 173420 30982 173450 31034
rect 173450 30982 173476 31034
rect 173180 30980 173236 30982
rect 173260 30980 173316 30982
rect 173340 30980 173396 30982
rect 173420 30980 173476 30982
rect 157820 30490 157876 30492
rect 157900 30490 157956 30492
rect 157980 30490 158036 30492
rect 158060 30490 158116 30492
rect 157820 30438 157846 30490
rect 157846 30438 157876 30490
rect 157900 30438 157910 30490
rect 157910 30438 157956 30490
rect 157980 30438 158026 30490
rect 158026 30438 158036 30490
rect 158060 30438 158090 30490
rect 158090 30438 158116 30490
rect 157820 30436 157876 30438
rect 157900 30436 157956 30438
rect 157980 30436 158036 30438
rect 158060 30436 158116 30438
rect 173180 29946 173236 29948
rect 173260 29946 173316 29948
rect 173340 29946 173396 29948
rect 173420 29946 173476 29948
rect 173180 29894 173206 29946
rect 173206 29894 173236 29946
rect 173260 29894 173270 29946
rect 173270 29894 173316 29946
rect 173340 29894 173386 29946
rect 173386 29894 173396 29946
rect 173420 29894 173450 29946
rect 173450 29894 173476 29946
rect 173180 29892 173236 29894
rect 173260 29892 173316 29894
rect 173340 29892 173396 29894
rect 173420 29892 173476 29894
rect 157820 29402 157876 29404
rect 157900 29402 157956 29404
rect 157980 29402 158036 29404
rect 158060 29402 158116 29404
rect 157820 29350 157846 29402
rect 157846 29350 157876 29402
rect 157900 29350 157910 29402
rect 157910 29350 157956 29402
rect 157980 29350 158026 29402
rect 158026 29350 158036 29402
rect 158060 29350 158090 29402
rect 158090 29350 158116 29402
rect 157820 29348 157876 29350
rect 157900 29348 157956 29350
rect 157980 29348 158036 29350
rect 158060 29348 158116 29350
rect 173180 28858 173236 28860
rect 173260 28858 173316 28860
rect 173340 28858 173396 28860
rect 173420 28858 173476 28860
rect 173180 28806 173206 28858
rect 173206 28806 173236 28858
rect 173260 28806 173270 28858
rect 173270 28806 173316 28858
rect 173340 28806 173386 28858
rect 173386 28806 173396 28858
rect 173420 28806 173450 28858
rect 173450 28806 173476 28858
rect 173180 28804 173236 28806
rect 173260 28804 173316 28806
rect 173340 28804 173396 28806
rect 173420 28804 173476 28806
rect 157820 28314 157876 28316
rect 157900 28314 157956 28316
rect 157980 28314 158036 28316
rect 158060 28314 158116 28316
rect 157820 28262 157846 28314
rect 157846 28262 157876 28314
rect 157900 28262 157910 28314
rect 157910 28262 157956 28314
rect 157980 28262 158026 28314
rect 158026 28262 158036 28314
rect 158060 28262 158090 28314
rect 158090 28262 158116 28314
rect 157820 28260 157876 28262
rect 157900 28260 157956 28262
rect 157980 28260 158036 28262
rect 158060 28260 158116 28262
rect 173180 27770 173236 27772
rect 173260 27770 173316 27772
rect 173340 27770 173396 27772
rect 173420 27770 173476 27772
rect 173180 27718 173206 27770
rect 173206 27718 173236 27770
rect 173260 27718 173270 27770
rect 173270 27718 173316 27770
rect 173340 27718 173386 27770
rect 173386 27718 173396 27770
rect 173420 27718 173450 27770
rect 173450 27718 173476 27770
rect 173180 27716 173236 27718
rect 173260 27716 173316 27718
rect 173340 27716 173396 27718
rect 173420 27716 173476 27718
rect 157820 27226 157876 27228
rect 157900 27226 157956 27228
rect 157980 27226 158036 27228
rect 158060 27226 158116 27228
rect 157820 27174 157846 27226
rect 157846 27174 157876 27226
rect 157900 27174 157910 27226
rect 157910 27174 157956 27226
rect 157980 27174 158026 27226
rect 158026 27174 158036 27226
rect 158060 27174 158090 27226
rect 158090 27174 158116 27226
rect 157820 27172 157876 27174
rect 157900 27172 157956 27174
rect 157980 27172 158036 27174
rect 158060 27172 158116 27174
rect 173180 26682 173236 26684
rect 173260 26682 173316 26684
rect 173340 26682 173396 26684
rect 173420 26682 173476 26684
rect 173180 26630 173206 26682
rect 173206 26630 173236 26682
rect 173260 26630 173270 26682
rect 173270 26630 173316 26682
rect 173340 26630 173386 26682
rect 173386 26630 173396 26682
rect 173420 26630 173450 26682
rect 173450 26630 173476 26682
rect 173180 26628 173236 26630
rect 173260 26628 173316 26630
rect 173340 26628 173396 26630
rect 173420 26628 173476 26630
rect 157820 26138 157876 26140
rect 157900 26138 157956 26140
rect 157980 26138 158036 26140
rect 158060 26138 158116 26140
rect 157820 26086 157846 26138
rect 157846 26086 157876 26138
rect 157900 26086 157910 26138
rect 157910 26086 157956 26138
rect 157980 26086 158026 26138
rect 158026 26086 158036 26138
rect 158060 26086 158090 26138
rect 158090 26086 158116 26138
rect 157820 26084 157876 26086
rect 157900 26084 157956 26086
rect 157980 26084 158036 26086
rect 158060 26084 158116 26086
rect 173180 25594 173236 25596
rect 173260 25594 173316 25596
rect 173340 25594 173396 25596
rect 173420 25594 173476 25596
rect 173180 25542 173206 25594
rect 173206 25542 173236 25594
rect 173260 25542 173270 25594
rect 173270 25542 173316 25594
rect 173340 25542 173386 25594
rect 173386 25542 173396 25594
rect 173420 25542 173450 25594
rect 173450 25542 173476 25594
rect 173180 25540 173236 25542
rect 173260 25540 173316 25542
rect 173340 25540 173396 25542
rect 173420 25540 173476 25542
rect 157820 25050 157876 25052
rect 157900 25050 157956 25052
rect 157980 25050 158036 25052
rect 158060 25050 158116 25052
rect 157820 24998 157846 25050
rect 157846 24998 157876 25050
rect 157900 24998 157910 25050
rect 157910 24998 157956 25050
rect 157980 24998 158026 25050
rect 158026 24998 158036 25050
rect 158060 24998 158090 25050
rect 158090 24998 158116 25050
rect 157820 24996 157876 24998
rect 157900 24996 157956 24998
rect 157980 24996 158036 24998
rect 158060 24996 158116 24998
rect 173180 24506 173236 24508
rect 173260 24506 173316 24508
rect 173340 24506 173396 24508
rect 173420 24506 173476 24508
rect 173180 24454 173206 24506
rect 173206 24454 173236 24506
rect 173260 24454 173270 24506
rect 173270 24454 173316 24506
rect 173340 24454 173386 24506
rect 173386 24454 173396 24506
rect 173420 24454 173450 24506
rect 173450 24454 173476 24506
rect 173180 24452 173236 24454
rect 173260 24452 173316 24454
rect 173340 24452 173396 24454
rect 173420 24452 173476 24454
rect 157820 23962 157876 23964
rect 157900 23962 157956 23964
rect 157980 23962 158036 23964
rect 158060 23962 158116 23964
rect 157820 23910 157846 23962
rect 157846 23910 157876 23962
rect 157900 23910 157910 23962
rect 157910 23910 157956 23962
rect 157980 23910 158026 23962
rect 158026 23910 158036 23962
rect 158060 23910 158090 23962
rect 158090 23910 158116 23962
rect 157820 23908 157876 23910
rect 157900 23908 157956 23910
rect 157980 23908 158036 23910
rect 158060 23908 158116 23910
rect 173180 23418 173236 23420
rect 173260 23418 173316 23420
rect 173340 23418 173396 23420
rect 173420 23418 173476 23420
rect 173180 23366 173206 23418
rect 173206 23366 173236 23418
rect 173260 23366 173270 23418
rect 173270 23366 173316 23418
rect 173340 23366 173386 23418
rect 173386 23366 173396 23418
rect 173420 23366 173450 23418
rect 173450 23366 173476 23418
rect 173180 23364 173236 23366
rect 173260 23364 173316 23366
rect 173340 23364 173396 23366
rect 173420 23364 173476 23366
rect 157820 22874 157876 22876
rect 157900 22874 157956 22876
rect 157980 22874 158036 22876
rect 158060 22874 158116 22876
rect 157820 22822 157846 22874
rect 157846 22822 157876 22874
rect 157900 22822 157910 22874
rect 157910 22822 157956 22874
rect 157980 22822 158026 22874
rect 158026 22822 158036 22874
rect 158060 22822 158090 22874
rect 158090 22822 158116 22874
rect 157820 22820 157876 22822
rect 157900 22820 157956 22822
rect 157980 22820 158036 22822
rect 158060 22820 158116 22822
rect 173180 22330 173236 22332
rect 173260 22330 173316 22332
rect 173340 22330 173396 22332
rect 173420 22330 173476 22332
rect 173180 22278 173206 22330
rect 173206 22278 173236 22330
rect 173260 22278 173270 22330
rect 173270 22278 173316 22330
rect 173340 22278 173386 22330
rect 173386 22278 173396 22330
rect 173420 22278 173450 22330
rect 173450 22278 173476 22330
rect 173180 22276 173236 22278
rect 173260 22276 173316 22278
rect 173340 22276 173396 22278
rect 173420 22276 173476 22278
rect 157820 21786 157876 21788
rect 157900 21786 157956 21788
rect 157980 21786 158036 21788
rect 158060 21786 158116 21788
rect 157820 21734 157846 21786
rect 157846 21734 157876 21786
rect 157900 21734 157910 21786
rect 157910 21734 157956 21786
rect 157980 21734 158026 21786
rect 158026 21734 158036 21786
rect 158060 21734 158090 21786
rect 158090 21734 158116 21786
rect 157820 21732 157876 21734
rect 157900 21732 157956 21734
rect 157980 21732 158036 21734
rect 158060 21732 158116 21734
rect 173180 21242 173236 21244
rect 173260 21242 173316 21244
rect 173340 21242 173396 21244
rect 173420 21242 173476 21244
rect 173180 21190 173206 21242
rect 173206 21190 173236 21242
rect 173260 21190 173270 21242
rect 173270 21190 173316 21242
rect 173340 21190 173386 21242
rect 173386 21190 173396 21242
rect 173420 21190 173450 21242
rect 173450 21190 173476 21242
rect 173180 21188 173236 21190
rect 173260 21188 173316 21190
rect 173340 21188 173396 21190
rect 173420 21188 173476 21190
rect 157820 20698 157876 20700
rect 157900 20698 157956 20700
rect 157980 20698 158036 20700
rect 158060 20698 158116 20700
rect 157820 20646 157846 20698
rect 157846 20646 157876 20698
rect 157900 20646 157910 20698
rect 157910 20646 157956 20698
rect 157980 20646 158026 20698
rect 158026 20646 158036 20698
rect 158060 20646 158090 20698
rect 158090 20646 158116 20698
rect 157820 20644 157876 20646
rect 157900 20644 157956 20646
rect 157980 20644 158036 20646
rect 158060 20644 158116 20646
rect 173180 20154 173236 20156
rect 173260 20154 173316 20156
rect 173340 20154 173396 20156
rect 173420 20154 173476 20156
rect 173180 20102 173206 20154
rect 173206 20102 173236 20154
rect 173260 20102 173270 20154
rect 173270 20102 173316 20154
rect 173340 20102 173386 20154
rect 173386 20102 173396 20154
rect 173420 20102 173450 20154
rect 173450 20102 173476 20154
rect 173180 20100 173236 20102
rect 173260 20100 173316 20102
rect 173340 20100 173396 20102
rect 173420 20100 173476 20102
rect 157820 19610 157876 19612
rect 157900 19610 157956 19612
rect 157980 19610 158036 19612
rect 158060 19610 158116 19612
rect 157820 19558 157846 19610
rect 157846 19558 157876 19610
rect 157900 19558 157910 19610
rect 157910 19558 157956 19610
rect 157980 19558 158026 19610
rect 158026 19558 158036 19610
rect 158060 19558 158090 19610
rect 158090 19558 158116 19610
rect 157820 19556 157876 19558
rect 157900 19556 157956 19558
rect 157980 19556 158036 19558
rect 158060 19556 158116 19558
rect 173180 19066 173236 19068
rect 173260 19066 173316 19068
rect 173340 19066 173396 19068
rect 173420 19066 173476 19068
rect 173180 19014 173206 19066
rect 173206 19014 173236 19066
rect 173260 19014 173270 19066
rect 173270 19014 173316 19066
rect 173340 19014 173386 19066
rect 173386 19014 173396 19066
rect 173420 19014 173450 19066
rect 173450 19014 173476 19066
rect 173180 19012 173236 19014
rect 173260 19012 173316 19014
rect 173340 19012 173396 19014
rect 173420 19012 173476 19014
rect 96380 18522 96436 18524
rect 96460 18522 96516 18524
rect 96540 18522 96596 18524
rect 96620 18522 96676 18524
rect 96380 18470 96406 18522
rect 96406 18470 96436 18522
rect 96460 18470 96470 18522
rect 96470 18470 96516 18522
rect 96540 18470 96586 18522
rect 96586 18470 96596 18522
rect 96620 18470 96650 18522
rect 96650 18470 96676 18522
rect 96380 18468 96436 18470
rect 96460 18468 96516 18470
rect 96540 18468 96596 18470
rect 96620 18468 96676 18470
rect 127100 18522 127156 18524
rect 127180 18522 127236 18524
rect 127260 18522 127316 18524
rect 127340 18522 127396 18524
rect 127100 18470 127126 18522
rect 127126 18470 127156 18522
rect 127180 18470 127190 18522
rect 127190 18470 127236 18522
rect 127260 18470 127306 18522
rect 127306 18470 127316 18522
rect 127340 18470 127370 18522
rect 127370 18470 127396 18522
rect 127100 18468 127156 18470
rect 127180 18468 127236 18470
rect 127260 18468 127316 18470
rect 127340 18468 127396 18470
rect 157820 18522 157876 18524
rect 157900 18522 157956 18524
rect 157980 18522 158036 18524
rect 158060 18522 158116 18524
rect 157820 18470 157846 18522
rect 157846 18470 157876 18522
rect 157900 18470 157910 18522
rect 157910 18470 157956 18522
rect 157980 18470 158026 18522
rect 158026 18470 158036 18522
rect 158060 18470 158090 18522
rect 158090 18470 158116 18522
rect 157820 18468 157876 18470
rect 157900 18468 157956 18470
rect 157980 18468 158036 18470
rect 158060 18468 158116 18470
rect 81020 17978 81076 17980
rect 81100 17978 81156 17980
rect 81180 17978 81236 17980
rect 81260 17978 81316 17980
rect 81020 17926 81046 17978
rect 81046 17926 81076 17978
rect 81100 17926 81110 17978
rect 81110 17926 81156 17978
rect 81180 17926 81226 17978
rect 81226 17926 81236 17978
rect 81260 17926 81290 17978
rect 81290 17926 81316 17978
rect 81020 17924 81076 17926
rect 81100 17924 81156 17926
rect 81180 17924 81236 17926
rect 81260 17924 81316 17926
rect 111740 17978 111796 17980
rect 111820 17978 111876 17980
rect 111900 17978 111956 17980
rect 111980 17978 112036 17980
rect 111740 17926 111766 17978
rect 111766 17926 111796 17978
rect 111820 17926 111830 17978
rect 111830 17926 111876 17978
rect 111900 17926 111946 17978
rect 111946 17926 111956 17978
rect 111980 17926 112010 17978
rect 112010 17926 112036 17978
rect 111740 17924 111796 17926
rect 111820 17924 111876 17926
rect 111900 17924 111956 17926
rect 111980 17924 112036 17926
rect 142460 17978 142516 17980
rect 142540 17978 142596 17980
rect 142620 17978 142676 17980
rect 142700 17978 142756 17980
rect 142460 17926 142486 17978
rect 142486 17926 142516 17978
rect 142540 17926 142550 17978
rect 142550 17926 142596 17978
rect 142620 17926 142666 17978
rect 142666 17926 142676 17978
rect 142700 17926 142730 17978
rect 142730 17926 142756 17978
rect 142460 17924 142516 17926
rect 142540 17924 142596 17926
rect 142620 17924 142676 17926
rect 142700 17924 142756 17926
rect 173180 17978 173236 17980
rect 173260 17978 173316 17980
rect 173340 17978 173396 17980
rect 173420 17978 173476 17980
rect 173180 17926 173206 17978
rect 173206 17926 173236 17978
rect 173260 17926 173270 17978
rect 173270 17926 173316 17978
rect 173340 17926 173386 17978
rect 173386 17926 173396 17978
rect 173420 17926 173450 17978
rect 173450 17926 173476 17978
rect 173180 17924 173236 17926
rect 173260 17924 173316 17926
rect 173340 17924 173396 17926
rect 173420 17924 173476 17926
rect 96380 17434 96436 17436
rect 96460 17434 96516 17436
rect 96540 17434 96596 17436
rect 96620 17434 96676 17436
rect 96380 17382 96406 17434
rect 96406 17382 96436 17434
rect 96460 17382 96470 17434
rect 96470 17382 96516 17434
rect 96540 17382 96586 17434
rect 96586 17382 96596 17434
rect 96620 17382 96650 17434
rect 96650 17382 96676 17434
rect 96380 17380 96436 17382
rect 96460 17380 96516 17382
rect 96540 17380 96596 17382
rect 96620 17380 96676 17382
rect 127100 17434 127156 17436
rect 127180 17434 127236 17436
rect 127260 17434 127316 17436
rect 127340 17434 127396 17436
rect 127100 17382 127126 17434
rect 127126 17382 127156 17434
rect 127180 17382 127190 17434
rect 127190 17382 127236 17434
rect 127260 17382 127306 17434
rect 127306 17382 127316 17434
rect 127340 17382 127370 17434
rect 127370 17382 127396 17434
rect 127100 17380 127156 17382
rect 127180 17380 127236 17382
rect 127260 17380 127316 17382
rect 127340 17380 127396 17382
rect 157820 17434 157876 17436
rect 157900 17434 157956 17436
rect 157980 17434 158036 17436
rect 158060 17434 158116 17436
rect 157820 17382 157846 17434
rect 157846 17382 157876 17434
rect 157900 17382 157910 17434
rect 157910 17382 157956 17434
rect 157980 17382 158026 17434
rect 158026 17382 158036 17434
rect 158060 17382 158090 17434
rect 158090 17382 158116 17434
rect 157820 17380 157876 17382
rect 157900 17380 157956 17382
rect 157980 17380 158036 17382
rect 158060 17380 158116 17382
rect 81020 16890 81076 16892
rect 81100 16890 81156 16892
rect 81180 16890 81236 16892
rect 81260 16890 81316 16892
rect 81020 16838 81046 16890
rect 81046 16838 81076 16890
rect 81100 16838 81110 16890
rect 81110 16838 81156 16890
rect 81180 16838 81226 16890
rect 81226 16838 81236 16890
rect 81260 16838 81290 16890
rect 81290 16838 81316 16890
rect 81020 16836 81076 16838
rect 81100 16836 81156 16838
rect 81180 16836 81236 16838
rect 81260 16836 81316 16838
rect 111740 16890 111796 16892
rect 111820 16890 111876 16892
rect 111900 16890 111956 16892
rect 111980 16890 112036 16892
rect 111740 16838 111766 16890
rect 111766 16838 111796 16890
rect 111820 16838 111830 16890
rect 111830 16838 111876 16890
rect 111900 16838 111946 16890
rect 111946 16838 111956 16890
rect 111980 16838 112010 16890
rect 112010 16838 112036 16890
rect 111740 16836 111796 16838
rect 111820 16836 111876 16838
rect 111900 16836 111956 16838
rect 111980 16836 112036 16838
rect 142460 16890 142516 16892
rect 142540 16890 142596 16892
rect 142620 16890 142676 16892
rect 142700 16890 142756 16892
rect 142460 16838 142486 16890
rect 142486 16838 142516 16890
rect 142540 16838 142550 16890
rect 142550 16838 142596 16890
rect 142620 16838 142666 16890
rect 142666 16838 142676 16890
rect 142700 16838 142730 16890
rect 142730 16838 142756 16890
rect 142460 16836 142516 16838
rect 142540 16836 142596 16838
rect 142620 16836 142676 16838
rect 142700 16836 142756 16838
rect 173180 16890 173236 16892
rect 173260 16890 173316 16892
rect 173340 16890 173396 16892
rect 173420 16890 173476 16892
rect 173180 16838 173206 16890
rect 173206 16838 173236 16890
rect 173260 16838 173270 16890
rect 173270 16838 173316 16890
rect 173340 16838 173386 16890
rect 173386 16838 173396 16890
rect 173420 16838 173450 16890
rect 173450 16838 173476 16890
rect 173180 16836 173236 16838
rect 173260 16836 173316 16838
rect 173340 16836 173396 16838
rect 173420 16836 173476 16838
rect 96380 16346 96436 16348
rect 96460 16346 96516 16348
rect 96540 16346 96596 16348
rect 96620 16346 96676 16348
rect 96380 16294 96406 16346
rect 96406 16294 96436 16346
rect 96460 16294 96470 16346
rect 96470 16294 96516 16346
rect 96540 16294 96586 16346
rect 96586 16294 96596 16346
rect 96620 16294 96650 16346
rect 96650 16294 96676 16346
rect 96380 16292 96436 16294
rect 96460 16292 96516 16294
rect 96540 16292 96596 16294
rect 96620 16292 96676 16294
rect 127100 16346 127156 16348
rect 127180 16346 127236 16348
rect 127260 16346 127316 16348
rect 127340 16346 127396 16348
rect 127100 16294 127126 16346
rect 127126 16294 127156 16346
rect 127180 16294 127190 16346
rect 127190 16294 127236 16346
rect 127260 16294 127306 16346
rect 127306 16294 127316 16346
rect 127340 16294 127370 16346
rect 127370 16294 127396 16346
rect 127100 16292 127156 16294
rect 127180 16292 127236 16294
rect 127260 16292 127316 16294
rect 127340 16292 127396 16294
rect 157820 16346 157876 16348
rect 157900 16346 157956 16348
rect 157980 16346 158036 16348
rect 158060 16346 158116 16348
rect 157820 16294 157846 16346
rect 157846 16294 157876 16346
rect 157900 16294 157910 16346
rect 157910 16294 157956 16346
rect 157980 16294 158026 16346
rect 158026 16294 158036 16346
rect 158060 16294 158090 16346
rect 158090 16294 158116 16346
rect 157820 16292 157876 16294
rect 157900 16292 157956 16294
rect 157980 16292 158036 16294
rect 158060 16292 158116 16294
rect 81020 15802 81076 15804
rect 81100 15802 81156 15804
rect 81180 15802 81236 15804
rect 81260 15802 81316 15804
rect 81020 15750 81046 15802
rect 81046 15750 81076 15802
rect 81100 15750 81110 15802
rect 81110 15750 81156 15802
rect 81180 15750 81226 15802
rect 81226 15750 81236 15802
rect 81260 15750 81290 15802
rect 81290 15750 81316 15802
rect 81020 15748 81076 15750
rect 81100 15748 81156 15750
rect 81180 15748 81236 15750
rect 81260 15748 81316 15750
rect 111740 15802 111796 15804
rect 111820 15802 111876 15804
rect 111900 15802 111956 15804
rect 111980 15802 112036 15804
rect 111740 15750 111766 15802
rect 111766 15750 111796 15802
rect 111820 15750 111830 15802
rect 111830 15750 111876 15802
rect 111900 15750 111946 15802
rect 111946 15750 111956 15802
rect 111980 15750 112010 15802
rect 112010 15750 112036 15802
rect 111740 15748 111796 15750
rect 111820 15748 111876 15750
rect 111900 15748 111956 15750
rect 111980 15748 112036 15750
rect 142460 15802 142516 15804
rect 142540 15802 142596 15804
rect 142620 15802 142676 15804
rect 142700 15802 142756 15804
rect 142460 15750 142486 15802
rect 142486 15750 142516 15802
rect 142540 15750 142550 15802
rect 142550 15750 142596 15802
rect 142620 15750 142666 15802
rect 142666 15750 142676 15802
rect 142700 15750 142730 15802
rect 142730 15750 142756 15802
rect 142460 15748 142516 15750
rect 142540 15748 142596 15750
rect 142620 15748 142676 15750
rect 142700 15748 142756 15750
rect 173180 15802 173236 15804
rect 173260 15802 173316 15804
rect 173340 15802 173396 15804
rect 173420 15802 173476 15804
rect 173180 15750 173206 15802
rect 173206 15750 173236 15802
rect 173260 15750 173270 15802
rect 173270 15750 173316 15802
rect 173340 15750 173386 15802
rect 173386 15750 173396 15802
rect 173420 15750 173450 15802
rect 173450 15750 173476 15802
rect 173180 15748 173236 15750
rect 173260 15748 173316 15750
rect 173340 15748 173396 15750
rect 173420 15748 173476 15750
rect 96380 15258 96436 15260
rect 96460 15258 96516 15260
rect 96540 15258 96596 15260
rect 96620 15258 96676 15260
rect 96380 15206 96406 15258
rect 96406 15206 96436 15258
rect 96460 15206 96470 15258
rect 96470 15206 96516 15258
rect 96540 15206 96586 15258
rect 96586 15206 96596 15258
rect 96620 15206 96650 15258
rect 96650 15206 96676 15258
rect 96380 15204 96436 15206
rect 96460 15204 96516 15206
rect 96540 15204 96596 15206
rect 96620 15204 96676 15206
rect 127100 15258 127156 15260
rect 127180 15258 127236 15260
rect 127260 15258 127316 15260
rect 127340 15258 127396 15260
rect 127100 15206 127126 15258
rect 127126 15206 127156 15258
rect 127180 15206 127190 15258
rect 127190 15206 127236 15258
rect 127260 15206 127306 15258
rect 127306 15206 127316 15258
rect 127340 15206 127370 15258
rect 127370 15206 127396 15258
rect 127100 15204 127156 15206
rect 127180 15204 127236 15206
rect 127260 15204 127316 15206
rect 127340 15204 127396 15206
rect 157820 15258 157876 15260
rect 157900 15258 157956 15260
rect 157980 15258 158036 15260
rect 158060 15258 158116 15260
rect 157820 15206 157846 15258
rect 157846 15206 157876 15258
rect 157900 15206 157910 15258
rect 157910 15206 157956 15258
rect 157980 15206 158026 15258
rect 158026 15206 158036 15258
rect 158060 15206 158090 15258
rect 158090 15206 158116 15258
rect 157820 15204 157876 15206
rect 157900 15204 157956 15206
rect 157980 15204 158036 15206
rect 158060 15204 158116 15206
rect 81020 14714 81076 14716
rect 81100 14714 81156 14716
rect 81180 14714 81236 14716
rect 81260 14714 81316 14716
rect 81020 14662 81046 14714
rect 81046 14662 81076 14714
rect 81100 14662 81110 14714
rect 81110 14662 81156 14714
rect 81180 14662 81226 14714
rect 81226 14662 81236 14714
rect 81260 14662 81290 14714
rect 81290 14662 81316 14714
rect 81020 14660 81076 14662
rect 81100 14660 81156 14662
rect 81180 14660 81236 14662
rect 81260 14660 81316 14662
rect 111740 14714 111796 14716
rect 111820 14714 111876 14716
rect 111900 14714 111956 14716
rect 111980 14714 112036 14716
rect 111740 14662 111766 14714
rect 111766 14662 111796 14714
rect 111820 14662 111830 14714
rect 111830 14662 111876 14714
rect 111900 14662 111946 14714
rect 111946 14662 111956 14714
rect 111980 14662 112010 14714
rect 112010 14662 112036 14714
rect 111740 14660 111796 14662
rect 111820 14660 111876 14662
rect 111900 14660 111956 14662
rect 111980 14660 112036 14662
rect 142460 14714 142516 14716
rect 142540 14714 142596 14716
rect 142620 14714 142676 14716
rect 142700 14714 142756 14716
rect 142460 14662 142486 14714
rect 142486 14662 142516 14714
rect 142540 14662 142550 14714
rect 142550 14662 142596 14714
rect 142620 14662 142666 14714
rect 142666 14662 142676 14714
rect 142700 14662 142730 14714
rect 142730 14662 142756 14714
rect 142460 14660 142516 14662
rect 142540 14660 142596 14662
rect 142620 14660 142676 14662
rect 142700 14660 142756 14662
rect 173180 14714 173236 14716
rect 173260 14714 173316 14716
rect 173340 14714 173396 14716
rect 173420 14714 173476 14716
rect 173180 14662 173206 14714
rect 173206 14662 173236 14714
rect 173260 14662 173270 14714
rect 173270 14662 173316 14714
rect 173340 14662 173386 14714
rect 173386 14662 173396 14714
rect 173420 14662 173450 14714
rect 173450 14662 173476 14714
rect 173180 14660 173236 14662
rect 173260 14660 173316 14662
rect 173340 14660 173396 14662
rect 173420 14660 173476 14662
rect 96380 14170 96436 14172
rect 96460 14170 96516 14172
rect 96540 14170 96596 14172
rect 96620 14170 96676 14172
rect 96380 14118 96406 14170
rect 96406 14118 96436 14170
rect 96460 14118 96470 14170
rect 96470 14118 96516 14170
rect 96540 14118 96586 14170
rect 96586 14118 96596 14170
rect 96620 14118 96650 14170
rect 96650 14118 96676 14170
rect 96380 14116 96436 14118
rect 96460 14116 96516 14118
rect 96540 14116 96596 14118
rect 96620 14116 96676 14118
rect 81020 13626 81076 13628
rect 81100 13626 81156 13628
rect 81180 13626 81236 13628
rect 81260 13626 81316 13628
rect 81020 13574 81046 13626
rect 81046 13574 81076 13626
rect 81100 13574 81110 13626
rect 81110 13574 81156 13626
rect 81180 13574 81226 13626
rect 81226 13574 81236 13626
rect 81260 13574 81290 13626
rect 81290 13574 81316 13626
rect 81020 13572 81076 13574
rect 81100 13572 81156 13574
rect 81180 13572 81236 13574
rect 81260 13572 81316 13574
rect 70398 6160 70454 6216
rect 70030 3068 70032 3088
rect 70032 3068 70084 3088
rect 70084 3068 70086 3088
rect 70030 3032 70086 3068
rect 70490 2896 70546 2952
rect 70674 3168 70730 3224
rect 71502 3884 71504 3904
rect 71504 3884 71556 3904
rect 71556 3884 71558 3904
rect 71502 3848 71558 3884
rect 71318 2916 71374 2952
rect 71318 2896 71320 2916
rect 71320 2896 71372 2916
rect 71372 2896 71374 2916
rect 71962 3032 72018 3088
rect 72146 3576 72202 3632
rect 73250 6160 73306 6216
rect 73250 3984 73306 4040
rect 73434 3032 73490 3088
rect 96380 13082 96436 13084
rect 96460 13082 96516 13084
rect 96540 13082 96596 13084
rect 96620 13082 96676 13084
rect 96380 13030 96406 13082
rect 96406 13030 96436 13082
rect 96460 13030 96470 13082
rect 96470 13030 96516 13082
rect 96540 13030 96586 13082
rect 96586 13030 96596 13082
rect 96620 13030 96650 13082
rect 96650 13030 96676 13082
rect 96380 13028 96436 13030
rect 96460 13028 96516 13030
rect 96540 13028 96596 13030
rect 96620 13028 96676 13030
rect 81020 12538 81076 12540
rect 81100 12538 81156 12540
rect 81180 12538 81236 12540
rect 81260 12538 81316 12540
rect 81020 12486 81046 12538
rect 81046 12486 81076 12538
rect 81100 12486 81110 12538
rect 81110 12486 81156 12538
rect 81180 12486 81226 12538
rect 81226 12486 81236 12538
rect 81260 12486 81290 12538
rect 81290 12486 81316 12538
rect 81020 12484 81076 12486
rect 81100 12484 81156 12486
rect 81180 12484 81236 12486
rect 81260 12484 81316 12486
rect 81020 11450 81076 11452
rect 81100 11450 81156 11452
rect 81180 11450 81236 11452
rect 81260 11450 81316 11452
rect 81020 11398 81046 11450
rect 81046 11398 81076 11450
rect 81100 11398 81110 11450
rect 81110 11398 81156 11450
rect 81180 11398 81226 11450
rect 81226 11398 81236 11450
rect 81260 11398 81290 11450
rect 81290 11398 81316 11450
rect 81020 11396 81076 11398
rect 81100 11396 81156 11398
rect 81180 11396 81236 11398
rect 81260 11396 81316 11398
rect 81020 10362 81076 10364
rect 81100 10362 81156 10364
rect 81180 10362 81236 10364
rect 81260 10362 81316 10364
rect 81020 10310 81046 10362
rect 81046 10310 81076 10362
rect 81100 10310 81110 10362
rect 81110 10310 81156 10362
rect 81180 10310 81226 10362
rect 81226 10310 81236 10362
rect 81260 10310 81290 10362
rect 81290 10310 81316 10362
rect 81020 10308 81076 10310
rect 81100 10308 81156 10310
rect 81180 10308 81236 10310
rect 81260 10308 81316 10310
rect 81020 9274 81076 9276
rect 81100 9274 81156 9276
rect 81180 9274 81236 9276
rect 81260 9274 81316 9276
rect 81020 9222 81046 9274
rect 81046 9222 81076 9274
rect 81100 9222 81110 9274
rect 81110 9222 81156 9274
rect 81180 9222 81226 9274
rect 81226 9222 81236 9274
rect 81260 9222 81290 9274
rect 81290 9222 81316 9274
rect 81020 9220 81076 9222
rect 81100 9220 81156 9222
rect 81180 9220 81236 9222
rect 81260 9220 81316 9222
rect 81020 8186 81076 8188
rect 81100 8186 81156 8188
rect 81180 8186 81236 8188
rect 81260 8186 81316 8188
rect 81020 8134 81046 8186
rect 81046 8134 81076 8186
rect 81100 8134 81110 8186
rect 81110 8134 81156 8186
rect 81180 8134 81226 8186
rect 81226 8134 81236 8186
rect 81260 8134 81290 8186
rect 81290 8134 81316 8186
rect 81020 8132 81076 8134
rect 81100 8132 81156 8134
rect 81180 8132 81236 8134
rect 81260 8132 81316 8134
rect 81020 7098 81076 7100
rect 81100 7098 81156 7100
rect 81180 7098 81236 7100
rect 81260 7098 81316 7100
rect 81020 7046 81046 7098
rect 81046 7046 81076 7098
rect 81100 7046 81110 7098
rect 81110 7046 81156 7098
rect 81180 7046 81226 7098
rect 81226 7046 81236 7098
rect 81260 7046 81290 7098
rect 81290 7046 81316 7098
rect 81020 7044 81076 7046
rect 81100 7044 81156 7046
rect 81180 7044 81236 7046
rect 81260 7044 81316 7046
rect 74630 2896 74686 2952
rect 74906 2352 74962 2408
rect 75090 3440 75146 3496
rect 75274 4528 75330 4584
rect 75550 3032 75606 3088
rect 75826 3576 75882 3632
rect 75642 2760 75698 2816
rect 75826 3476 75828 3496
rect 75828 3476 75880 3496
rect 75880 3476 75882 3496
rect 75826 3440 75882 3476
rect 76286 3612 76288 3632
rect 76288 3612 76340 3632
rect 76340 3612 76342 3632
rect 76286 3576 76342 3612
rect 76654 3032 76710 3088
rect 77390 3304 77446 3360
rect 77850 3848 77906 3904
rect 77758 3304 77814 3360
rect 78402 4392 78458 4448
rect 78586 3168 78642 3224
rect 79046 5616 79102 5672
rect 78862 5344 78918 5400
rect 79046 3304 79102 3360
rect 78770 3168 78826 3224
rect 78862 2624 78918 2680
rect 79046 2916 79102 2952
rect 79046 2896 79048 2916
rect 79048 2896 79100 2916
rect 79100 2896 79102 2916
rect 79690 4256 79746 4312
rect 79414 4120 79470 4176
rect 79690 3712 79746 3768
rect 79690 2796 79692 2816
rect 79692 2796 79744 2816
rect 79744 2796 79746 2816
rect 79690 2760 79746 2796
rect 78954 2216 79010 2272
rect 80334 5072 80390 5128
rect 79874 3440 79930 3496
rect 80426 4256 80482 4312
rect 80426 2080 80482 2136
rect 80610 3460 80666 3496
rect 80610 3440 80612 3460
rect 80612 3440 80664 3460
rect 80664 3440 80666 3460
rect 81020 6010 81076 6012
rect 81100 6010 81156 6012
rect 81180 6010 81236 6012
rect 81260 6010 81316 6012
rect 81020 5958 81046 6010
rect 81046 5958 81076 6010
rect 81100 5958 81110 6010
rect 81110 5958 81156 6010
rect 81180 5958 81226 6010
rect 81226 5958 81236 6010
rect 81260 5958 81290 6010
rect 81290 5958 81316 6010
rect 81020 5956 81076 5958
rect 81100 5956 81156 5958
rect 81180 5956 81236 5958
rect 81260 5956 81316 5958
rect 81020 4922 81076 4924
rect 81100 4922 81156 4924
rect 81180 4922 81236 4924
rect 81260 4922 81316 4924
rect 81020 4870 81046 4922
rect 81046 4870 81076 4922
rect 81100 4870 81110 4922
rect 81110 4870 81156 4922
rect 81180 4870 81226 4922
rect 81226 4870 81236 4922
rect 81260 4870 81290 4922
rect 81290 4870 81316 4922
rect 81020 4868 81076 4870
rect 81100 4868 81156 4870
rect 81180 4868 81236 4870
rect 81260 4868 81316 4870
rect 81020 3834 81076 3836
rect 81100 3834 81156 3836
rect 81180 3834 81236 3836
rect 81260 3834 81316 3836
rect 81020 3782 81046 3834
rect 81046 3782 81076 3834
rect 81100 3782 81110 3834
rect 81110 3782 81156 3834
rect 81180 3782 81226 3834
rect 81226 3782 81236 3834
rect 81260 3782 81290 3834
rect 81290 3782 81316 3834
rect 81020 3780 81076 3782
rect 81100 3780 81156 3782
rect 81180 3780 81236 3782
rect 81260 3780 81316 3782
rect 81070 3440 81126 3496
rect 80886 2760 80942 2816
rect 81020 2746 81076 2748
rect 81100 2746 81156 2748
rect 81180 2746 81236 2748
rect 81260 2746 81316 2748
rect 81020 2694 81046 2746
rect 81046 2694 81076 2746
rect 81100 2694 81110 2746
rect 81110 2694 81156 2746
rect 81180 2694 81226 2746
rect 81226 2694 81236 2746
rect 81260 2694 81290 2746
rect 81290 2694 81316 2746
rect 81020 2692 81076 2694
rect 81100 2692 81156 2694
rect 81180 2692 81236 2694
rect 81260 2692 81316 2694
rect 81806 5208 81862 5264
rect 81714 4800 81770 4856
rect 81714 2624 81770 2680
rect 82542 5752 82598 5808
rect 82266 5092 82322 5128
rect 82266 5072 82268 5092
rect 82268 5072 82320 5092
rect 82320 5072 82322 5092
rect 82818 3848 82874 3904
rect 83002 4392 83058 4448
rect 83370 5480 83426 5536
rect 83738 5344 83794 5400
rect 83738 2760 83794 2816
rect 83186 2352 83242 2408
rect 84566 5752 84622 5808
rect 84014 5616 84070 5672
rect 83922 4392 83978 4448
rect 84198 4256 84254 4312
rect 84106 3712 84162 3768
rect 84198 2760 84254 2816
rect 84750 5364 84806 5400
rect 84750 5344 84752 5364
rect 84752 5344 84804 5364
rect 84804 5344 84806 5364
rect 84842 4936 84898 4992
rect 84842 4256 84898 4312
rect 84566 2352 84622 2408
rect 85026 5208 85082 5264
rect 85762 5480 85818 5536
rect 85394 3848 85450 3904
rect 85486 3712 85542 3768
rect 85210 2080 85266 2136
rect 85854 4392 85910 4448
rect 85670 3440 85726 3496
rect 85762 3032 85818 3088
rect 86222 3984 86278 4040
rect 86222 3884 86224 3904
rect 86224 3884 86276 3904
rect 86276 3884 86278 3904
rect 86222 3848 86278 3884
rect 86498 4664 86554 4720
rect 86774 4256 86830 4312
rect 86774 3984 86830 4040
rect 86498 3032 86554 3088
rect 86958 3032 87014 3088
rect 86406 2760 86462 2816
rect 86774 2760 86830 2816
rect 86682 2352 86738 2408
rect 86498 2080 86554 2136
rect 86774 1944 86830 2000
rect 87878 4800 87934 4856
rect 88522 4800 88578 4856
rect 87234 3068 87236 3088
rect 87236 3068 87288 3088
rect 87288 3068 87290 3088
rect 87234 3032 87290 3068
rect 87326 2760 87382 2816
rect 87602 4392 87658 4448
rect 87694 2216 87750 2272
rect 87970 4256 88026 4312
rect 87970 3304 88026 3360
rect 88062 3032 88118 3088
rect 88430 4548 88486 4584
rect 88430 4528 88432 4548
rect 88432 4528 88484 4548
rect 88484 4528 88486 4548
rect 88614 4004 88670 4040
rect 88614 3984 88616 4004
rect 88616 3984 88668 4004
rect 88668 3984 88670 4004
rect 88706 3732 88762 3768
rect 88706 3712 88708 3732
rect 88708 3712 88760 3732
rect 88760 3712 88762 3732
rect 88614 3576 88670 3632
rect 88430 3440 88486 3496
rect 89626 4800 89682 4856
rect 89166 2896 89222 2952
rect 89718 4392 89774 4448
rect 89626 2760 89682 2816
rect 92202 5072 92258 5128
rect 91006 4140 91062 4176
rect 91006 4120 91008 4140
rect 91008 4120 91060 4140
rect 91060 4120 91062 4140
rect 90822 3168 90878 3224
rect 91834 2080 91890 2136
rect 93214 3304 93270 3360
rect 93582 2216 93638 2272
rect 96380 11994 96436 11996
rect 96460 11994 96516 11996
rect 96540 11994 96596 11996
rect 96620 11994 96676 11996
rect 96380 11942 96406 11994
rect 96406 11942 96436 11994
rect 96460 11942 96470 11994
rect 96470 11942 96516 11994
rect 96540 11942 96586 11994
rect 96586 11942 96596 11994
rect 96620 11942 96650 11994
rect 96650 11942 96676 11994
rect 96380 11940 96436 11942
rect 96460 11940 96516 11942
rect 96540 11940 96596 11942
rect 96620 11940 96676 11942
rect 96380 10906 96436 10908
rect 96460 10906 96516 10908
rect 96540 10906 96596 10908
rect 96620 10906 96676 10908
rect 96380 10854 96406 10906
rect 96406 10854 96436 10906
rect 96460 10854 96470 10906
rect 96470 10854 96516 10906
rect 96540 10854 96586 10906
rect 96586 10854 96596 10906
rect 96620 10854 96650 10906
rect 96650 10854 96676 10906
rect 96380 10852 96436 10854
rect 96460 10852 96516 10854
rect 96540 10852 96596 10854
rect 96620 10852 96676 10854
rect 96380 9818 96436 9820
rect 96460 9818 96516 9820
rect 96540 9818 96596 9820
rect 96620 9818 96676 9820
rect 96380 9766 96406 9818
rect 96406 9766 96436 9818
rect 96460 9766 96470 9818
rect 96470 9766 96516 9818
rect 96540 9766 96586 9818
rect 96586 9766 96596 9818
rect 96620 9766 96650 9818
rect 96650 9766 96676 9818
rect 96380 9764 96436 9766
rect 96460 9764 96516 9766
rect 96540 9764 96596 9766
rect 96620 9764 96676 9766
rect 96380 8730 96436 8732
rect 96460 8730 96516 8732
rect 96540 8730 96596 8732
rect 96620 8730 96676 8732
rect 96380 8678 96406 8730
rect 96406 8678 96436 8730
rect 96460 8678 96470 8730
rect 96470 8678 96516 8730
rect 96540 8678 96586 8730
rect 96586 8678 96596 8730
rect 96620 8678 96650 8730
rect 96650 8678 96676 8730
rect 96380 8676 96436 8678
rect 96460 8676 96516 8678
rect 96540 8676 96596 8678
rect 96620 8676 96676 8678
rect 96380 7642 96436 7644
rect 96460 7642 96516 7644
rect 96540 7642 96596 7644
rect 96620 7642 96676 7644
rect 96380 7590 96406 7642
rect 96406 7590 96436 7642
rect 96460 7590 96470 7642
rect 96470 7590 96516 7642
rect 96540 7590 96586 7642
rect 96586 7590 96596 7642
rect 96620 7590 96650 7642
rect 96650 7590 96676 7642
rect 96380 7588 96436 7590
rect 96460 7588 96516 7590
rect 96540 7588 96596 7590
rect 96620 7588 96676 7590
rect 96380 6554 96436 6556
rect 96460 6554 96516 6556
rect 96540 6554 96596 6556
rect 96620 6554 96676 6556
rect 96380 6502 96406 6554
rect 96406 6502 96436 6554
rect 96460 6502 96470 6554
rect 96470 6502 96516 6554
rect 96540 6502 96586 6554
rect 96586 6502 96596 6554
rect 96620 6502 96650 6554
rect 96650 6502 96676 6554
rect 96380 6500 96436 6502
rect 96460 6500 96516 6502
rect 96540 6500 96596 6502
rect 96620 6500 96676 6502
rect 96380 5466 96436 5468
rect 96460 5466 96516 5468
rect 96540 5466 96596 5468
rect 96620 5466 96676 5468
rect 96380 5414 96406 5466
rect 96406 5414 96436 5466
rect 96460 5414 96470 5466
rect 96470 5414 96516 5466
rect 96540 5414 96586 5466
rect 96586 5414 96596 5466
rect 96620 5414 96650 5466
rect 96650 5414 96676 5466
rect 96380 5412 96436 5414
rect 96460 5412 96516 5414
rect 96540 5412 96596 5414
rect 96620 5412 96676 5414
rect 96380 4378 96436 4380
rect 96460 4378 96516 4380
rect 96540 4378 96596 4380
rect 96620 4378 96676 4380
rect 96380 4326 96406 4378
rect 96406 4326 96436 4378
rect 96460 4326 96470 4378
rect 96470 4326 96516 4378
rect 96540 4326 96586 4378
rect 96586 4326 96596 4378
rect 96620 4326 96650 4378
rect 96650 4326 96676 4378
rect 96380 4324 96436 4326
rect 96460 4324 96516 4326
rect 96540 4324 96596 4326
rect 96620 4324 96676 4326
rect 95054 4256 95110 4312
rect 94686 2488 94742 2544
rect 95606 3612 95608 3632
rect 95608 3612 95660 3632
rect 95660 3612 95662 3632
rect 95606 3576 95662 3612
rect 95146 2624 95202 2680
rect 96380 3290 96436 3292
rect 96460 3290 96516 3292
rect 96540 3290 96596 3292
rect 96620 3290 96676 3292
rect 96380 3238 96406 3290
rect 96406 3238 96436 3290
rect 96460 3238 96470 3290
rect 96470 3238 96516 3290
rect 96540 3238 96586 3290
rect 96586 3238 96596 3290
rect 96620 3238 96650 3290
rect 96650 3238 96676 3290
rect 96380 3236 96436 3238
rect 96460 3236 96516 3238
rect 96540 3236 96596 3238
rect 96620 3236 96676 3238
rect 96380 2202 96436 2204
rect 96460 2202 96516 2204
rect 96540 2202 96596 2204
rect 96620 2202 96676 2204
rect 96380 2150 96406 2202
rect 96406 2150 96436 2202
rect 96460 2150 96470 2202
rect 96470 2150 96516 2202
rect 96540 2150 96586 2202
rect 96586 2150 96596 2202
rect 96620 2150 96650 2202
rect 96650 2150 96676 2202
rect 96380 2148 96436 2150
rect 96460 2148 96516 2150
rect 96540 2148 96596 2150
rect 96620 2148 96676 2150
rect 97998 3848 98054 3904
rect 127100 14170 127156 14172
rect 127180 14170 127236 14172
rect 127260 14170 127316 14172
rect 127340 14170 127396 14172
rect 127100 14118 127126 14170
rect 127126 14118 127156 14170
rect 127180 14118 127190 14170
rect 127190 14118 127236 14170
rect 127260 14118 127306 14170
rect 127306 14118 127316 14170
rect 127340 14118 127370 14170
rect 127370 14118 127396 14170
rect 127100 14116 127156 14118
rect 127180 14116 127236 14118
rect 127260 14116 127316 14118
rect 127340 14116 127396 14118
rect 157820 14170 157876 14172
rect 157900 14170 157956 14172
rect 157980 14170 158036 14172
rect 158060 14170 158116 14172
rect 157820 14118 157846 14170
rect 157846 14118 157876 14170
rect 157900 14118 157910 14170
rect 157910 14118 157956 14170
rect 157980 14118 158026 14170
rect 158026 14118 158036 14170
rect 158060 14118 158090 14170
rect 158090 14118 158116 14170
rect 157820 14116 157876 14118
rect 157900 14116 157956 14118
rect 157980 14116 158036 14118
rect 158060 14116 158116 14118
rect 111740 13626 111796 13628
rect 111820 13626 111876 13628
rect 111900 13626 111956 13628
rect 111980 13626 112036 13628
rect 111740 13574 111766 13626
rect 111766 13574 111796 13626
rect 111820 13574 111830 13626
rect 111830 13574 111876 13626
rect 111900 13574 111946 13626
rect 111946 13574 111956 13626
rect 111980 13574 112010 13626
rect 112010 13574 112036 13626
rect 111740 13572 111796 13574
rect 111820 13572 111876 13574
rect 111900 13572 111956 13574
rect 111980 13572 112036 13574
rect 142460 13626 142516 13628
rect 142540 13626 142596 13628
rect 142620 13626 142676 13628
rect 142700 13626 142756 13628
rect 142460 13574 142486 13626
rect 142486 13574 142516 13626
rect 142540 13574 142550 13626
rect 142550 13574 142596 13626
rect 142620 13574 142666 13626
rect 142666 13574 142676 13626
rect 142700 13574 142730 13626
rect 142730 13574 142756 13626
rect 142460 13572 142516 13574
rect 142540 13572 142596 13574
rect 142620 13572 142676 13574
rect 142700 13572 142756 13574
rect 173180 13626 173236 13628
rect 173260 13626 173316 13628
rect 173340 13626 173396 13628
rect 173420 13626 173476 13628
rect 173180 13574 173206 13626
rect 173206 13574 173236 13626
rect 173260 13574 173270 13626
rect 173270 13574 173316 13626
rect 173340 13574 173386 13626
rect 173386 13574 173396 13626
rect 173420 13574 173450 13626
rect 173450 13574 173476 13626
rect 173180 13572 173236 13574
rect 173260 13572 173316 13574
rect 173340 13572 173396 13574
rect 173420 13572 173476 13574
rect 127100 13082 127156 13084
rect 127180 13082 127236 13084
rect 127260 13082 127316 13084
rect 127340 13082 127396 13084
rect 127100 13030 127126 13082
rect 127126 13030 127156 13082
rect 127180 13030 127190 13082
rect 127190 13030 127236 13082
rect 127260 13030 127306 13082
rect 127306 13030 127316 13082
rect 127340 13030 127370 13082
rect 127370 13030 127396 13082
rect 127100 13028 127156 13030
rect 127180 13028 127236 13030
rect 127260 13028 127316 13030
rect 127340 13028 127396 13030
rect 157820 13082 157876 13084
rect 157900 13082 157956 13084
rect 157980 13082 158036 13084
rect 158060 13082 158116 13084
rect 157820 13030 157846 13082
rect 157846 13030 157876 13082
rect 157900 13030 157910 13082
rect 157910 13030 157956 13082
rect 157980 13030 158026 13082
rect 158026 13030 158036 13082
rect 158060 13030 158090 13082
rect 158090 13030 158116 13082
rect 157820 13028 157876 13030
rect 157900 13028 157956 13030
rect 157980 13028 158036 13030
rect 158060 13028 158116 13030
rect 111740 12538 111796 12540
rect 111820 12538 111876 12540
rect 111900 12538 111956 12540
rect 111980 12538 112036 12540
rect 111740 12486 111766 12538
rect 111766 12486 111796 12538
rect 111820 12486 111830 12538
rect 111830 12486 111876 12538
rect 111900 12486 111946 12538
rect 111946 12486 111956 12538
rect 111980 12486 112010 12538
rect 112010 12486 112036 12538
rect 111740 12484 111796 12486
rect 111820 12484 111876 12486
rect 111900 12484 111956 12486
rect 111980 12484 112036 12486
rect 142460 12538 142516 12540
rect 142540 12538 142596 12540
rect 142620 12538 142676 12540
rect 142700 12538 142756 12540
rect 142460 12486 142486 12538
rect 142486 12486 142516 12538
rect 142540 12486 142550 12538
rect 142550 12486 142596 12538
rect 142620 12486 142666 12538
rect 142666 12486 142676 12538
rect 142700 12486 142730 12538
rect 142730 12486 142756 12538
rect 142460 12484 142516 12486
rect 142540 12484 142596 12486
rect 142620 12484 142676 12486
rect 142700 12484 142756 12486
rect 173180 12538 173236 12540
rect 173260 12538 173316 12540
rect 173340 12538 173396 12540
rect 173420 12538 173476 12540
rect 173180 12486 173206 12538
rect 173206 12486 173236 12538
rect 173260 12486 173270 12538
rect 173270 12486 173316 12538
rect 173340 12486 173386 12538
rect 173386 12486 173396 12538
rect 173420 12486 173450 12538
rect 173450 12486 173476 12538
rect 173180 12484 173236 12486
rect 173260 12484 173316 12486
rect 173340 12484 173396 12486
rect 173420 12484 173476 12486
rect 127100 11994 127156 11996
rect 127180 11994 127236 11996
rect 127260 11994 127316 11996
rect 127340 11994 127396 11996
rect 127100 11942 127126 11994
rect 127126 11942 127156 11994
rect 127180 11942 127190 11994
rect 127190 11942 127236 11994
rect 127260 11942 127306 11994
rect 127306 11942 127316 11994
rect 127340 11942 127370 11994
rect 127370 11942 127396 11994
rect 127100 11940 127156 11942
rect 127180 11940 127236 11942
rect 127260 11940 127316 11942
rect 127340 11940 127396 11942
rect 157820 11994 157876 11996
rect 157900 11994 157956 11996
rect 157980 11994 158036 11996
rect 158060 11994 158116 11996
rect 157820 11942 157846 11994
rect 157846 11942 157876 11994
rect 157900 11942 157910 11994
rect 157910 11942 157956 11994
rect 157980 11942 158026 11994
rect 158026 11942 158036 11994
rect 158060 11942 158090 11994
rect 158090 11942 158116 11994
rect 157820 11940 157876 11942
rect 157900 11940 157956 11942
rect 157980 11940 158036 11942
rect 158060 11940 158116 11942
rect 111740 11450 111796 11452
rect 111820 11450 111876 11452
rect 111900 11450 111956 11452
rect 111980 11450 112036 11452
rect 111740 11398 111766 11450
rect 111766 11398 111796 11450
rect 111820 11398 111830 11450
rect 111830 11398 111876 11450
rect 111900 11398 111946 11450
rect 111946 11398 111956 11450
rect 111980 11398 112010 11450
rect 112010 11398 112036 11450
rect 111740 11396 111796 11398
rect 111820 11396 111876 11398
rect 111900 11396 111956 11398
rect 111980 11396 112036 11398
rect 142460 11450 142516 11452
rect 142540 11450 142596 11452
rect 142620 11450 142676 11452
rect 142700 11450 142756 11452
rect 142460 11398 142486 11450
rect 142486 11398 142516 11450
rect 142540 11398 142550 11450
rect 142550 11398 142596 11450
rect 142620 11398 142666 11450
rect 142666 11398 142676 11450
rect 142700 11398 142730 11450
rect 142730 11398 142756 11450
rect 142460 11396 142516 11398
rect 142540 11396 142596 11398
rect 142620 11396 142676 11398
rect 142700 11396 142756 11398
rect 173180 11450 173236 11452
rect 173260 11450 173316 11452
rect 173340 11450 173396 11452
rect 173420 11450 173476 11452
rect 173180 11398 173206 11450
rect 173206 11398 173236 11450
rect 173260 11398 173270 11450
rect 173270 11398 173316 11450
rect 173340 11398 173386 11450
rect 173386 11398 173396 11450
rect 173420 11398 173450 11450
rect 173450 11398 173476 11450
rect 173180 11396 173236 11398
rect 173260 11396 173316 11398
rect 173340 11396 173396 11398
rect 173420 11396 173476 11398
rect 127100 10906 127156 10908
rect 127180 10906 127236 10908
rect 127260 10906 127316 10908
rect 127340 10906 127396 10908
rect 127100 10854 127126 10906
rect 127126 10854 127156 10906
rect 127180 10854 127190 10906
rect 127190 10854 127236 10906
rect 127260 10854 127306 10906
rect 127306 10854 127316 10906
rect 127340 10854 127370 10906
rect 127370 10854 127396 10906
rect 127100 10852 127156 10854
rect 127180 10852 127236 10854
rect 127260 10852 127316 10854
rect 127340 10852 127396 10854
rect 157820 10906 157876 10908
rect 157900 10906 157956 10908
rect 157980 10906 158036 10908
rect 158060 10906 158116 10908
rect 157820 10854 157846 10906
rect 157846 10854 157876 10906
rect 157900 10854 157910 10906
rect 157910 10854 157956 10906
rect 157980 10854 158026 10906
rect 158026 10854 158036 10906
rect 158060 10854 158090 10906
rect 158090 10854 158116 10906
rect 157820 10852 157876 10854
rect 157900 10852 157956 10854
rect 157980 10852 158036 10854
rect 158060 10852 158116 10854
rect 111740 10362 111796 10364
rect 111820 10362 111876 10364
rect 111900 10362 111956 10364
rect 111980 10362 112036 10364
rect 111740 10310 111766 10362
rect 111766 10310 111796 10362
rect 111820 10310 111830 10362
rect 111830 10310 111876 10362
rect 111900 10310 111946 10362
rect 111946 10310 111956 10362
rect 111980 10310 112010 10362
rect 112010 10310 112036 10362
rect 111740 10308 111796 10310
rect 111820 10308 111876 10310
rect 111900 10308 111956 10310
rect 111980 10308 112036 10310
rect 142460 10362 142516 10364
rect 142540 10362 142596 10364
rect 142620 10362 142676 10364
rect 142700 10362 142756 10364
rect 142460 10310 142486 10362
rect 142486 10310 142516 10362
rect 142540 10310 142550 10362
rect 142550 10310 142596 10362
rect 142620 10310 142666 10362
rect 142666 10310 142676 10362
rect 142700 10310 142730 10362
rect 142730 10310 142756 10362
rect 142460 10308 142516 10310
rect 142540 10308 142596 10310
rect 142620 10308 142676 10310
rect 142700 10308 142756 10310
rect 173180 10362 173236 10364
rect 173260 10362 173316 10364
rect 173340 10362 173396 10364
rect 173420 10362 173476 10364
rect 173180 10310 173206 10362
rect 173206 10310 173236 10362
rect 173260 10310 173270 10362
rect 173270 10310 173316 10362
rect 173340 10310 173386 10362
rect 173386 10310 173396 10362
rect 173420 10310 173450 10362
rect 173450 10310 173476 10362
rect 173180 10308 173236 10310
rect 173260 10308 173316 10310
rect 173340 10308 173396 10310
rect 173420 10308 173476 10310
rect 127100 9818 127156 9820
rect 127180 9818 127236 9820
rect 127260 9818 127316 9820
rect 127340 9818 127396 9820
rect 127100 9766 127126 9818
rect 127126 9766 127156 9818
rect 127180 9766 127190 9818
rect 127190 9766 127236 9818
rect 127260 9766 127306 9818
rect 127306 9766 127316 9818
rect 127340 9766 127370 9818
rect 127370 9766 127396 9818
rect 127100 9764 127156 9766
rect 127180 9764 127236 9766
rect 127260 9764 127316 9766
rect 127340 9764 127396 9766
rect 157820 9818 157876 9820
rect 157900 9818 157956 9820
rect 157980 9818 158036 9820
rect 158060 9818 158116 9820
rect 157820 9766 157846 9818
rect 157846 9766 157876 9818
rect 157900 9766 157910 9818
rect 157910 9766 157956 9818
rect 157980 9766 158026 9818
rect 158026 9766 158036 9818
rect 158060 9766 158090 9818
rect 158090 9766 158116 9818
rect 157820 9764 157876 9766
rect 157900 9764 157956 9766
rect 157980 9764 158036 9766
rect 158060 9764 158116 9766
rect 111740 9274 111796 9276
rect 111820 9274 111876 9276
rect 111900 9274 111956 9276
rect 111980 9274 112036 9276
rect 111740 9222 111766 9274
rect 111766 9222 111796 9274
rect 111820 9222 111830 9274
rect 111830 9222 111876 9274
rect 111900 9222 111946 9274
rect 111946 9222 111956 9274
rect 111980 9222 112010 9274
rect 112010 9222 112036 9274
rect 111740 9220 111796 9222
rect 111820 9220 111876 9222
rect 111900 9220 111956 9222
rect 111980 9220 112036 9222
rect 142460 9274 142516 9276
rect 142540 9274 142596 9276
rect 142620 9274 142676 9276
rect 142700 9274 142756 9276
rect 142460 9222 142486 9274
rect 142486 9222 142516 9274
rect 142540 9222 142550 9274
rect 142550 9222 142596 9274
rect 142620 9222 142666 9274
rect 142666 9222 142676 9274
rect 142700 9222 142730 9274
rect 142730 9222 142756 9274
rect 142460 9220 142516 9222
rect 142540 9220 142596 9222
rect 142620 9220 142676 9222
rect 142700 9220 142756 9222
rect 173180 9274 173236 9276
rect 173260 9274 173316 9276
rect 173340 9274 173396 9276
rect 173420 9274 173476 9276
rect 173180 9222 173206 9274
rect 173206 9222 173236 9274
rect 173260 9222 173270 9274
rect 173270 9222 173316 9274
rect 173340 9222 173386 9274
rect 173386 9222 173396 9274
rect 173420 9222 173450 9274
rect 173450 9222 173476 9274
rect 173180 9220 173236 9222
rect 173260 9220 173316 9222
rect 173340 9220 173396 9222
rect 173420 9220 173476 9222
rect 127100 8730 127156 8732
rect 127180 8730 127236 8732
rect 127260 8730 127316 8732
rect 127340 8730 127396 8732
rect 127100 8678 127126 8730
rect 127126 8678 127156 8730
rect 127180 8678 127190 8730
rect 127190 8678 127236 8730
rect 127260 8678 127306 8730
rect 127306 8678 127316 8730
rect 127340 8678 127370 8730
rect 127370 8678 127396 8730
rect 127100 8676 127156 8678
rect 127180 8676 127236 8678
rect 127260 8676 127316 8678
rect 127340 8676 127396 8678
rect 157820 8730 157876 8732
rect 157900 8730 157956 8732
rect 157980 8730 158036 8732
rect 158060 8730 158116 8732
rect 157820 8678 157846 8730
rect 157846 8678 157876 8730
rect 157900 8678 157910 8730
rect 157910 8678 157956 8730
rect 157980 8678 158026 8730
rect 158026 8678 158036 8730
rect 158060 8678 158090 8730
rect 158090 8678 158116 8730
rect 157820 8676 157876 8678
rect 157900 8676 157956 8678
rect 157980 8676 158036 8678
rect 158060 8676 158116 8678
rect 111740 8186 111796 8188
rect 111820 8186 111876 8188
rect 111900 8186 111956 8188
rect 111980 8186 112036 8188
rect 111740 8134 111766 8186
rect 111766 8134 111796 8186
rect 111820 8134 111830 8186
rect 111830 8134 111876 8186
rect 111900 8134 111946 8186
rect 111946 8134 111956 8186
rect 111980 8134 112010 8186
rect 112010 8134 112036 8186
rect 111740 8132 111796 8134
rect 111820 8132 111876 8134
rect 111900 8132 111956 8134
rect 111980 8132 112036 8134
rect 142460 8186 142516 8188
rect 142540 8186 142596 8188
rect 142620 8186 142676 8188
rect 142700 8186 142756 8188
rect 142460 8134 142486 8186
rect 142486 8134 142516 8186
rect 142540 8134 142550 8186
rect 142550 8134 142596 8186
rect 142620 8134 142666 8186
rect 142666 8134 142676 8186
rect 142700 8134 142730 8186
rect 142730 8134 142756 8186
rect 142460 8132 142516 8134
rect 142540 8132 142596 8134
rect 142620 8132 142676 8134
rect 142700 8132 142756 8134
rect 173180 8186 173236 8188
rect 173260 8186 173316 8188
rect 173340 8186 173396 8188
rect 173420 8186 173476 8188
rect 173180 8134 173206 8186
rect 173206 8134 173236 8186
rect 173260 8134 173270 8186
rect 173270 8134 173316 8186
rect 173340 8134 173386 8186
rect 173386 8134 173396 8186
rect 173420 8134 173450 8186
rect 173450 8134 173476 8186
rect 173180 8132 173236 8134
rect 173260 8132 173316 8134
rect 173340 8132 173396 8134
rect 173420 8132 173476 8134
rect 127100 7642 127156 7644
rect 127180 7642 127236 7644
rect 127260 7642 127316 7644
rect 127340 7642 127396 7644
rect 127100 7590 127126 7642
rect 127126 7590 127156 7642
rect 127180 7590 127190 7642
rect 127190 7590 127236 7642
rect 127260 7590 127306 7642
rect 127306 7590 127316 7642
rect 127340 7590 127370 7642
rect 127370 7590 127396 7642
rect 127100 7588 127156 7590
rect 127180 7588 127236 7590
rect 127260 7588 127316 7590
rect 127340 7588 127396 7590
rect 157820 7642 157876 7644
rect 157900 7642 157956 7644
rect 157980 7642 158036 7644
rect 158060 7642 158116 7644
rect 157820 7590 157846 7642
rect 157846 7590 157876 7642
rect 157900 7590 157910 7642
rect 157910 7590 157956 7642
rect 157980 7590 158026 7642
rect 158026 7590 158036 7642
rect 158060 7590 158090 7642
rect 158090 7590 158116 7642
rect 157820 7588 157876 7590
rect 157900 7588 157956 7590
rect 157980 7588 158036 7590
rect 158060 7588 158116 7590
rect 111740 7098 111796 7100
rect 111820 7098 111876 7100
rect 111900 7098 111956 7100
rect 111980 7098 112036 7100
rect 111740 7046 111766 7098
rect 111766 7046 111796 7098
rect 111820 7046 111830 7098
rect 111830 7046 111876 7098
rect 111900 7046 111946 7098
rect 111946 7046 111956 7098
rect 111980 7046 112010 7098
rect 112010 7046 112036 7098
rect 111740 7044 111796 7046
rect 111820 7044 111876 7046
rect 111900 7044 111956 7046
rect 111980 7044 112036 7046
rect 142460 7098 142516 7100
rect 142540 7098 142596 7100
rect 142620 7098 142676 7100
rect 142700 7098 142756 7100
rect 142460 7046 142486 7098
rect 142486 7046 142516 7098
rect 142540 7046 142550 7098
rect 142550 7046 142596 7098
rect 142620 7046 142666 7098
rect 142666 7046 142676 7098
rect 142700 7046 142730 7098
rect 142730 7046 142756 7098
rect 142460 7044 142516 7046
rect 142540 7044 142596 7046
rect 142620 7044 142676 7046
rect 142700 7044 142756 7046
rect 173180 7098 173236 7100
rect 173260 7098 173316 7100
rect 173340 7098 173396 7100
rect 173420 7098 173476 7100
rect 173180 7046 173206 7098
rect 173206 7046 173236 7098
rect 173260 7046 173270 7098
rect 173270 7046 173316 7098
rect 173340 7046 173386 7098
rect 173386 7046 173396 7098
rect 173420 7046 173450 7098
rect 173450 7046 173476 7098
rect 173180 7044 173236 7046
rect 173260 7044 173316 7046
rect 173340 7044 173396 7046
rect 173420 7044 173476 7046
rect 127100 6554 127156 6556
rect 127180 6554 127236 6556
rect 127260 6554 127316 6556
rect 127340 6554 127396 6556
rect 127100 6502 127126 6554
rect 127126 6502 127156 6554
rect 127180 6502 127190 6554
rect 127190 6502 127236 6554
rect 127260 6502 127306 6554
rect 127306 6502 127316 6554
rect 127340 6502 127370 6554
rect 127370 6502 127396 6554
rect 127100 6500 127156 6502
rect 127180 6500 127236 6502
rect 127260 6500 127316 6502
rect 127340 6500 127396 6502
rect 157820 6554 157876 6556
rect 157900 6554 157956 6556
rect 157980 6554 158036 6556
rect 158060 6554 158116 6556
rect 157820 6502 157846 6554
rect 157846 6502 157876 6554
rect 157900 6502 157910 6554
rect 157910 6502 157956 6554
rect 157980 6502 158026 6554
rect 158026 6502 158036 6554
rect 158060 6502 158090 6554
rect 158090 6502 158116 6554
rect 157820 6500 157876 6502
rect 157900 6500 157956 6502
rect 157980 6500 158036 6502
rect 158060 6500 158116 6502
rect 111740 6010 111796 6012
rect 111820 6010 111876 6012
rect 111900 6010 111956 6012
rect 111980 6010 112036 6012
rect 111740 5958 111766 6010
rect 111766 5958 111796 6010
rect 111820 5958 111830 6010
rect 111830 5958 111876 6010
rect 111900 5958 111946 6010
rect 111946 5958 111956 6010
rect 111980 5958 112010 6010
rect 112010 5958 112036 6010
rect 111740 5956 111796 5958
rect 111820 5956 111876 5958
rect 111900 5956 111956 5958
rect 111980 5956 112036 5958
rect 142460 6010 142516 6012
rect 142540 6010 142596 6012
rect 142620 6010 142676 6012
rect 142700 6010 142756 6012
rect 142460 5958 142486 6010
rect 142486 5958 142516 6010
rect 142540 5958 142550 6010
rect 142550 5958 142596 6010
rect 142620 5958 142666 6010
rect 142666 5958 142676 6010
rect 142700 5958 142730 6010
rect 142730 5958 142756 6010
rect 142460 5956 142516 5958
rect 142540 5956 142596 5958
rect 142620 5956 142676 5958
rect 142700 5956 142756 5958
rect 173180 6010 173236 6012
rect 173260 6010 173316 6012
rect 173340 6010 173396 6012
rect 173420 6010 173476 6012
rect 173180 5958 173206 6010
rect 173206 5958 173236 6010
rect 173260 5958 173270 6010
rect 173270 5958 173316 6010
rect 173340 5958 173386 6010
rect 173386 5958 173396 6010
rect 173420 5958 173450 6010
rect 173450 5958 173476 6010
rect 173180 5956 173236 5958
rect 173260 5956 173316 5958
rect 173340 5956 173396 5958
rect 173420 5956 173476 5958
rect 127100 5466 127156 5468
rect 127180 5466 127236 5468
rect 127260 5466 127316 5468
rect 127340 5466 127396 5468
rect 127100 5414 127126 5466
rect 127126 5414 127156 5466
rect 127180 5414 127190 5466
rect 127190 5414 127236 5466
rect 127260 5414 127306 5466
rect 127306 5414 127316 5466
rect 127340 5414 127370 5466
rect 127370 5414 127396 5466
rect 127100 5412 127156 5414
rect 127180 5412 127236 5414
rect 127260 5412 127316 5414
rect 127340 5412 127396 5414
rect 157820 5466 157876 5468
rect 157900 5466 157956 5468
rect 157980 5466 158036 5468
rect 158060 5466 158116 5468
rect 157820 5414 157846 5466
rect 157846 5414 157876 5466
rect 157900 5414 157910 5466
rect 157910 5414 157956 5466
rect 157980 5414 158026 5466
rect 158026 5414 158036 5466
rect 158060 5414 158090 5466
rect 158090 5414 158116 5466
rect 157820 5412 157876 5414
rect 157900 5412 157956 5414
rect 157980 5412 158036 5414
rect 158060 5412 158116 5414
rect 111740 4922 111796 4924
rect 111820 4922 111876 4924
rect 111900 4922 111956 4924
rect 111980 4922 112036 4924
rect 111740 4870 111766 4922
rect 111766 4870 111796 4922
rect 111820 4870 111830 4922
rect 111830 4870 111876 4922
rect 111900 4870 111946 4922
rect 111946 4870 111956 4922
rect 111980 4870 112010 4922
rect 112010 4870 112036 4922
rect 111740 4868 111796 4870
rect 111820 4868 111876 4870
rect 111900 4868 111956 4870
rect 111980 4868 112036 4870
rect 142460 4922 142516 4924
rect 142540 4922 142596 4924
rect 142620 4922 142676 4924
rect 142700 4922 142756 4924
rect 142460 4870 142486 4922
rect 142486 4870 142516 4922
rect 142540 4870 142550 4922
rect 142550 4870 142596 4922
rect 142620 4870 142666 4922
rect 142666 4870 142676 4922
rect 142700 4870 142730 4922
rect 142730 4870 142756 4922
rect 142460 4868 142516 4870
rect 142540 4868 142596 4870
rect 142620 4868 142676 4870
rect 142700 4868 142756 4870
rect 173180 4922 173236 4924
rect 173260 4922 173316 4924
rect 173340 4922 173396 4924
rect 173420 4922 173476 4924
rect 173180 4870 173206 4922
rect 173206 4870 173236 4922
rect 173260 4870 173270 4922
rect 173270 4870 173316 4922
rect 173340 4870 173386 4922
rect 173386 4870 173396 4922
rect 173420 4870 173450 4922
rect 173450 4870 173476 4922
rect 173180 4868 173236 4870
rect 173260 4868 173316 4870
rect 173340 4868 173396 4870
rect 173420 4868 173476 4870
rect 101034 2760 101090 2816
rect 101402 2896 101458 2952
rect 101586 3984 101642 4040
rect 101862 3712 101918 3768
rect 101770 3576 101826 3632
rect 102138 3052 102194 3088
rect 102138 3032 102140 3052
rect 102140 3032 102192 3052
rect 102192 3032 102194 3052
rect 127100 4378 127156 4380
rect 127180 4378 127236 4380
rect 127260 4378 127316 4380
rect 127340 4378 127396 4380
rect 127100 4326 127126 4378
rect 127126 4326 127156 4378
rect 127180 4326 127190 4378
rect 127190 4326 127236 4378
rect 127260 4326 127306 4378
rect 127306 4326 127316 4378
rect 127340 4326 127370 4378
rect 127370 4326 127396 4378
rect 127100 4324 127156 4326
rect 127180 4324 127236 4326
rect 127260 4324 127316 4326
rect 127340 4324 127396 4326
rect 157820 4378 157876 4380
rect 157900 4378 157956 4380
rect 157980 4378 158036 4380
rect 158060 4378 158116 4380
rect 157820 4326 157846 4378
rect 157846 4326 157876 4378
rect 157900 4326 157910 4378
rect 157910 4326 157956 4378
rect 157980 4326 158026 4378
rect 158026 4326 158036 4378
rect 158060 4326 158090 4378
rect 158090 4326 158116 4378
rect 157820 4324 157876 4326
rect 157900 4324 157956 4326
rect 157980 4324 158036 4326
rect 158060 4324 158116 4326
rect 102874 2916 102930 2952
rect 102874 2896 102876 2916
rect 102876 2896 102928 2916
rect 102928 2896 102930 2916
rect 103518 3168 103574 3224
rect 111740 3834 111796 3836
rect 111820 3834 111876 3836
rect 111900 3834 111956 3836
rect 111980 3834 112036 3836
rect 111740 3782 111766 3834
rect 111766 3782 111796 3834
rect 111820 3782 111830 3834
rect 111830 3782 111876 3834
rect 111900 3782 111946 3834
rect 111946 3782 111956 3834
rect 111980 3782 112010 3834
rect 112010 3782 112036 3834
rect 111740 3780 111796 3782
rect 111820 3780 111876 3782
rect 111900 3780 111956 3782
rect 111980 3780 112036 3782
rect 111740 2746 111796 2748
rect 111820 2746 111876 2748
rect 111900 2746 111956 2748
rect 111980 2746 112036 2748
rect 111740 2694 111766 2746
rect 111766 2694 111796 2746
rect 111820 2694 111830 2746
rect 111830 2694 111876 2746
rect 111900 2694 111946 2746
rect 111946 2694 111956 2746
rect 111980 2694 112010 2746
rect 112010 2694 112036 2746
rect 111740 2692 111796 2694
rect 111820 2692 111876 2694
rect 111900 2692 111956 2694
rect 111980 2692 112036 2694
rect 127100 3290 127156 3292
rect 127180 3290 127236 3292
rect 127260 3290 127316 3292
rect 127340 3290 127396 3292
rect 127100 3238 127126 3290
rect 127126 3238 127156 3290
rect 127180 3238 127190 3290
rect 127190 3238 127236 3290
rect 127260 3238 127306 3290
rect 127306 3238 127316 3290
rect 127340 3238 127370 3290
rect 127370 3238 127396 3290
rect 127100 3236 127156 3238
rect 127180 3236 127236 3238
rect 127260 3236 127316 3238
rect 127340 3236 127396 3238
rect 127100 2202 127156 2204
rect 127180 2202 127236 2204
rect 127260 2202 127316 2204
rect 127340 2202 127396 2204
rect 127100 2150 127126 2202
rect 127126 2150 127156 2202
rect 127180 2150 127190 2202
rect 127190 2150 127236 2202
rect 127260 2150 127306 2202
rect 127306 2150 127316 2202
rect 127340 2150 127370 2202
rect 127370 2150 127396 2202
rect 127100 2148 127156 2150
rect 127180 2148 127236 2150
rect 127260 2148 127316 2150
rect 127340 2148 127396 2150
rect 142460 3834 142516 3836
rect 142540 3834 142596 3836
rect 142620 3834 142676 3836
rect 142700 3834 142756 3836
rect 142460 3782 142486 3834
rect 142486 3782 142516 3834
rect 142540 3782 142550 3834
rect 142550 3782 142596 3834
rect 142620 3782 142666 3834
rect 142666 3782 142676 3834
rect 142700 3782 142730 3834
rect 142730 3782 142756 3834
rect 142460 3780 142516 3782
rect 142540 3780 142596 3782
rect 142620 3780 142676 3782
rect 142700 3780 142756 3782
rect 142460 2746 142516 2748
rect 142540 2746 142596 2748
rect 142620 2746 142676 2748
rect 142700 2746 142756 2748
rect 142460 2694 142486 2746
rect 142486 2694 142516 2746
rect 142540 2694 142550 2746
rect 142550 2694 142596 2746
rect 142620 2694 142666 2746
rect 142666 2694 142676 2746
rect 142700 2694 142730 2746
rect 142730 2694 142756 2746
rect 142460 2692 142516 2694
rect 142540 2692 142596 2694
rect 142620 2692 142676 2694
rect 142700 2692 142756 2694
rect 157820 3290 157876 3292
rect 157900 3290 157956 3292
rect 157980 3290 158036 3292
rect 158060 3290 158116 3292
rect 157820 3238 157846 3290
rect 157846 3238 157876 3290
rect 157900 3238 157910 3290
rect 157910 3238 157956 3290
rect 157980 3238 158026 3290
rect 158026 3238 158036 3290
rect 158060 3238 158090 3290
rect 158090 3238 158116 3290
rect 157820 3236 157876 3238
rect 157900 3236 157956 3238
rect 157980 3236 158036 3238
rect 158060 3236 158116 3238
rect 157820 2202 157876 2204
rect 157900 2202 157956 2204
rect 157980 2202 158036 2204
rect 158060 2202 158116 2204
rect 157820 2150 157846 2202
rect 157846 2150 157876 2202
rect 157900 2150 157910 2202
rect 157910 2150 157956 2202
rect 157980 2150 158026 2202
rect 158026 2150 158036 2202
rect 158060 2150 158090 2202
rect 158090 2150 158116 2202
rect 157820 2148 157876 2150
rect 157900 2148 157956 2150
rect 157980 2148 158036 2150
rect 158060 2148 158116 2150
rect 173180 3834 173236 3836
rect 173260 3834 173316 3836
rect 173340 3834 173396 3836
rect 173420 3834 173476 3836
rect 173180 3782 173206 3834
rect 173206 3782 173236 3834
rect 173260 3782 173270 3834
rect 173270 3782 173316 3834
rect 173340 3782 173386 3834
rect 173386 3782 173396 3834
rect 173420 3782 173450 3834
rect 173450 3782 173476 3834
rect 173180 3780 173236 3782
rect 173260 3780 173316 3782
rect 173340 3780 173396 3782
rect 173420 3780 173476 3782
rect 173180 2746 173236 2748
rect 173260 2746 173316 2748
rect 173340 2746 173396 2748
rect 173420 2746 173476 2748
rect 173180 2694 173206 2746
rect 173206 2694 173236 2746
rect 173260 2694 173270 2746
rect 173270 2694 173316 2746
rect 173340 2694 173386 2746
rect 173386 2694 173396 2746
rect 173420 2694 173450 2746
rect 173450 2694 173476 2746
rect 173180 2692 173236 2694
rect 173260 2692 173316 2694
rect 173340 2692 173396 2694
rect 173420 2692 173476 2694
<< metal3 >>
rect 4208 117536 4528 117537
rect 4208 117472 4216 117536
rect 4280 117472 4296 117536
rect 4360 117472 4376 117536
rect 4440 117472 4456 117536
rect 4520 117472 4528 117536
rect 4208 117471 4528 117472
rect 34928 117536 35248 117537
rect 34928 117472 34936 117536
rect 35000 117472 35016 117536
rect 35080 117472 35096 117536
rect 35160 117472 35176 117536
rect 35240 117472 35248 117536
rect 34928 117471 35248 117472
rect 65648 117536 65968 117537
rect 65648 117472 65656 117536
rect 65720 117472 65736 117536
rect 65800 117472 65816 117536
rect 65880 117472 65896 117536
rect 65960 117472 65968 117536
rect 65648 117471 65968 117472
rect 96368 117536 96688 117537
rect 96368 117472 96376 117536
rect 96440 117472 96456 117536
rect 96520 117472 96536 117536
rect 96600 117472 96616 117536
rect 96680 117472 96688 117536
rect 96368 117471 96688 117472
rect 127088 117536 127408 117537
rect 127088 117472 127096 117536
rect 127160 117472 127176 117536
rect 127240 117472 127256 117536
rect 127320 117472 127336 117536
rect 127400 117472 127408 117536
rect 127088 117471 127408 117472
rect 157808 117536 158128 117537
rect 157808 117472 157816 117536
rect 157880 117472 157896 117536
rect 157960 117472 157976 117536
rect 158040 117472 158056 117536
rect 158120 117472 158128 117536
rect 157808 117471 158128 117472
rect 19568 116992 19888 116993
rect 19568 116928 19576 116992
rect 19640 116928 19656 116992
rect 19720 116928 19736 116992
rect 19800 116928 19816 116992
rect 19880 116928 19888 116992
rect 19568 116927 19888 116928
rect 50288 116992 50608 116993
rect 50288 116928 50296 116992
rect 50360 116928 50376 116992
rect 50440 116928 50456 116992
rect 50520 116928 50536 116992
rect 50600 116928 50608 116992
rect 50288 116927 50608 116928
rect 81008 116992 81328 116993
rect 81008 116928 81016 116992
rect 81080 116928 81096 116992
rect 81160 116928 81176 116992
rect 81240 116928 81256 116992
rect 81320 116928 81328 116992
rect 81008 116927 81328 116928
rect 111728 116992 112048 116993
rect 111728 116928 111736 116992
rect 111800 116928 111816 116992
rect 111880 116928 111896 116992
rect 111960 116928 111976 116992
rect 112040 116928 112048 116992
rect 111728 116927 112048 116928
rect 142448 116992 142768 116993
rect 142448 116928 142456 116992
rect 142520 116928 142536 116992
rect 142600 116928 142616 116992
rect 142680 116928 142696 116992
rect 142760 116928 142768 116992
rect 142448 116927 142768 116928
rect 173168 116992 173488 116993
rect 173168 116928 173176 116992
rect 173240 116928 173256 116992
rect 173320 116928 173336 116992
rect 173400 116928 173416 116992
rect 173480 116928 173488 116992
rect 173168 116927 173488 116928
rect 4208 116448 4528 116449
rect 4208 116384 4216 116448
rect 4280 116384 4296 116448
rect 4360 116384 4376 116448
rect 4440 116384 4456 116448
rect 4520 116384 4528 116448
rect 4208 116383 4528 116384
rect 34928 116448 35248 116449
rect 34928 116384 34936 116448
rect 35000 116384 35016 116448
rect 35080 116384 35096 116448
rect 35160 116384 35176 116448
rect 35240 116384 35248 116448
rect 34928 116383 35248 116384
rect 65648 116448 65968 116449
rect 65648 116384 65656 116448
rect 65720 116384 65736 116448
rect 65800 116384 65816 116448
rect 65880 116384 65896 116448
rect 65960 116384 65968 116448
rect 65648 116383 65968 116384
rect 96368 116448 96688 116449
rect 96368 116384 96376 116448
rect 96440 116384 96456 116448
rect 96520 116384 96536 116448
rect 96600 116384 96616 116448
rect 96680 116384 96688 116448
rect 96368 116383 96688 116384
rect 127088 116448 127408 116449
rect 127088 116384 127096 116448
rect 127160 116384 127176 116448
rect 127240 116384 127256 116448
rect 127320 116384 127336 116448
rect 127400 116384 127408 116448
rect 127088 116383 127408 116384
rect 157808 116448 158128 116449
rect 157808 116384 157816 116448
rect 157880 116384 157896 116448
rect 157960 116384 157976 116448
rect 158040 116384 158056 116448
rect 158120 116384 158128 116448
rect 157808 116383 158128 116384
rect 19568 115904 19888 115905
rect 19568 115840 19576 115904
rect 19640 115840 19656 115904
rect 19720 115840 19736 115904
rect 19800 115840 19816 115904
rect 19880 115840 19888 115904
rect 19568 115839 19888 115840
rect 50288 115904 50608 115905
rect 50288 115840 50296 115904
rect 50360 115840 50376 115904
rect 50440 115840 50456 115904
rect 50520 115840 50536 115904
rect 50600 115840 50608 115904
rect 50288 115839 50608 115840
rect 81008 115904 81328 115905
rect 81008 115840 81016 115904
rect 81080 115840 81096 115904
rect 81160 115840 81176 115904
rect 81240 115840 81256 115904
rect 81320 115840 81328 115904
rect 81008 115839 81328 115840
rect 111728 115904 112048 115905
rect 111728 115840 111736 115904
rect 111800 115840 111816 115904
rect 111880 115840 111896 115904
rect 111960 115840 111976 115904
rect 112040 115840 112048 115904
rect 111728 115839 112048 115840
rect 142448 115904 142768 115905
rect 142448 115840 142456 115904
rect 142520 115840 142536 115904
rect 142600 115840 142616 115904
rect 142680 115840 142696 115904
rect 142760 115840 142768 115904
rect 142448 115839 142768 115840
rect 173168 115904 173488 115905
rect 173168 115840 173176 115904
rect 173240 115840 173256 115904
rect 173320 115840 173336 115904
rect 173400 115840 173416 115904
rect 173480 115840 173488 115904
rect 173168 115839 173488 115840
rect 4208 115360 4528 115361
rect 4208 115296 4216 115360
rect 4280 115296 4296 115360
rect 4360 115296 4376 115360
rect 4440 115296 4456 115360
rect 4520 115296 4528 115360
rect 4208 115295 4528 115296
rect 34928 115360 35248 115361
rect 34928 115296 34936 115360
rect 35000 115296 35016 115360
rect 35080 115296 35096 115360
rect 35160 115296 35176 115360
rect 35240 115296 35248 115360
rect 34928 115295 35248 115296
rect 65648 115360 65968 115361
rect 65648 115296 65656 115360
rect 65720 115296 65736 115360
rect 65800 115296 65816 115360
rect 65880 115296 65896 115360
rect 65960 115296 65968 115360
rect 65648 115295 65968 115296
rect 96368 115360 96688 115361
rect 96368 115296 96376 115360
rect 96440 115296 96456 115360
rect 96520 115296 96536 115360
rect 96600 115296 96616 115360
rect 96680 115296 96688 115360
rect 96368 115295 96688 115296
rect 127088 115360 127408 115361
rect 127088 115296 127096 115360
rect 127160 115296 127176 115360
rect 127240 115296 127256 115360
rect 127320 115296 127336 115360
rect 127400 115296 127408 115360
rect 127088 115295 127408 115296
rect 157808 115360 158128 115361
rect 157808 115296 157816 115360
rect 157880 115296 157896 115360
rect 157960 115296 157976 115360
rect 158040 115296 158056 115360
rect 158120 115296 158128 115360
rect 157808 115295 158128 115296
rect 19568 114816 19888 114817
rect 19568 114752 19576 114816
rect 19640 114752 19656 114816
rect 19720 114752 19736 114816
rect 19800 114752 19816 114816
rect 19880 114752 19888 114816
rect 19568 114751 19888 114752
rect 50288 114816 50608 114817
rect 50288 114752 50296 114816
rect 50360 114752 50376 114816
rect 50440 114752 50456 114816
rect 50520 114752 50536 114816
rect 50600 114752 50608 114816
rect 50288 114751 50608 114752
rect 81008 114816 81328 114817
rect 81008 114752 81016 114816
rect 81080 114752 81096 114816
rect 81160 114752 81176 114816
rect 81240 114752 81256 114816
rect 81320 114752 81328 114816
rect 81008 114751 81328 114752
rect 111728 114816 112048 114817
rect 111728 114752 111736 114816
rect 111800 114752 111816 114816
rect 111880 114752 111896 114816
rect 111960 114752 111976 114816
rect 112040 114752 112048 114816
rect 111728 114751 112048 114752
rect 142448 114816 142768 114817
rect 142448 114752 142456 114816
rect 142520 114752 142536 114816
rect 142600 114752 142616 114816
rect 142680 114752 142696 114816
rect 142760 114752 142768 114816
rect 142448 114751 142768 114752
rect 173168 114816 173488 114817
rect 173168 114752 173176 114816
rect 173240 114752 173256 114816
rect 173320 114752 173336 114816
rect 173400 114752 173416 114816
rect 173480 114752 173488 114816
rect 173168 114751 173488 114752
rect 4208 114272 4528 114273
rect 4208 114208 4216 114272
rect 4280 114208 4296 114272
rect 4360 114208 4376 114272
rect 4440 114208 4456 114272
rect 4520 114208 4528 114272
rect 4208 114207 4528 114208
rect 34928 114272 35248 114273
rect 34928 114208 34936 114272
rect 35000 114208 35016 114272
rect 35080 114208 35096 114272
rect 35160 114208 35176 114272
rect 35240 114208 35248 114272
rect 34928 114207 35248 114208
rect 65648 114272 65968 114273
rect 65648 114208 65656 114272
rect 65720 114208 65736 114272
rect 65800 114208 65816 114272
rect 65880 114208 65896 114272
rect 65960 114208 65968 114272
rect 65648 114207 65968 114208
rect 96368 114272 96688 114273
rect 96368 114208 96376 114272
rect 96440 114208 96456 114272
rect 96520 114208 96536 114272
rect 96600 114208 96616 114272
rect 96680 114208 96688 114272
rect 96368 114207 96688 114208
rect 127088 114272 127408 114273
rect 127088 114208 127096 114272
rect 127160 114208 127176 114272
rect 127240 114208 127256 114272
rect 127320 114208 127336 114272
rect 127400 114208 127408 114272
rect 127088 114207 127408 114208
rect 157808 114272 158128 114273
rect 157808 114208 157816 114272
rect 157880 114208 157896 114272
rect 157960 114208 157976 114272
rect 158040 114208 158056 114272
rect 158120 114208 158128 114272
rect 157808 114207 158128 114208
rect 19568 113728 19888 113729
rect 19568 113664 19576 113728
rect 19640 113664 19656 113728
rect 19720 113664 19736 113728
rect 19800 113664 19816 113728
rect 19880 113664 19888 113728
rect 19568 113663 19888 113664
rect 50288 113728 50608 113729
rect 50288 113664 50296 113728
rect 50360 113664 50376 113728
rect 50440 113664 50456 113728
rect 50520 113664 50536 113728
rect 50600 113664 50608 113728
rect 50288 113663 50608 113664
rect 81008 113728 81328 113729
rect 81008 113664 81016 113728
rect 81080 113664 81096 113728
rect 81160 113664 81176 113728
rect 81240 113664 81256 113728
rect 81320 113664 81328 113728
rect 81008 113663 81328 113664
rect 111728 113728 112048 113729
rect 111728 113664 111736 113728
rect 111800 113664 111816 113728
rect 111880 113664 111896 113728
rect 111960 113664 111976 113728
rect 112040 113664 112048 113728
rect 111728 113663 112048 113664
rect 142448 113728 142768 113729
rect 142448 113664 142456 113728
rect 142520 113664 142536 113728
rect 142600 113664 142616 113728
rect 142680 113664 142696 113728
rect 142760 113664 142768 113728
rect 142448 113663 142768 113664
rect 173168 113728 173488 113729
rect 173168 113664 173176 113728
rect 173240 113664 173256 113728
rect 173320 113664 173336 113728
rect 173400 113664 173416 113728
rect 173480 113664 173488 113728
rect 173168 113663 173488 113664
rect 4208 113184 4528 113185
rect 4208 113120 4216 113184
rect 4280 113120 4296 113184
rect 4360 113120 4376 113184
rect 4440 113120 4456 113184
rect 4520 113120 4528 113184
rect 4208 113119 4528 113120
rect 34928 113184 35248 113185
rect 34928 113120 34936 113184
rect 35000 113120 35016 113184
rect 35080 113120 35096 113184
rect 35160 113120 35176 113184
rect 35240 113120 35248 113184
rect 34928 113119 35248 113120
rect 65648 113184 65968 113185
rect 65648 113120 65656 113184
rect 65720 113120 65736 113184
rect 65800 113120 65816 113184
rect 65880 113120 65896 113184
rect 65960 113120 65968 113184
rect 65648 113119 65968 113120
rect 96368 113184 96688 113185
rect 96368 113120 96376 113184
rect 96440 113120 96456 113184
rect 96520 113120 96536 113184
rect 96600 113120 96616 113184
rect 96680 113120 96688 113184
rect 96368 113119 96688 113120
rect 127088 113184 127408 113185
rect 127088 113120 127096 113184
rect 127160 113120 127176 113184
rect 127240 113120 127256 113184
rect 127320 113120 127336 113184
rect 127400 113120 127408 113184
rect 127088 113119 127408 113120
rect 157808 113184 158128 113185
rect 157808 113120 157816 113184
rect 157880 113120 157896 113184
rect 157960 113120 157976 113184
rect 158040 113120 158056 113184
rect 158120 113120 158128 113184
rect 157808 113119 158128 113120
rect 19568 112640 19888 112641
rect 19568 112576 19576 112640
rect 19640 112576 19656 112640
rect 19720 112576 19736 112640
rect 19800 112576 19816 112640
rect 19880 112576 19888 112640
rect 19568 112575 19888 112576
rect 50288 112640 50608 112641
rect 50288 112576 50296 112640
rect 50360 112576 50376 112640
rect 50440 112576 50456 112640
rect 50520 112576 50536 112640
rect 50600 112576 50608 112640
rect 50288 112575 50608 112576
rect 81008 112640 81328 112641
rect 81008 112576 81016 112640
rect 81080 112576 81096 112640
rect 81160 112576 81176 112640
rect 81240 112576 81256 112640
rect 81320 112576 81328 112640
rect 81008 112575 81328 112576
rect 111728 112640 112048 112641
rect 111728 112576 111736 112640
rect 111800 112576 111816 112640
rect 111880 112576 111896 112640
rect 111960 112576 111976 112640
rect 112040 112576 112048 112640
rect 111728 112575 112048 112576
rect 142448 112640 142768 112641
rect 142448 112576 142456 112640
rect 142520 112576 142536 112640
rect 142600 112576 142616 112640
rect 142680 112576 142696 112640
rect 142760 112576 142768 112640
rect 142448 112575 142768 112576
rect 173168 112640 173488 112641
rect 173168 112576 173176 112640
rect 173240 112576 173256 112640
rect 173320 112576 173336 112640
rect 173400 112576 173416 112640
rect 173480 112576 173488 112640
rect 173168 112575 173488 112576
rect 4208 112096 4528 112097
rect 4208 112032 4216 112096
rect 4280 112032 4296 112096
rect 4360 112032 4376 112096
rect 4440 112032 4456 112096
rect 4520 112032 4528 112096
rect 4208 112031 4528 112032
rect 34928 112096 35248 112097
rect 34928 112032 34936 112096
rect 35000 112032 35016 112096
rect 35080 112032 35096 112096
rect 35160 112032 35176 112096
rect 35240 112032 35248 112096
rect 34928 112031 35248 112032
rect 65648 112096 65968 112097
rect 65648 112032 65656 112096
rect 65720 112032 65736 112096
rect 65800 112032 65816 112096
rect 65880 112032 65896 112096
rect 65960 112032 65968 112096
rect 65648 112031 65968 112032
rect 96368 112096 96688 112097
rect 96368 112032 96376 112096
rect 96440 112032 96456 112096
rect 96520 112032 96536 112096
rect 96600 112032 96616 112096
rect 96680 112032 96688 112096
rect 96368 112031 96688 112032
rect 127088 112096 127408 112097
rect 127088 112032 127096 112096
rect 127160 112032 127176 112096
rect 127240 112032 127256 112096
rect 127320 112032 127336 112096
rect 127400 112032 127408 112096
rect 127088 112031 127408 112032
rect 157808 112096 158128 112097
rect 157808 112032 157816 112096
rect 157880 112032 157896 112096
rect 157960 112032 157976 112096
rect 158040 112032 158056 112096
rect 158120 112032 158128 112096
rect 157808 112031 158128 112032
rect 19568 111552 19888 111553
rect 19568 111488 19576 111552
rect 19640 111488 19656 111552
rect 19720 111488 19736 111552
rect 19800 111488 19816 111552
rect 19880 111488 19888 111552
rect 19568 111487 19888 111488
rect 50288 111552 50608 111553
rect 50288 111488 50296 111552
rect 50360 111488 50376 111552
rect 50440 111488 50456 111552
rect 50520 111488 50536 111552
rect 50600 111488 50608 111552
rect 50288 111487 50608 111488
rect 81008 111552 81328 111553
rect 81008 111488 81016 111552
rect 81080 111488 81096 111552
rect 81160 111488 81176 111552
rect 81240 111488 81256 111552
rect 81320 111488 81328 111552
rect 81008 111487 81328 111488
rect 111728 111552 112048 111553
rect 111728 111488 111736 111552
rect 111800 111488 111816 111552
rect 111880 111488 111896 111552
rect 111960 111488 111976 111552
rect 112040 111488 112048 111552
rect 111728 111487 112048 111488
rect 142448 111552 142768 111553
rect 142448 111488 142456 111552
rect 142520 111488 142536 111552
rect 142600 111488 142616 111552
rect 142680 111488 142696 111552
rect 142760 111488 142768 111552
rect 142448 111487 142768 111488
rect 173168 111552 173488 111553
rect 173168 111488 173176 111552
rect 173240 111488 173256 111552
rect 173320 111488 173336 111552
rect 173400 111488 173416 111552
rect 173480 111488 173488 111552
rect 173168 111487 173488 111488
rect 4208 111008 4528 111009
rect 4208 110944 4216 111008
rect 4280 110944 4296 111008
rect 4360 110944 4376 111008
rect 4440 110944 4456 111008
rect 4520 110944 4528 111008
rect 4208 110943 4528 110944
rect 34928 111008 35248 111009
rect 34928 110944 34936 111008
rect 35000 110944 35016 111008
rect 35080 110944 35096 111008
rect 35160 110944 35176 111008
rect 35240 110944 35248 111008
rect 34928 110943 35248 110944
rect 65648 111008 65968 111009
rect 65648 110944 65656 111008
rect 65720 110944 65736 111008
rect 65800 110944 65816 111008
rect 65880 110944 65896 111008
rect 65960 110944 65968 111008
rect 65648 110943 65968 110944
rect 96368 111008 96688 111009
rect 96368 110944 96376 111008
rect 96440 110944 96456 111008
rect 96520 110944 96536 111008
rect 96600 110944 96616 111008
rect 96680 110944 96688 111008
rect 96368 110943 96688 110944
rect 127088 111008 127408 111009
rect 127088 110944 127096 111008
rect 127160 110944 127176 111008
rect 127240 110944 127256 111008
rect 127320 110944 127336 111008
rect 127400 110944 127408 111008
rect 127088 110943 127408 110944
rect 157808 111008 158128 111009
rect 157808 110944 157816 111008
rect 157880 110944 157896 111008
rect 157960 110944 157976 111008
rect 158040 110944 158056 111008
rect 158120 110944 158128 111008
rect 157808 110943 158128 110944
rect 19568 110464 19888 110465
rect 19568 110400 19576 110464
rect 19640 110400 19656 110464
rect 19720 110400 19736 110464
rect 19800 110400 19816 110464
rect 19880 110400 19888 110464
rect 19568 110399 19888 110400
rect 50288 110464 50608 110465
rect 50288 110400 50296 110464
rect 50360 110400 50376 110464
rect 50440 110400 50456 110464
rect 50520 110400 50536 110464
rect 50600 110400 50608 110464
rect 50288 110399 50608 110400
rect 81008 110464 81328 110465
rect 81008 110400 81016 110464
rect 81080 110400 81096 110464
rect 81160 110400 81176 110464
rect 81240 110400 81256 110464
rect 81320 110400 81328 110464
rect 81008 110399 81328 110400
rect 111728 110464 112048 110465
rect 111728 110400 111736 110464
rect 111800 110400 111816 110464
rect 111880 110400 111896 110464
rect 111960 110400 111976 110464
rect 112040 110400 112048 110464
rect 111728 110399 112048 110400
rect 142448 110464 142768 110465
rect 142448 110400 142456 110464
rect 142520 110400 142536 110464
rect 142600 110400 142616 110464
rect 142680 110400 142696 110464
rect 142760 110400 142768 110464
rect 142448 110399 142768 110400
rect 173168 110464 173488 110465
rect 173168 110400 173176 110464
rect 173240 110400 173256 110464
rect 173320 110400 173336 110464
rect 173400 110400 173416 110464
rect 173480 110400 173488 110464
rect 173168 110399 173488 110400
rect 4208 109920 4528 109921
rect 4208 109856 4216 109920
rect 4280 109856 4296 109920
rect 4360 109856 4376 109920
rect 4440 109856 4456 109920
rect 4520 109856 4528 109920
rect 4208 109855 4528 109856
rect 34928 109920 35248 109921
rect 34928 109856 34936 109920
rect 35000 109856 35016 109920
rect 35080 109856 35096 109920
rect 35160 109856 35176 109920
rect 35240 109856 35248 109920
rect 34928 109855 35248 109856
rect 65648 109920 65968 109921
rect 65648 109856 65656 109920
rect 65720 109856 65736 109920
rect 65800 109856 65816 109920
rect 65880 109856 65896 109920
rect 65960 109856 65968 109920
rect 65648 109855 65968 109856
rect 96368 109920 96688 109921
rect 96368 109856 96376 109920
rect 96440 109856 96456 109920
rect 96520 109856 96536 109920
rect 96600 109856 96616 109920
rect 96680 109856 96688 109920
rect 96368 109855 96688 109856
rect 127088 109920 127408 109921
rect 127088 109856 127096 109920
rect 127160 109856 127176 109920
rect 127240 109856 127256 109920
rect 127320 109856 127336 109920
rect 127400 109856 127408 109920
rect 127088 109855 127408 109856
rect 157808 109920 158128 109921
rect 157808 109856 157816 109920
rect 157880 109856 157896 109920
rect 157960 109856 157976 109920
rect 158040 109856 158056 109920
rect 158120 109856 158128 109920
rect 157808 109855 158128 109856
rect 19568 109376 19888 109377
rect 19568 109312 19576 109376
rect 19640 109312 19656 109376
rect 19720 109312 19736 109376
rect 19800 109312 19816 109376
rect 19880 109312 19888 109376
rect 19568 109311 19888 109312
rect 50288 109376 50608 109377
rect 50288 109312 50296 109376
rect 50360 109312 50376 109376
rect 50440 109312 50456 109376
rect 50520 109312 50536 109376
rect 50600 109312 50608 109376
rect 50288 109311 50608 109312
rect 81008 109376 81328 109377
rect 81008 109312 81016 109376
rect 81080 109312 81096 109376
rect 81160 109312 81176 109376
rect 81240 109312 81256 109376
rect 81320 109312 81328 109376
rect 81008 109311 81328 109312
rect 111728 109376 112048 109377
rect 111728 109312 111736 109376
rect 111800 109312 111816 109376
rect 111880 109312 111896 109376
rect 111960 109312 111976 109376
rect 112040 109312 112048 109376
rect 111728 109311 112048 109312
rect 142448 109376 142768 109377
rect 142448 109312 142456 109376
rect 142520 109312 142536 109376
rect 142600 109312 142616 109376
rect 142680 109312 142696 109376
rect 142760 109312 142768 109376
rect 142448 109311 142768 109312
rect 173168 109376 173488 109377
rect 173168 109312 173176 109376
rect 173240 109312 173256 109376
rect 173320 109312 173336 109376
rect 173400 109312 173416 109376
rect 173480 109312 173488 109376
rect 173168 109311 173488 109312
rect 4208 108832 4528 108833
rect 4208 108768 4216 108832
rect 4280 108768 4296 108832
rect 4360 108768 4376 108832
rect 4440 108768 4456 108832
rect 4520 108768 4528 108832
rect 4208 108767 4528 108768
rect 34928 108832 35248 108833
rect 34928 108768 34936 108832
rect 35000 108768 35016 108832
rect 35080 108768 35096 108832
rect 35160 108768 35176 108832
rect 35240 108768 35248 108832
rect 34928 108767 35248 108768
rect 65648 108832 65968 108833
rect 65648 108768 65656 108832
rect 65720 108768 65736 108832
rect 65800 108768 65816 108832
rect 65880 108768 65896 108832
rect 65960 108768 65968 108832
rect 65648 108767 65968 108768
rect 96368 108832 96688 108833
rect 96368 108768 96376 108832
rect 96440 108768 96456 108832
rect 96520 108768 96536 108832
rect 96600 108768 96616 108832
rect 96680 108768 96688 108832
rect 96368 108767 96688 108768
rect 127088 108832 127408 108833
rect 127088 108768 127096 108832
rect 127160 108768 127176 108832
rect 127240 108768 127256 108832
rect 127320 108768 127336 108832
rect 127400 108768 127408 108832
rect 127088 108767 127408 108768
rect 157808 108832 158128 108833
rect 157808 108768 157816 108832
rect 157880 108768 157896 108832
rect 157960 108768 157976 108832
rect 158040 108768 158056 108832
rect 158120 108768 158128 108832
rect 157808 108767 158128 108768
rect 19568 108288 19888 108289
rect 19568 108224 19576 108288
rect 19640 108224 19656 108288
rect 19720 108224 19736 108288
rect 19800 108224 19816 108288
rect 19880 108224 19888 108288
rect 19568 108223 19888 108224
rect 50288 108288 50608 108289
rect 50288 108224 50296 108288
rect 50360 108224 50376 108288
rect 50440 108224 50456 108288
rect 50520 108224 50536 108288
rect 50600 108224 50608 108288
rect 50288 108223 50608 108224
rect 81008 108288 81328 108289
rect 81008 108224 81016 108288
rect 81080 108224 81096 108288
rect 81160 108224 81176 108288
rect 81240 108224 81256 108288
rect 81320 108224 81328 108288
rect 81008 108223 81328 108224
rect 111728 108288 112048 108289
rect 111728 108224 111736 108288
rect 111800 108224 111816 108288
rect 111880 108224 111896 108288
rect 111960 108224 111976 108288
rect 112040 108224 112048 108288
rect 111728 108223 112048 108224
rect 142448 108288 142768 108289
rect 142448 108224 142456 108288
rect 142520 108224 142536 108288
rect 142600 108224 142616 108288
rect 142680 108224 142696 108288
rect 142760 108224 142768 108288
rect 142448 108223 142768 108224
rect 173168 108288 173488 108289
rect 173168 108224 173176 108288
rect 173240 108224 173256 108288
rect 173320 108224 173336 108288
rect 173400 108224 173416 108288
rect 173480 108224 173488 108288
rect 173168 108223 173488 108224
rect 4208 107744 4528 107745
rect 4208 107680 4216 107744
rect 4280 107680 4296 107744
rect 4360 107680 4376 107744
rect 4440 107680 4456 107744
rect 4520 107680 4528 107744
rect 4208 107679 4528 107680
rect 34928 107744 35248 107745
rect 34928 107680 34936 107744
rect 35000 107680 35016 107744
rect 35080 107680 35096 107744
rect 35160 107680 35176 107744
rect 35240 107680 35248 107744
rect 34928 107679 35248 107680
rect 65648 107744 65968 107745
rect 65648 107680 65656 107744
rect 65720 107680 65736 107744
rect 65800 107680 65816 107744
rect 65880 107680 65896 107744
rect 65960 107680 65968 107744
rect 65648 107679 65968 107680
rect 96368 107744 96688 107745
rect 96368 107680 96376 107744
rect 96440 107680 96456 107744
rect 96520 107680 96536 107744
rect 96600 107680 96616 107744
rect 96680 107680 96688 107744
rect 96368 107679 96688 107680
rect 127088 107744 127408 107745
rect 127088 107680 127096 107744
rect 127160 107680 127176 107744
rect 127240 107680 127256 107744
rect 127320 107680 127336 107744
rect 127400 107680 127408 107744
rect 127088 107679 127408 107680
rect 157808 107744 158128 107745
rect 157808 107680 157816 107744
rect 157880 107680 157896 107744
rect 157960 107680 157976 107744
rect 158040 107680 158056 107744
rect 158120 107680 158128 107744
rect 157808 107679 158128 107680
rect 19568 107200 19888 107201
rect 19568 107136 19576 107200
rect 19640 107136 19656 107200
rect 19720 107136 19736 107200
rect 19800 107136 19816 107200
rect 19880 107136 19888 107200
rect 19568 107135 19888 107136
rect 50288 107200 50608 107201
rect 50288 107136 50296 107200
rect 50360 107136 50376 107200
rect 50440 107136 50456 107200
rect 50520 107136 50536 107200
rect 50600 107136 50608 107200
rect 50288 107135 50608 107136
rect 81008 107200 81328 107201
rect 81008 107136 81016 107200
rect 81080 107136 81096 107200
rect 81160 107136 81176 107200
rect 81240 107136 81256 107200
rect 81320 107136 81328 107200
rect 81008 107135 81328 107136
rect 111728 107200 112048 107201
rect 111728 107136 111736 107200
rect 111800 107136 111816 107200
rect 111880 107136 111896 107200
rect 111960 107136 111976 107200
rect 112040 107136 112048 107200
rect 111728 107135 112048 107136
rect 142448 107200 142768 107201
rect 142448 107136 142456 107200
rect 142520 107136 142536 107200
rect 142600 107136 142616 107200
rect 142680 107136 142696 107200
rect 142760 107136 142768 107200
rect 142448 107135 142768 107136
rect 173168 107200 173488 107201
rect 173168 107136 173176 107200
rect 173240 107136 173256 107200
rect 173320 107136 173336 107200
rect 173400 107136 173416 107200
rect 173480 107136 173488 107200
rect 173168 107135 173488 107136
rect 4208 106656 4528 106657
rect 4208 106592 4216 106656
rect 4280 106592 4296 106656
rect 4360 106592 4376 106656
rect 4440 106592 4456 106656
rect 4520 106592 4528 106656
rect 4208 106591 4528 106592
rect 34928 106656 35248 106657
rect 34928 106592 34936 106656
rect 35000 106592 35016 106656
rect 35080 106592 35096 106656
rect 35160 106592 35176 106656
rect 35240 106592 35248 106656
rect 34928 106591 35248 106592
rect 65648 106656 65968 106657
rect 65648 106592 65656 106656
rect 65720 106592 65736 106656
rect 65800 106592 65816 106656
rect 65880 106592 65896 106656
rect 65960 106592 65968 106656
rect 65648 106591 65968 106592
rect 96368 106656 96688 106657
rect 96368 106592 96376 106656
rect 96440 106592 96456 106656
rect 96520 106592 96536 106656
rect 96600 106592 96616 106656
rect 96680 106592 96688 106656
rect 96368 106591 96688 106592
rect 127088 106656 127408 106657
rect 127088 106592 127096 106656
rect 127160 106592 127176 106656
rect 127240 106592 127256 106656
rect 127320 106592 127336 106656
rect 127400 106592 127408 106656
rect 127088 106591 127408 106592
rect 157808 106656 158128 106657
rect 157808 106592 157816 106656
rect 157880 106592 157896 106656
rect 157960 106592 157976 106656
rect 158040 106592 158056 106656
rect 158120 106592 158128 106656
rect 157808 106591 158128 106592
rect 19568 106112 19888 106113
rect 19568 106048 19576 106112
rect 19640 106048 19656 106112
rect 19720 106048 19736 106112
rect 19800 106048 19816 106112
rect 19880 106048 19888 106112
rect 19568 106047 19888 106048
rect 50288 106112 50608 106113
rect 50288 106048 50296 106112
rect 50360 106048 50376 106112
rect 50440 106048 50456 106112
rect 50520 106048 50536 106112
rect 50600 106048 50608 106112
rect 50288 106047 50608 106048
rect 81008 106112 81328 106113
rect 81008 106048 81016 106112
rect 81080 106048 81096 106112
rect 81160 106048 81176 106112
rect 81240 106048 81256 106112
rect 81320 106048 81328 106112
rect 81008 106047 81328 106048
rect 111728 106112 112048 106113
rect 111728 106048 111736 106112
rect 111800 106048 111816 106112
rect 111880 106048 111896 106112
rect 111960 106048 111976 106112
rect 112040 106048 112048 106112
rect 111728 106047 112048 106048
rect 142448 106112 142768 106113
rect 142448 106048 142456 106112
rect 142520 106048 142536 106112
rect 142600 106048 142616 106112
rect 142680 106048 142696 106112
rect 142760 106048 142768 106112
rect 142448 106047 142768 106048
rect 173168 106112 173488 106113
rect 173168 106048 173176 106112
rect 173240 106048 173256 106112
rect 173320 106048 173336 106112
rect 173400 106048 173416 106112
rect 173480 106048 173488 106112
rect 173168 106047 173488 106048
rect 4208 105568 4528 105569
rect 4208 105504 4216 105568
rect 4280 105504 4296 105568
rect 4360 105504 4376 105568
rect 4440 105504 4456 105568
rect 4520 105504 4528 105568
rect 4208 105503 4528 105504
rect 34928 105568 35248 105569
rect 34928 105504 34936 105568
rect 35000 105504 35016 105568
rect 35080 105504 35096 105568
rect 35160 105504 35176 105568
rect 35240 105504 35248 105568
rect 34928 105503 35248 105504
rect 65648 105568 65968 105569
rect 65648 105504 65656 105568
rect 65720 105504 65736 105568
rect 65800 105504 65816 105568
rect 65880 105504 65896 105568
rect 65960 105504 65968 105568
rect 65648 105503 65968 105504
rect 96368 105568 96688 105569
rect 96368 105504 96376 105568
rect 96440 105504 96456 105568
rect 96520 105504 96536 105568
rect 96600 105504 96616 105568
rect 96680 105504 96688 105568
rect 96368 105503 96688 105504
rect 127088 105568 127408 105569
rect 127088 105504 127096 105568
rect 127160 105504 127176 105568
rect 127240 105504 127256 105568
rect 127320 105504 127336 105568
rect 127400 105504 127408 105568
rect 127088 105503 127408 105504
rect 157808 105568 158128 105569
rect 157808 105504 157816 105568
rect 157880 105504 157896 105568
rect 157960 105504 157976 105568
rect 158040 105504 158056 105568
rect 158120 105504 158128 105568
rect 157808 105503 158128 105504
rect 19568 105024 19888 105025
rect 19568 104960 19576 105024
rect 19640 104960 19656 105024
rect 19720 104960 19736 105024
rect 19800 104960 19816 105024
rect 19880 104960 19888 105024
rect 19568 104959 19888 104960
rect 50288 105024 50608 105025
rect 50288 104960 50296 105024
rect 50360 104960 50376 105024
rect 50440 104960 50456 105024
rect 50520 104960 50536 105024
rect 50600 104960 50608 105024
rect 50288 104959 50608 104960
rect 81008 105024 81328 105025
rect 81008 104960 81016 105024
rect 81080 104960 81096 105024
rect 81160 104960 81176 105024
rect 81240 104960 81256 105024
rect 81320 104960 81328 105024
rect 81008 104959 81328 104960
rect 111728 105024 112048 105025
rect 111728 104960 111736 105024
rect 111800 104960 111816 105024
rect 111880 104960 111896 105024
rect 111960 104960 111976 105024
rect 112040 104960 112048 105024
rect 111728 104959 112048 104960
rect 142448 105024 142768 105025
rect 142448 104960 142456 105024
rect 142520 104960 142536 105024
rect 142600 104960 142616 105024
rect 142680 104960 142696 105024
rect 142760 104960 142768 105024
rect 142448 104959 142768 104960
rect 173168 105024 173488 105025
rect 173168 104960 173176 105024
rect 173240 104960 173256 105024
rect 173320 104960 173336 105024
rect 173400 104960 173416 105024
rect 173480 104960 173488 105024
rect 173168 104959 173488 104960
rect 4208 104480 4528 104481
rect 4208 104416 4216 104480
rect 4280 104416 4296 104480
rect 4360 104416 4376 104480
rect 4440 104416 4456 104480
rect 4520 104416 4528 104480
rect 4208 104415 4528 104416
rect 34928 104480 35248 104481
rect 34928 104416 34936 104480
rect 35000 104416 35016 104480
rect 35080 104416 35096 104480
rect 35160 104416 35176 104480
rect 35240 104416 35248 104480
rect 34928 104415 35248 104416
rect 65648 104480 65968 104481
rect 65648 104416 65656 104480
rect 65720 104416 65736 104480
rect 65800 104416 65816 104480
rect 65880 104416 65896 104480
rect 65960 104416 65968 104480
rect 65648 104415 65968 104416
rect 96368 104480 96688 104481
rect 96368 104416 96376 104480
rect 96440 104416 96456 104480
rect 96520 104416 96536 104480
rect 96600 104416 96616 104480
rect 96680 104416 96688 104480
rect 96368 104415 96688 104416
rect 127088 104480 127408 104481
rect 127088 104416 127096 104480
rect 127160 104416 127176 104480
rect 127240 104416 127256 104480
rect 127320 104416 127336 104480
rect 127400 104416 127408 104480
rect 127088 104415 127408 104416
rect 157808 104480 158128 104481
rect 157808 104416 157816 104480
rect 157880 104416 157896 104480
rect 157960 104416 157976 104480
rect 158040 104416 158056 104480
rect 158120 104416 158128 104480
rect 157808 104415 158128 104416
rect 19568 103936 19888 103937
rect 19568 103872 19576 103936
rect 19640 103872 19656 103936
rect 19720 103872 19736 103936
rect 19800 103872 19816 103936
rect 19880 103872 19888 103936
rect 19568 103871 19888 103872
rect 50288 103936 50608 103937
rect 50288 103872 50296 103936
rect 50360 103872 50376 103936
rect 50440 103872 50456 103936
rect 50520 103872 50536 103936
rect 50600 103872 50608 103936
rect 50288 103871 50608 103872
rect 81008 103936 81328 103937
rect 81008 103872 81016 103936
rect 81080 103872 81096 103936
rect 81160 103872 81176 103936
rect 81240 103872 81256 103936
rect 81320 103872 81328 103936
rect 81008 103871 81328 103872
rect 111728 103936 112048 103937
rect 111728 103872 111736 103936
rect 111800 103872 111816 103936
rect 111880 103872 111896 103936
rect 111960 103872 111976 103936
rect 112040 103872 112048 103936
rect 111728 103871 112048 103872
rect 142448 103936 142768 103937
rect 142448 103872 142456 103936
rect 142520 103872 142536 103936
rect 142600 103872 142616 103936
rect 142680 103872 142696 103936
rect 142760 103872 142768 103936
rect 142448 103871 142768 103872
rect 173168 103936 173488 103937
rect 173168 103872 173176 103936
rect 173240 103872 173256 103936
rect 173320 103872 173336 103936
rect 173400 103872 173416 103936
rect 173480 103872 173488 103936
rect 173168 103871 173488 103872
rect 4208 103392 4528 103393
rect 4208 103328 4216 103392
rect 4280 103328 4296 103392
rect 4360 103328 4376 103392
rect 4440 103328 4456 103392
rect 4520 103328 4528 103392
rect 4208 103327 4528 103328
rect 34928 103392 35248 103393
rect 34928 103328 34936 103392
rect 35000 103328 35016 103392
rect 35080 103328 35096 103392
rect 35160 103328 35176 103392
rect 35240 103328 35248 103392
rect 34928 103327 35248 103328
rect 65648 103392 65968 103393
rect 65648 103328 65656 103392
rect 65720 103328 65736 103392
rect 65800 103328 65816 103392
rect 65880 103328 65896 103392
rect 65960 103328 65968 103392
rect 65648 103327 65968 103328
rect 96368 103392 96688 103393
rect 96368 103328 96376 103392
rect 96440 103328 96456 103392
rect 96520 103328 96536 103392
rect 96600 103328 96616 103392
rect 96680 103328 96688 103392
rect 96368 103327 96688 103328
rect 127088 103392 127408 103393
rect 127088 103328 127096 103392
rect 127160 103328 127176 103392
rect 127240 103328 127256 103392
rect 127320 103328 127336 103392
rect 127400 103328 127408 103392
rect 127088 103327 127408 103328
rect 157808 103392 158128 103393
rect 157808 103328 157816 103392
rect 157880 103328 157896 103392
rect 157960 103328 157976 103392
rect 158040 103328 158056 103392
rect 158120 103328 158128 103392
rect 157808 103327 158128 103328
rect 19568 102848 19888 102849
rect 19568 102784 19576 102848
rect 19640 102784 19656 102848
rect 19720 102784 19736 102848
rect 19800 102784 19816 102848
rect 19880 102784 19888 102848
rect 19568 102783 19888 102784
rect 50288 102848 50608 102849
rect 50288 102784 50296 102848
rect 50360 102784 50376 102848
rect 50440 102784 50456 102848
rect 50520 102784 50536 102848
rect 50600 102784 50608 102848
rect 50288 102783 50608 102784
rect 81008 102848 81328 102849
rect 81008 102784 81016 102848
rect 81080 102784 81096 102848
rect 81160 102784 81176 102848
rect 81240 102784 81256 102848
rect 81320 102784 81328 102848
rect 81008 102783 81328 102784
rect 111728 102848 112048 102849
rect 111728 102784 111736 102848
rect 111800 102784 111816 102848
rect 111880 102784 111896 102848
rect 111960 102784 111976 102848
rect 112040 102784 112048 102848
rect 111728 102783 112048 102784
rect 142448 102848 142768 102849
rect 142448 102784 142456 102848
rect 142520 102784 142536 102848
rect 142600 102784 142616 102848
rect 142680 102784 142696 102848
rect 142760 102784 142768 102848
rect 142448 102783 142768 102784
rect 173168 102848 173488 102849
rect 173168 102784 173176 102848
rect 173240 102784 173256 102848
rect 173320 102784 173336 102848
rect 173400 102784 173416 102848
rect 173480 102784 173488 102848
rect 173168 102783 173488 102784
rect 4208 102304 4528 102305
rect 4208 102240 4216 102304
rect 4280 102240 4296 102304
rect 4360 102240 4376 102304
rect 4440 102240 4456 102304
rect 4520 102240 4528 102304
rect 4208 102239 4528 102240
rect 34928 102304 35248 102305
rect 34928 102240 34936 102304
rect 35000 102240 35016 102304
rect 35080 102240 35096 102304
rect 35160 102240 35176 102304
rect 35240 102240 35248 102304
rect 34928 102239 35248 102240
rect 65648 102304 65968 102305
rect 65648 102240 65656 102304
rect 65720 102240 65736 102304
rect 65800 102240 65816 102304
rect 65880 102240 65896 102304
rect 65960 102240 65968 102304
rect 65648 102239 65968 102240
rect 96368 102304 96688 102305
rect 96368 102240 96376 102304
rect 96440 102240 96456 102304
rect 96520 102240 96536 102304
rect 96600 102240 96616 102304
rect 96680 102240 96688 102304
rect 96368 102239 96688 102240
rect 127088 102304 127408 102305
rect 127088 102240 127096 102304
rect 127160 102240 127176 102304
rect 127240 102240 127256 102304
rect 127320 102240 127336 102304
rect 127400 102240 127408 102304
rect 127088 102239 127408 102240
rect 157808 102304 158128 102305
rect 157808 102240 157816 102304
rect 157880 102240 157896 102304
rect 157960 102240 157976 102304
rect 158040 102240 158056 102304
rect 158120 102240 158128 102304
rect 157808 102239 158128 102240
rect 19568 101760 19888 101761
rect 19568 101696 19576 101760
rect 19640 101696 19656 101760
rect 19720 101696 19736 101760
rect 19800 101696 19816 101760
rect 19880 101696 19888 101760
rect 19568 101695 19888 101696
rect 50288 101760 50608 101761
rect 50288 101696 50296 101760
rect 50360 101696 50376 101760
rect 50440 101696 50456 101760
rect 50520 101696 50536 101760
rect 50600 101696 50608 101760
rect 50288 101695 50608 101696
rect 81008 101760 81328 101761
rect 81008 101696 81016 101760
rect 81080 101696 81096 101760
rect 81160 101696 81176 101760
rect 81240 101696 81256 101760
rect 81320 101696 81328 101760
rect 81008 101695 81328 101696
rect 111728 101760 112048 101761
rect 111728 101696 111736 101760
rect 111800 101696 111816 101760
rect 111880 101696 111896 101760
rect 111960 101696 111976 101760
rect 112040 101696 112048 101760
rect 111728 101695 112048 101696
rect 142448 101760 142768 101761
rect 142448 101696 142456 101760
rect 142520 101696 142536 101760
rect 142600 101696 142616 101760
rect 142680 101696 142696 101760
rect 142760 101696 142768 101760
rect 142448 101695 142768 101696
rect 173168 101760 173488 101761
rect 173168 101696 173176 101760
rect 173240 101696 173256 101760
rect 173320 101696 173336 101760
rect 173400 101696 173416 101760
rect 173480 101696 173488 101760
rect 173168 101695 173488 101696
rect 4208 101216 4528 101217
rect 4208 101152 4216 101216
rect 4280 101152 4296 101216
rect 4360 101152 4376 101216
rect 4440 101152 4456 101216
rect 4520 101152 4528 101216
rect 4208 101151 4528 101152
rect 34928 101216 35248 101217
rect 34928 101152 34936 101216
rect 35000 101152 35016 101216
rect 35080 101152 35096 101216
rect 35160 101152 35176 101216
rect 35240 101152 35248 101216
rect 34928 101151 35248 101152
rect 65648 101216 65968 101217
rect 65648 101152 65656 101216
rect 65720 101152 65736 101216
rect 65800 101152 65816 101216
rect 65880 101152 65896 101216
rect 65960 101152 65968 101216
rect 65648 101151 65968 101152
rect 96368 101216 96688 101217
rect 96368 101152 96376 101216
rect 96440 101152 96456 101216
rect 96520 101152 96536 101216
rect 96600 101152 96616 101216
rect 96680 101152 96688 101216
rect 96368 101151 96688 101152
rect 127088 101216 127408 101217
rect 127088 101152 127096 101216
rect 127160 101152 127176 101216
rect 127240 101152 127256 101216
rect 127320 101152 127336 101216
rect 127400 101152 127408 101216
rect 127088 101151 127408 101152
rect 157808 101216 158128 101217
rect 157808 101152 157816 101216
rect 157880 101152 157896 101216
rect 157960 101152 157976 101216
rect 158040 101152 158056 101216
rect 158120 101152 158128 101216
rect 157808 101151 158128 101152
rect 19568 100672 19888 100673
rect 19568 100608 19576 100672
rect 19640 100608 19656 100672
rect 19720 100608 19736 100672
rect 19800 100608 19816 100672
rect 19880 100608 19888 100672
rect 19568 100607 19888 100608
rect 50288 100672 50608 100673
rect 50288 100608 50296 100672
rect 50360 100608 50376 100672
rect 50440 100608 50456 100672
rect 50520 100608 50536 100672
rect 50600 100608 50608 100672
rect 50288 100607 50608 100608
rect 81008 100672 81328 100673
rect 81008 100608 81016 100672
rect 81080 100608 81096 100672
rect 81160 100608 81176 100672
rect 81240 100608 81256 100672
rect 81320 100608 81328 100672
rect 81008 100607 81328 100608
rect 111728 100672 112048 100673
rect 111728 100608 111736 100672
rect 111800 100608 111816 100672
rect 111880 100608 111896 100672
rect 111960 100608 111976 100672
rect 112040 100608 112048 100672
rect 111728 100607 112048 100608
rect 142448 100672 142768 100673
rect 142448 100608 142456 100672
rect 142520 100608 142536 100672
rect 142600 100608 142616 100672
rect 142680 100608 142696 100672
rect 142760 100608 142768 100672
rect 142448 100607 142768 100608
rect 173168 100672 173488 100673
rect 173168 100608 173176 100672
rect 173240 100608 173256 100672
rect 173320 100608 173336 100672
rect 173400 100608 173416 100672
rect 173480 100608 173488 100672
rect 173168 100607 173488 100608
rect 4208 100128 4528 100129
rect 4208 100064 4216 100128
rect 4280 100064 4296 100128
rect 4360 100064 4376 100128
rect 4440 100064 4456 100128
rect 4520 100064 4528 100128
rect 4208 100063 4528 100064
rect 34928 100128 35248 100129
rect 34928 100064 34936 100128
rect 35000 100064 35016 100128
rect 35080 100064 35096 100128
rect 35160 100064 35176 100128
rect 35240 100064 35248 100128
rect 34928 100063 35248 100064
rect 65648 100128 65968 100129
rect 65648 100064 65656 100128
rect 65720 100064 65736 100128
rect 65800 100064 65816 100128
rect 65880 100064 65896 100128
rect 65960 100064 65968 100128
rect 65648 100063 65968 100064
rect 96368 100128 96688 100129
rect 96368 100064 96376 100128
rect 96440 100064 96456 100128
rect 96520 100064 96536 100128
rect 96600 100064 96616 100128
rect 96680 100064 96688 100128
rect 96368 100063 96688 100064
rect 127088 100128 127408 100129
rect 127088 100064 127096 100128
rect 127160 100064 127176 100128
rect 127240 100064 127256 100128
rect 127320 100064 127336 100128
rect 127400 100064 127408 100128
rect 127088 100063 127408 100064
rect 157808 100128 158128 100129
rect 157808 100064 157816 100128
rect 157880 100064 157896 100128
rect 157960 100064 157976 100128
rect 158040 100064 158056 100128
rect 158120 100064 158128 100128
rect 157808 100063 158128 100064
rect 19568 99584 19888 99585
rect 19568 99520 19576 99584
rect 19640 99520 19656 99584
rect 19720 99520 19736 99584
rect 19800 99520 19816 99584
rect 19880 99520 19888 99584
rect 19568 99519 19888 99520
rect 50288 99584 50608 99585
rect 50288 99520 50296 99584
rect 50360 99520 50376 99584
rect 50440 99520 50456 99584
rect 50520 99520 50536 99584
rect 50600 99520 50608 99584
rect 50288 99519 50608 99520
rect 81008 99584 81328 99585
rect 81008 99520 81016 99584
rect 81080 99520 81096 99584
rect 81160 99520 81176 99584
rect 81240 99520 81256 99584
rect 81320 99520 81328 99584
rect 81008 99519 81328 99520
rect 111728 99584 112048 99585
rect 111728 99520 111736 99584
rect 111800 99520 111816 99584
rect 111880 99520 111896 99584
rect 111960 99520 111976 99584
rect 112040 99520 112048 99584
rect 111728 99519 112048 99520
rect 142448 99584 142768 99585
rect 142448 99520 142456 99584
rect 142520 99520 142536 99584
rect 142600 99520 142616 99584
rect 142680 99520 142696 99584
rect 142760 99520 142768 99584
rect 142448 99519 142768 99520
rect 173168 99584 173488 99585
rect 173168 99520 173176 99584
rect 173240 99520 173256 99584
rect 173320 99520 173336 99584
rect 173400 99520 173416 99584
rect 173480 99520 173488 99584
rect 173168 99519 173488 99520
rect 4208 99040 4528 99041
rect 4208 98976 4216 99040
rect 4280 98976 4296 99040
rect 4360 98976 4376 99040
rect 4440 98976 4456 99040
rect 4520 98976 4528 99040
rect 4208 98975 4528 98976
rect 34928 99040 35248 99041
rect 34928 98976 34936 99040
rect 35000 98976 35016 99040
rect 35080 98976 35096 99040
rect 35160 98976 35176 99040
rect 35240 98976 35248 99040
rect 34928 98975 35248 98976
rect 65648 99040 65968 99041
rect 65648 98976 65656 99040
rect 65720 98976 65736 99040
rect 65800 98976 65816 99040
rect 65880 98976 65896 99040
rect 65960 98976 65968 99040
rect 65648 98975 65968 98976
rect 96368 99040 96688 99041
rect 96368 98976 96376 99040
rect 96440 98976 96456 99040
rect 96520 98976 96536 99040
rect 96600 98976 96616 99040
rect 96680 98976 96688 99040
rect 96368 98975 96688 98976
rect 127088 99040 127408 99041
rect 127088 98976 127096 99040
rect 127160 98976 127176 99040
rect 127240 98976 127256 99040
rect 127320 98976 127336 99040
rect 127400 98976 127408 99040
rect 127088 98975 127408 98976
rect 157808 99040 158128 99041
rect 157808 98976 157816 99040
rect 157880 98976 157896 99040
rect 157960 98976 157976 99040
rect 158040 98976 158056 99040
rect 158120 98976 158128 99040
rect 157808 98975 158128 98976
rect 19568 98496 19888 98497
rect 19568 98432 19576 98496
rect 19640 98432 19656 98496
rect 19720 98432 19736 98496
rect 19800 98432 19816 98496
rect 19880 98432 19888 98496
rect 19568 98431 19888 98432
rect 50288 98496 50608 98497
rect 50288 98432 50296 98496
rect 50360 98432 50376 98496
rect 50440 98432 50456 98496
rect 50520 98432 50536 98496
rect 50600 98432 50608 98496
rect 50288 98431 50608 98432
rect 81008 98496 81328 98497
rect 81008 98432 81016 98496
rect 81080 98432 81096 98496
rect 81160 98432 81176 98496
rect 81240 98432 81256 98496
rect 81320 98432 81328 98496
rect 81008 98431 81328 98432
rect 111728 98496 112048 98497
rect 111728 98432 111736 98496
rect 111800 98432 111816 98496
rect 111880 98432 111896 98496
rect 111960 98432 111976 98496
rect 112040 98432 112048 98496
rect 111728 98431 112048 98432
rect 142448 98496 142768 98497
rect 142448 98432 142456 98496
rect 142520 98432 142536 98496
rect 142600 98432 142616 98496
rect 142680 98432 142696 98496
rect 142760 98432 142768 98496
rect 142448 98431 142768 98432
rect 173168 98496 173488 98497
rect 173168 98432 173176 98496
rect 173240 98432 173256 98496
rect 173320 98432 173336 98496
rect 173400 98432 173416 98496
rect 173480 98432 173488 98496
rect 173168 98431 173488 98432
rect 4208 97952 4528 97953
rect 4208 97888 4216 97952
rect 4280 97888 4296 97952
rect 4360 97888 4376 97952
rect 4440 97888 4456 97952
rect 4520 97888 4528 97952
rect 4208 97887 4528 97888
rect 34928 97952 35248 97953
rect 34928 97888 34936 97952
rect 35000 97888 35016 97952
rect 35080 97888 35096 97952
rect 35160 97888 35176 97952
rect 35240 97888 35248 97952
rect 34928 97887 35248 97888
rect 65648 97952 65968 97953
rect 65648 97888 65656 97952
rect 65720 97888 65736 97952
rect 65800 97888 65816 97952
rect 65880 97888 65896 97952
rect 65960 97888 65968 97952
rect 65648 97887 65968 97888
rect 96368 97952 96688 97953
rect 96368 97888 96376 97952
rect 96440 97888 96456 97952
rect 96520 97888 96536 97952
rect 96600 97888 96616 97952
rect 96680 97888 96688 97952
rect 96368 97887 96688 97888
rect 127088 97952 127408 97953
rect 127088 97888 127096 97952
rect 127160 97888 127176 97952
rect 127240 97888 127256 97952
rect 127320 97888 127336 97952
rect 127400 97888 127408 97952
rect 127088 97887 127408 97888
rect 157808 97952 158128 97953
rect 157808 97888 157816 97952
rect 157880 97888 157896 97952
rect 157960 97888 157976 97952
rect 158040 97888 158056 97952
rect 158120 97888 158128 97952
rect 157808 97887 158128 97888
rect 19568 97408 19888 97409
rect 19568 97344 19576 97408
rect 19640 97344 19656 97408
rect 19720 97344 19736 97408
rect 19800 97344 19816 97408
rect 19880 97344 19888 97408
rect 19568 97343 19888 97344
rect 50288 97408 50608 97409
rect 50288 97344 50296 97408
rect 50360 97344 50376 97408
rect 50440 97344 50456 97408
rect 50520 97344 50536 97408
rect 50600 97344 50608 97408
rect 50288 97343 50608 97344
rect 81008 97408 81328 97409
rect 81008 97344 81016 97408
rect 81080 97344 81096 97408
rect 81160 97344 81176 97408
rect 81240 97344 81256 97408
rect 81320 97344 81328 97408
rect 81008 97343 81328 97344
rect 111728 97408 112048 97409
rect 111728 97344 111736 97408
rect 111800 97344 111816 97408
rect 111880 97344 111896 97408
rect 111960 97344 111976 97408
rect 112040 97344 112048 97408
rect 111728 97343 112048 97344
rect 142448 97408 142768 97409
rect 142448 97344 142456 97408
rect 142520 97344 142536 97408
rect 142600 97344 142616 97408
rect 142680 97344 142696 97408
rect 142760 97344 142768 97408
rect 142448 97343 142768 97344
rect 173168 97408 173488 97409
rect 173168 97344 173176 97408
rect 173240 97344 173256 97408
rect 173320 97344 173336 97408
rect 173400 97344 173416 97408
rect 173480 97344 173488 97408
rect 173168 97343 173488 97344
rect 4208 96864 4528 96865
rect 4208 96800 4216 96864
rect 4280 96800 4296 96864
rect 4360 96800 4376 96864
rect 4440 96800 4456 96864
rect 4520 96800 4528 96864
rect 4208 96799 4528 96800
rect 34928 96864 35248 96865
rect 34928 96800 34936 96864
rect 35000 96800 35016 96864
rect 35080 96800 35096 96864
rect 35160 96800 35176 96864
rect 35240 96800 35248 96864
rect 34928 96799 35248 96800
rect 65648 96864 65968 96865
rect 65648 96800 65656 96864
rect 65720 96800 65736 96864
rect 65800 96800 65816 96864
rect 65880 96800 65896 96864
rect 65960 96800 65968 96864
rect 65648 96799 65968 96800
rect 96368 96864 96688 96865
rect 96368 96800 96376 96864
rect 96440 96800 96456 96864
rect 96520 96800 96536 96864
rect 96600 96800 96616 96864
rect 96680 96800 96688 96864
rect 96368 96799 96688 96800
rect 127088 96864 127408 96865
rect 127088 96800 127096 96864
rect 127160 96800 127176 96864
rect 127240 96800 127256 96864
rect 127320 96800 127336 96864
rect 127400 96800 127408 96864
rect 127088 96799 127408 96800
rect 157808 96864 158128 96865
rect 157808 96800 157816 96864
rect 157880 96800 157896 96864
rect 157960 96800 157976 96864
rect 158040 96800 158056 96864
rect 158120 96800 158128 96864
rect 157808 96799 158128 96800
rect 19568 96320 19888 96321
rect 19568 96256 19576 96320
rect 19640 96256 19656 96320
rect 19720 96256 19736 96320
rect 19800 96256 19816 96320
rect 19880 96256 19888 96320
rect 19568 96255 19888 96256
rect 50288 96320 50608 96321
rect 50288 96256 50296 96320
rect 50360 96256 50376 96320
rect 50440 96256 50456 96320
rect 50520 96256 50536 96320
rect 50600 96256 50608 96320
rect 50288 96255 50608 96256
rect 81008 96320 81328 96321
rect 81008 96256 81016 96320
rect 81080 96256 81096 96320
rect 81160 96256 81176 96320
rect 81240 96256 81256 96320
rect 81320 96256 81328 96320
rect 81008 96255 81328 96256
rect 111728 96320 112048 96321
rect 111728 96256 111736 96320
rect 111800 96256 111816 96320
rect 111880 96256 111896 96320
rect 111960 96256 111976 96320
rect 112040 96256 112048 96320
rect 111728 96255 112048 96256
rect 142448 96320 142768 96321
rect 142448 96256 142456 96320
rect 142520 96256 142536 96320
rect 142600 96256 142616 96320
rect 142680 96256 142696 96320
rect 142760 96256 142768 96320
rect 142448 96255 142768 96256
rect 173168 96320 173488 96321
rect 173168 96256 173176 96320
rect 173240 96256 173256 96320
rect 173320 96256 173336 96320
rect 173400 96256 173416 96320
rect 173480 96256 173488 96320
rect 173168 96255 173488 96256
rect 4208 95776 4528 95777
rect 4208 95712 4216 95776
rect 4280 95712 4296 95776
rect 4360 95712 4376 95776
rect 4440 95712 4456 95776
rect 4520 95712 4528 95776
rect 4208 95711 4528 95712
rect 34928 95776 35248 95777
rect 34928 95712 34936 95776
rect 35000 95712 35016 95776
rect 35080 95712 35096 95776
rect 35160 95712 35176 95776
rect 35240 95712 35248 95776
rect 34928 95711 35248 95712
rect 65648 95776 65968 95777
rect 65648 95712 65656 95776
rect 65720 95712 65736 95776
rect 65800 95712 65816 95776
rect 65880 95712 65896 95776
rect 65960 95712 65968 95776
rect 65648 95711 65968 95712
rect 96368 95776 96688 95777
rect 96368 95712 96376 95776
rect 96440 95712 96456 95776
rect 96520 95712 96536 95776
rect 96600 95712 96616 95776
rect 96680 95712 96688 95776
rect 96368 95711 96688 95712
rect 127088 95776 127408 95777
rect 127088 95712 127096 95776
rect 127160 95712 127176 95776
rect 127240 95712 127256 95776
rect 127320 95712 127336 95776
rect 127400 95712 127408 95776
rect 127088 95711 127408 95712
rect 157808 95776 158128 95777
rect 157808 95712 157816 95776
rect 157880 95712 157896 95776
rect 157960 95712 157976 95776
rect 158040 95712 158056 95776
rect 158120 95712 158128 95776
rect 157808 95711 158128 95712
rect 19568 95232 19888 95233
rect 19568 95168 19576 95232
rect 19640 95168 19656 95232
rect 19720 95168 19736 95232
rect 19800 95168 19816 95232
rect 19880 95168 19888 95232
rect 19568 95167 19888 95168
rect 50288 95232 50608 95233
rect 50288 95168 50296 95232
rect 50360 95168 50376 95232
rect 50440 95168 50456 95232
rect 50520 95168 50536 95232
rect 50600 95168 50608 95232
rect 50288 95167 50608 95168
rect 81008 95232 81328 95233
rect 81008 95168 81016 95232
rect 81080 95168 81096 95232
rect 81160 95168 81176 95232
rect 81240 95168 81256 95232
rect 81320 95168 81328 95232
rect 81008 95167 81328 95168
rect 111728 95232 112048 95233
rect 111728 95168 111736 95232
rect 111800 95168 111816 95232
rect 111880 95168 111896 95232
rect 111960 95168 111976 95232
rect 112040 95168 112048 95232
rect 111728 95167 112048 95168
rect 142448 95232 142768 95233
rect 142448 95168 142456 95232
rect 142520 95168 142536 95232
rect 142600 95168 142616 95232
rect 142680 95168 142696 95232
rect 142760 95168 142768 95232
rect 142448 95167 142768 95168
rect 173168 95232 173488 95233
rect 173168 95168 173176 95232
rect 173240 95168 173256 95232
rect 173320 95168 173336 95232
rect 173400 95168 173416 95232
rect 173480 95168 173488 95232
rect 173168 95167 173488 95168
rect 4208 94688 4528 94689
rect 4208 94624 4216 94688
rect 4280 94624 4296 94688
rect 4360 94624 4376 94688
rect 4440 94624 4456 94688
rect 4520 94624 4528 94688
rect 4208 94623 4528 94624
rect 34928 94688 35248 94689
rect 34928 94624 34936 94688
rect 35000 94624 35016 94688
rect 35080 94624 35096 94688
rect 35160 94624 35176 94688
rect 35240 94624 35248 94688
rect 34928 94623 35248 94624
rect 65648 94688 65968 94689
rect 65648 94624 65656 94688
rect 65720 94624 65736 94688
rect 65800 94624 65816 94688
rect 65880 94624 65896 94688
rect 65960 94624 65968 94688
rect 65648 94623 65968 94624
rect 96368 94688 96688 94689
rect 96368 94624 96376 94688
rect 96440 94624 96456 94688
rect 96520 94624 96536 94688
rect 96600 94624 96616 94688
rect 96680 94624 96688 94688
rect 96368 94623 96688 94624
rect 127088 94688 127408 94689
rect 127088 94624 127096 94688
rect 127160 94624 127176 94688
rect 127240 94624 127256 94688
rect 127320 94624 127336 94688
rect 127400 94624 127408 94688
rect 127088 94623 127408 94624
rect 157808 94688 158128 94689
rect 157808 94624 157816 94688
rect 157880 94624 157896 94688
rect 157960 94624 157976 94688
rect 158040 94624 158056 94688
rect 158120 94624 158128 94688
rect 157808 94623 158128 94624
rect 19568 94144 19888 94145
rect 19568 94080 19576 94144
rect 19640 94080 19656 94144
rect 19720 94080 19736 94144
rect 19800 94080 19816 94144
rect 19880 94080 19888 94144
rect 19568 94079 19888 94080
rect 50288 94144 50608 94145
rect 50288 94080 50296 94144
rect 50360 94080 50376 94144
rect 50440 94080 50456 94144
rect 50520 94080 50536 94144
rect 50600 94080 50608 94144
rect 50288 94079 50608 94080
rect 81008 94144 81328 94145
rect 81008 94080 81016 94144
rect 81080 94080 81096 94144
rect 81160 94080 81176 94144
rect 81240 94080 81256 94144
rect 81320 94080 81328 94144
rect 81008 94079 81328 94080
rect 111728 94144 112048 94145
rect 111728 94080 111736 94144
rect 111800 94080 111816 94144
rect 111880 94080 111896 94144
rect 111960 94080 111976 94144
rect 112040 94080 112048 94144
rect 111728 94079 112048 94080
rect 142448 94144 142768 94145
rect 142448 94080 142456 94144
rect 142520 94080 142536 94144
rect 142600 94080 142616 94144
rect 142680 94080 142696 94144
rect 142760 94080 142768 94144
rect 142448 94079 142768 94080
rect 173168 94144 173488 94145
rect 173168 94080 173176 94144
rect 173240 94080 173256 94144
rect 173320 94080 173336 94144
rect 173400 94080 173416 94144
rect 173480 94080 173488 94144
rect 173168 94079 173488 94080
rect 4208 93600 4528 93601
rect 4208 93536 4216 93600
rect 4280 93536 4296 93600
rect 4360 93536 4376 93600
rect 4440 93536 4456 93600
rect 4520 93536 4528 93600
rect 4208 93535 4528 93536
rect 34928 93600 35248 93601
rect 34928 93536 34936 93600
rect 35000 93536 35016 93600
rect 35080 93536 35096 93600
rect 35160 93536 35176 93600
rect 35240 93536 35248 93600
rect 34928 93535 35248 93536
rect 65648 93600 65968 93601
rect 65648 93536 65656 93600
rect 65720 93536 65736 93600
rect 65800 93536 65816 93600
rect 65880 93536 65896 93600
rect 65960 93536 65968 93600
rect 65648 93535 65968 93536
rect 96368 93600 96688 93601
rect 96368 93536 96376 93600
rect 96440 93536 96456 93600
rect 96520 93536 96536 93600
rect 96600 93536 96616 93600
rect 96680 93536 96688 93600
rect 96368 93535 96688 93536
rect 127088 93600 127408 93601
rect 127088 93536 127096 93600
rect 127160 93536 127176 93600
rect 127240 93536 127256 93600
rect 127320 93536 127336 93600
rect 127400 93536 127408 93600
rect 127088 93535 127408 93536
rect 157808 93600 158128 93601
rect 157808 93536 157816 93600
rect 157880 93536 157896 93600
rect 157960 93536 157976 93600
rect 158040 93536 158056 93600
rect 158120 93536 158128 93600
rect 157808 93535 158128 93536
rect 19568 93056 19888 93057
rect 19568 92992 19576 93056
rect 19640 92992 19656 93056
rect 19720 92992 19736 93056
rect 19800 92992 19816 93056
rect 19880 92992 19888 93056
rect 19568 92991 19888 92992
rect 50288 93056 50608 93057
rect 50288 92992 50296 93056
rect 50360 92992 50376 93056
rect 50440 92992 50456 93056
rect 50520 92992 50536 93056
rect 50600 92992 50608 93056
rect 50288 92991 50608 92992
rect 81008 93056 81328 93057
rect 81008 92992 81016 93056
rect 81080 92992 81096 93056
rect 81160 92992 81176 93056
rect 81240 92992 81256 93056
rect 81320 92992 81328 93056
rect 81008 92991 81328 92992
rect 111728 93056 112048 93057
rect 111728 92992 111736 93056
rect 111800 92992 111816 93056
rect 111880 92992 111896 93056
rect 111960 92992 111976 93056
rect 112040 92992 112048 93056
rect 111728 92991 112048 92992
rect 142448 93056 142768 93057
rect 142448 92992 142456 93056
rect 142520 92992 142536 93056
rect 142600 92992 142616 93056
rect 142680 92992 142696 93056
rect 142760 92992 142768 93056
rect 142448 92991 142768 92992
rect 173168 93056 173488 93057
rect 173168 92992 173176 93056
rect 173240 92992 173256 93056
rect 173320 92992 173336 93056
rect 173400 92992 173416 93056
rect 173480 92992 173488 93056
rect 173168 92991 173488 92992
rect 4208 92512 4528 92513
rect 4208 92448 4216 92512
rect 4280 92448 4296 92512
rect 4360 92448 4376 92512
rect 4440 92448 4456 92512
rect 4520 92448 4528 92512
rect 4208 92447 4528 92448
rect 34928 92512 35248 92513
rect 34928 92448 34936 92512
rect 35000 92448 35016 92512
rect 35080 92448 35096 92512
rect 35160 92448 35176 92512
rect 35240 92448 35248 92512
rect 34928 92447 35248 92448
rect 65648 92512 65968 92513
rect 65648 92448 65656 92512
rect 65720 92448 65736 92512
rect 65800 92448 65816 92512
rect 65880 92448 65896 92512
rect 65960 92448 65968 92512
rect 65648 92447 65968 92448
rect 96368 92512 96688 92513
rect 96368 92448 96376 92512
rect 96440 92448 96456 92512
rect 96520 92448 96536 92512
rect 96600 92448 96616 92512
rect 96680 92448 96688 92512
rect 96368 92447 96688 92448
rect 127088 92512 127408 92513
rect 127088 92448 127096 92512
rect 127160 92448 127176 92512
rect 127240 92448 127256 92512
rect 127320 92448 127336 92512
rect 127400 92448 127408 92512
rect 127088 92447 127408 92448
rect 157808 92512 158128 92513
rect 157808 92448 157816 92512
rect 157880 92448 157896 92512
rect 157960 92448 157976 92512
rect 158040 92448 158056 92512
rect 158120 92448 158128 92512
rect 157808 92447 158128 92448
rect 19568 91968 19888 91969
rect 19568 91904 19576 91968
rect 19640 91904 19656 91968
rect 19720 91904 19736 91968
rect 19800 91904 19816 91968
rect 19880 91904 19888 91968
rect 19568 91903 19888 91904
rect 50288 91968 50608 91969
rect 50288 91904 50296 91968
rect 50360 91904 50376 91968
rect 50440 91904 50456 91968
rect 50520 91904 50536 91968
rect 50600 91904 50608 91968
rect 50288 91903 50608 91904
rect 81008 91968 81328 91969
rect 81008 91904 81016 91968
rect 81080 91904 81096 91968
rect 81160 91904 81176 91968
rect 81240 91904 81256 91968
rect 81320 91904 81328 91968
rect 81008 91903 81328 91904
rect 111728 91968 112048 91969
rect 111728 91904 111736 91968
rect 111800 91904 111816 91968
rect 111880 91904 111896 91968
rect 111960 91904 111976 91968
rect 112040 91904 112048 91968
rect 111728 91903 112048 91904
rect 142448 91968 142768 91969
rect 142448 91904 142456 91968
rect 142520 91904 142536 91968
rect 142600 91904 142616 91968
rect 142680 91904 142696 91968
rect 142760 91904 142768 91968
rect 142448 91903 142768 91904
rect 173168 91968 173488 91969
rect 173168 91904 173176 91968
rect 173240 91904 173256 91968
rect 173320 91904 173336 91968
rect 173400 91904 173416 91968
rect 173480 91904 173488 91968
rect 173168 91903 173488 91904
rect 4208 91424 4528 91425
rect 4208 91360 4216 91424
rect 4280 91360 4296 91424
rect 4360 91360 4376 91424
rect 4440 91360 4456 91424
rect 4520 91360 4528 91424
rect 4208 91359 4528 91360
rect 34928 91424 35248 91425
rect 34928 91360 34936 91424
rect 35000 91360 35016 91424
rect 35080 91360 35096 91424
rect 35160 91360 35176 91424
rect 35240 91360 35248 91424
rect 34928 91359 35248 91360
rect 65648 91424 65968 91425
rect 65648 91360 65656 91424
rect 65720 91360 65736 91424
rect 65800 91360 65816 91424
rect 65880 91360 65896 91424
rect 65960 91360 65968 91424
rect 65648 91359 65968 91360
rect 96368 91424 96688 91425
rect 96368 91360 96376 91424
rect 96440 91360 96456 91424
rect 96520 91360 96536 91424
rect 96600 91360 96616 91424
rect 96680 91360 96688 91424
rect 96368 91359 96688 91360
rect 127088 91424 127408 91425
rect 127088 91360 127096 91424
rect 127160 91360 127176 91424
rect 127240 91360 127256 91424
rect 127320 91360 127336 91424
rect 127400 91360 127408 91424
rect 127088 91359 127408 91360
rect 157808 91424 158128 91425
rect 157808 91360 157816 91424
rect 157880 91360 157896 91424
rect 157960 91360 157976 91424
rect 158040 91360 158056 91424
rect 158120 91360 158128 91424
rect 157808 91359 158128 91360
rect 19568 90880 19888 90881
rect 19568 90816 19576 90880
rect 19640 90816 19656 90880
rect 19720 90816 19736 90880
rect 19800 90816 19816 90880
rect 19880 90816 19888 90880
rect 19568 90815 19888 90816
rect 50288 90880 50608 90881
rect 50288 90816 50296 90880
rect 50360 90816 50376 90880
rect 50440 90816 50456 90880
rect 50520 90816 50536 90880
rect 50600 90816 50608 90880
rect 50288 90815 50608 90816
rect 81008 90880 81328 90881
rect 81008 90816 81016 90880
rect 81080 90816 81096 90880
rect 81160 90816 81176 90880
rect 81240 90816 81256 90880
rect 81320 90816 81328 90880
rect 81008 90815 81328 90816
rect 111728 90880 112048 90881
rect 111728 90816 111736 90880
rect 111800 90816 111816 90880
rect 111880 90816 111896 90880
rect 111960 90816 111976 90880
rect 112040 90816 112048 90880
rect 111728 90815 112048 90816
rect 142448 90880 142768 90881
rect 142448 90816 142456 90880
rect 142520 90816 142536 90880
rect 142600 90816 142616 90880
rect 142680 90816 142696 90880
rect 142760 90816 142768 90880
rect 142448 90815 142768 90816
rect 173168 90880 173488 90881
rect 173168 90816 173176 90880
rect 173240 90816 173256 90880
rect 173320 90816 173336 90880
rect 173400 90816 173416 90880
rect 173480 90816 173488 90880
rect 173168 90815 173488 90816
rect 4208 90336 4528 90337
rect 4208 90272 4216 90336
rect 4280 90272 4296 90336
rect 4360 90272 4376 90336
rect 4440 90272 4456 90336
rect 4520 90272 4528 90336
rect 4208 90271 4528 90272
rect 34928 90336 35248 90337
rect 34928 90272 34936 90336
rect 35000 90272 35016 90336
rect 35080 90272 35096 90336
rect 35160 90272 35176 90336
rect 35240 90272 35248 90336
rect 34928 90271 35248 90272
rect 65648 90336 65968 90337
rect 65648 90272 65656 90336
rect 65720 90272 65736 90336
rect 65800 90272 65816 90336
rect 65880 90272 65896 90336
rect 65960 90272 65968 90336
rect 65648 90271 65968 90272
rect 96368 90336 96688 90337
rect 96368 90272 96376 90336
rect 96440 90272 96456 90336
rect 96520 90272 96536 90336
rect 96600 90272 96616 90336
rect 96680 90272 96688 90336
rect 96368 90271 96688 90272
rect 127088 90336 127408 90337
rect 127088 90272 127096 90336
rect 127160 90272 127176 90336
rect 127240 90272 127256 90336
rect 127320 90272 127336 90336
rect 127400 90272 127408 90336
rect 127088 90271 127408 90272
rect 157808 90336 158128 90337
rect 157808 90272 157816 90336
rect 157880 90272 157896 90336
rect 157960 90272 157976 90336
rect 158040 90272 158056 90336
rect 158120 90272 158128 90336
rect 157808 90271 158128 90272
rect 19568 89792 19888 89793
rect 19568 89728 19576 89792
rect 19640 89728 19656 89792
rect 19720 89728 19736 89792
rect 19800 89728 19816 89792
rect 19880 89728 19888 89792
rect 19568 89727 19888 89728
rect 50288 89792 50608 89793
rect 50288 89728 50296 89792
rect 50360 89728 50376 89792
rect 50440 89728 50456 89792
rect 50520 89728 50536 89792
rect 50600 89728 50608 89792
rect 50288 89727 50608 89728
rect 81008 89792 81328 89793
rect 81008 89728 81016 89792
rect 81080 89728 81096 89792
rect 81160 89728 81176 89792
rect 81240 89728 81256 89792
rect 81320 89728 81328 89792
rect 81008 89727 81328 89728
rect 111728 89792 112048 89793
rect 111728 89728 111736 89792
rect 111800 89728 111816 89792
rect 111880 89728 111896 89792
rect 111960 89728 111976 89792
rect 112040 89728 112048 89792
rect 111728 89727 112048 89728
rect 142448 89792 142768 89793
rect 142448 89728 142456 89792
rect 142520 89728 142536 89792
rect 142600 89728 142616 89792
rect 142680 89728 142696 89792
rect 142760 89728 142768 89792
rect 142448 89727 142768 89728
rect 173168 89792 173488 89793
rect 173168 89728 173176 89792
rect 173240 89728 173256 89792
rect 173320 89728 173336 89792
rect 173400 89728 173416 89792
rect 173480 89728 173488 89792
rect 173168 89727 173488 89728
rect 4208 89248 4528 89249
rect 4208 89184 4216 89248
rect 4280 89184 4296 89248
rect 4360 89184 4376 89248
rect 4440 89184 4456 89248
rect 4520 89184 4528 89248
rect 4208 89183 4528 89184
rect 34928 89248 35248 89249
rect 34928 89184 34936 89248
rect 35000 89184 35016 89248
rect 35080 89184 35096 89248
rect 35160 89184 35176 89248
rect 35240 89184 35248 89248
rect 34928 89183 35248 89184
rect 65648 89248 65968 89249
rect 65648 89184 65656 89248
rect 65720 89184 65736 89248
rect 65800 89184 65816 89248
rect 65880 89184 65896 89248
rect 65960 89184 65968 89248
rect 65648 89183 65968 89184
rect 96368 89248 96688 89249
rect 96368 89184 96376 89248
rect 96440 89184 96456 89248
rect 96520 89184 96536 89248
rect 96600 89184 96616 89248
rect 96680 89184 96688 89248
rect 96368 89183 96688 89184
rect 127088 89248 127408 89249
rect 127088 89184 127096 89248
rect 127160 89184 127176 89248
rect 127240 89184 127256 89248
rect 127320 89184 127336 89248
rect 127400 89184 127408 89248
rect 127088 89183 127408 89184
rect 157808 89248 158128 89249
rect 157808 89184 157816 89248
rect 157880 89184 157896 89248
rect 157960 89184 157976 89248
rect 158040 89184 158056 89248
rect 158120 89184 158128 89248
rect 157808 89183 158128 89184
rect 19568 88704 19888 88705
rect 19568 88640 19576 88704
rect 19640 88640 19656 88704
rect 19720 88640 19736 88704
rect 19800 88640 19816 88704
rect 19880 88640 19888 88704
rect 19568 88639 19888 88640
rect 50288 88704 50608 88705
rect 50288 88640 50296 88704
rect 50360 88640 50376 88704
rect 50440 88640 50456 88704
rect 50520 88640 50536 88704
rect 50600 88640 50608 88704
rect 50288 88639 50608 88640
rect 81008 88704 81328 88705
rect 81008 88640 81016 88704
rect 81080 88640 81096 88704
rect 81160 88640 81176 88704
rect 81240 88640 81256 88704
rect 81320 88640 81328 88704
rect 81008 88639 81328 88640
rect 111728 88704 112048 88705
rect 111728 88640 111736 88704
rect 111800 88640 111816 88704
rect 111880 88640 111896 88704
rect 111960 88640 111976 88704
rect 112040 88640 112048 88704
rect 111728 88639 112048 88640
rect 142448 88704 142768 88705
rect 142448 88640 142456 88704
rect 142520 88640 142536 88704
rect 142600 88640 142616 88704
rect 142680 88640 142696 88704
rect 142760 88640 142768 88704
rect 142448 88639 142768 88640
rect 173168 88704 173488 88705
rect 173168 88640 173176 88704
rect 173240 88640 173256 88704
rect 173320 88640 173336 88704
rect 173400 88640 173416 88704
rect 173480 88640 173488 88704
rect 173168 88639 173488 88640
rect 4208 88160 4528 88161
rect 4208 88096 4216 88160
rect 4280 88096 4296 88160
rect 4360 88096 4376 88160
rect 4440 88096 4456 88160
rect 4520 88096 4528 88160
rect 4208 88095 4528 88096
rect 34928 88160 35248 88161
rect 34928 88096 34936 88160
rect 35000 88096 35016 88160
rect 35080 88096 35096 88160
rect 35160 88096 35176 88160
rect 35240 88096 35248 88160
rect 34928 88095 35248 88096
rect 65648 88160 65968 88161
rect 65648 88096 65656 88160
rect 65720 88096 65736 88160
rect 65800 88096 65816 88160
rect 65880 88096 65896 88160
rect 65960 88096 65968 88160
rect 65648 88095 65968 88096
rect 96368 88160 96688 88161
rect 96368 88096 96376 88160
rect 96440 88096 96456 88160
rect 96520 88096 96536 88160
rect 96600 88096 96616 88160
rect 96680 88096 96688 88160
rect 96368 88095 96688 88096
rect 127088 88160 127408 88161
rect 127088 88096 127096 88160
rect 127160 88096 127176 88160
rect 127240 88096 127256 88160
rect 127320 88096 127336 88160
rect 127400 88096 127408 88160
rect 127088 88095 127408 88096
rect 157808 88160 158128 88161
rect 157808 88096 157816 88160
rect 157880 88096 157896 88160
rect 157960 88096 157976 88160
rect 158040 88096 158056 88160
rect 158120 88096 158128 88160
rect 157808 88095 158128 88096
rect 19568 87616 19888 87617
rect 19568 87552 19576 87616
rect 19640 87552 19656 87616
rect 19720 87552 19736 87616
rect 19800 87552 19816 87616
rect 19880 87552 19888 87616
rect 19568 87551 19888 87552
rect 50288 87616 50608 87617
rect 50288 87552 50296 87616
rect 50360 87552 50376 87616
rect 50440 87552 50456 87616
rect 50520 87552 50536 87616
rect 50600 87552 50608 87616
rect 50288 87551 50608 87552
rect 81008 87616 81328 87617
rect 81008 87552 81016 87616
rect 81080 87552 81096 87616
rect 81160 87552 81176 87616
rect 81240 87552 81256 87616
rect 81320 87552 81328 87616
rect 81008 87551 81328 87552
rect 111728 87616 112048 87617
rect 111728 87552 111736 87616
rect 111800 87552 111816 87616
rect 111880 87552 111896 87616
rect 111960 87552 111976 87616
rect 112040 87552 112048 87616
rect 111728 87551 112048 87552
rect 142448 87616 142768 87617
rect 142448 87552 142456 87616
rect 142520 87552 142536 87616
rect 142600 87552 142616 87616
rect 142680 87552 142696 87616
rect 142760 87552 142768 87616
rect 142448 87551 142768 87552
rect 173168 87616 173488 87617
rect 173168 87552 173176 87616
rect 173240 87552 173256 87616
rect 173320 87552 173336 87616
rect 173400 87552 173416 87616
rect 173480 87552 173488 87616
rect 173168 87551 173488 87552
rect 4208 87072 4528 87073
rect 4208 87008 4216 87072
rect 4280 87008 4296 87072
rect 4360 87008 4376 87072
rect 4440 87008 4456 87072
rect 4520 87008 4528 87072
rect 4208 87007 4528 87008
rect 34928 87072 35248 87073
rect 34928 87008 34936 87072
rect 35000 87008 35016 87072
rect 35080 87008 35096 87072
rect 35160 87008 35176 87072
rect 35240 87008 35248 87072
rect 34928 87007 35248 87008
rect 65648 87072 65968 87073
rect 65648 87008 65656 87072
rect 65720 87008 65736 87072
rect 65800 87008 65816 87072
rect 65880 87008 65896 87072
rect 65960 87008 65968 87072
rect 65648 87007 65968 87008
rect 96368 87072 96688 87073
rect 96368 87008 96376 87072
rect 96440 87008 96456 87072
rect 96520 87008 96536 87072
rect 96600 87008 96616 87072
rect 96680 87008 96688 87072
rect 96368 87007 96688 87008
rect 127088 87072 127408 87073
rect 127088 87008 127096 87072
rect 127160 87008 127176 87072
rect 127240 87008 127256 87072
rect 127320 87008 127336 87072
rect 127400 87008 127408 87072
rect 127088 87007 127408 87008
rect 157808 87072 158128 87073
rect 157808 87008 157816 87072
rect 157880 87008 157896 87072
rect 157960 87008 157976 87072
rect 158040 87008 158056 87072
rect 158120 87008 158128 87072
rect 157808 87007 158128 87008
rect 19568 86528 19888 86529
rect 19568 86464 19576 86528
rect 19640 86464 19656 86528
rect 19720 86464 19736 86528
rect 19800 86464 19816 86528
rect 19880 86464 19888 86528
rect 19568 86463 19888 86464
rect 50288 86528 50608 86529
rect 50288 86464 50296 86528
rect 50360 86464 50376 86528
rect 50440 86464 50456 86528
rect 50520 86464 50536 86528
rect 50600 86464 50608 86528
rect 50288 86463 50608 86464
rect 81008 86528 81328 86529
rect 81008 86464 81016 86528
rect 81080 86464 81096 86528
rect 81160 86464 81176 86528
rect 81240 86464 81256 86528
rect 81320 86464 81328 86528
rect 81008 86463 81328 86464
rect 111728 86528 112048 86529
rect 111728 86464 111736 86528
rect 111800 86464 111816 86528
rect 111880 86464 111896 86528
rect 111960 86464 111976 86528
rect 112040 86464 112048 86528
rect 111728 86463 112048 86464
rect 142448 86528 142768 86529
rect 142448 86464 142456 86528
rect 142520 86464 142536 86528
rect 142600 86464 142616 86528
rect 142680 86464 142696 86528
rect 142760 86464 142768 86528
rect 142448 86463 142768 86464
rect 173168 86528 173488 86529
rect 173168 86464 173176 86528
rect 173240 86464 173256 86528
rect 173320 86464 173336 86528
rect 173400 86464 173416 86528
rect 173480 86464 173488 86528
rect 173168 86463 173488 86464
rect 4208 85984 4528 85985
rect 4208 85920 4216 85984
rect 4280 85920 4296 85984
rect 4360 85920 4376 85984
rect 4440 85920 4456 85984
rect 4520 85920 4528 85984
rect 4208 85919 4528 85920
rect 34928 85984 35248 85985
rect 34928 85920 34936 85984
rect 35000 85920 35016 85984
rect 35080 85920 35096 85984
rect 35160 85920 35176 85984
rect 35240 85920 35248 85984
rect 34928 85919 35248 85920
rect 65648 85984 65968 85985
rect 65648 85920 65656 85984
rect 65720 85920 65736 85984
rect 65800 85920 65816 85984
rect 65880 85920 65896 85984
rect 65960 85920 65968 85984
rect 65648 85919 65968 85920
rect 96368 85984 96688 85985
rect 96368 85920 96376 85984
rect 96440 85920 96456 85984
rect 96520 85920 96536 85984
rect 96600 85920 96616 85984
rect 96680 85920 96688 85984
rect 96368 85919 96688 85920
rect 127088 85984 127408 85985
rect 127088 85920 127096 85984
rect 127160 85920 127176 85984
rect 127240 85920 127256 85984
rect 127320 85920 127336 85984
rect 127400 85920 127408 85984
rect 127088 85919 127408 85920
rect 157808 85984 158128 85985
rect 157808 85920 157816 85984
rect 157880 85920 157896 85984
rect 157960 85920 157976 85984
rect 158040 85920 158056 85984
rect 158120 85920 158128 85984
rect 157808 85919 158128 85920
rect 19568 85440 19888 85441
rect 19568 85376 19576 85440
rect 19640 85376 19656 85440
rect 19720 85376 19736 85440
rect 19800 85376 19816 85440
rect 19880 85376 19888 85440
rect 19568 85375 19888 85376
rect 50288 85440 50608 85441
rect 50288 85376 50296 85440
rect 50360 85376 50376 85440
rect 50440 85376 50456 85440
rect 50520 85376 50536 85440
rect 50600 85376 50608 85440
rect 50288 85375 50608 85376
rect 81008 85440 81328 85441
rect 81008 85376 81016 85440
rect 81080 85376 81096 85440
rect 81160 85376 81176 85440
rect 81240 85376 81256 85440
rect 81320 85376 81328 85440
rect 81008 85375 81328 85376
rect 111728 85440 112048 85441
rect 111728 85376 111736 85440
rect 111800 85376 111816 85440
rect 111880 85376 111896 85440
rect 111960 85376 111976 85440
rect 112040 85376 112048 85440
rect 111728 85375 112048 85376
rect 142448 85440 142768 85441
rect 142448 85376 142456 85440
rect 142520 85376 142536 85440
rect 142600 85376 142616 85440
rect 142680 85376 142696 85440
rect 142760 85376 142768 85440
rect 142448 85375 142768 85376
rect 173168 85440 173488 85441
rect 173168 85376 173176 85440
rect 173240 85376 173256 85440
rect 173320 85376 173336 85440
rect 173400 85376 173416 85440
rect 173480 85376 173488 85440
rect 173168 85375 173488 85376
rect 4208 84896 4528 84897
rect 4208 84832 4216 84896
rect 4280 84832 4296 84896
rect 4360 84832 4376 84896
rect 4440 84832 4456 84896
rect 4520 84832 4528 84896
rect 4208 84831 4528 84832
rect 34928 84896 35248 84897
rect 34928 84832 34936 84896
rect 35000 84832 35016 84896
rect 35080 84832 35096 84896
rect 35160 84832 35176 84896
rect 35240 84832 35248 84896
rect 34928 84831 35248 84832
rect 65648 84896 65968 84897
rect 65648 84832 65656 84896
rect 65720 84832 65736 84896
rect 65800 84832 65816 84896
rect 65880 84832 65896 84896
rect 65960 84832 65968 84896
rect 65648 84831 65968 84832
rect 96368 84896 96688 84897
rect 96368 84832 96376 84896
rect 96440 84832 96456 84896
rect 96520 84832 96536 84896
rect 96600 84832 96616 84896
rect 96680 84832 96688 84896
rect 96368 84831 96688 84832
rect 127088 84896 127408 84897
rect 127088 84832 127096 84896
rect 127160 84832 127176 84896
rect 127240 84832 127256 84896
rect 127320 84832 127336 84896
rect 127400 84832 127408 84896
rect 127088 84831 127408 84832
rect 157808 84896 158128 84897
rect 157808 84832 157816 84896
rect 157880 84832 157896 84896
rect 157960 84832 157976 84896
rect 158040 84832 158056 84896
rect 158120 84832 158128 84896
rect 157808 84831 158128 84832
rect 19568 84352 19888 84353
rect 19568 84288 19576 84352
rect 19640 84288 19656 84352
rect 19720 84288 19736 84352
rect 19800 84288 19816 84352
rect 19880 84288 19888 84352
rect 19568 84287 19888 84288
rect 50288 84352 50608 84353
rect 50288 84288 50296 84352
rect 50360 84288 50376 84352
rect 50440 84288 50456 84352
rect 50520 84288 50536 84352
rect 50600 84288 50608 84352
rect 50288 84287 50608 84288
rect 81008 84352 81328 84353
rect 81008 84288 81016 84352
rect 81080 84288 81096 84352
rect 81160 84288 81176 84352
rect 81240 84288 81256 84352
rect 81320 84288 81328 84352
rect 81008 84287 81328 84288
rect 111728 84352 112048 84353
rect 111728 84288 111736 84352
rect 111800 84288 111816 84352
rect 111880 84288 111896 84352
rect 111960 84288 111976 84352
rect 112040 84288 112048 84352
rect 111728 84287 112048 84288
rect 142448 84352 142768 84353
rect 142448 84288 142456 84352
rect 142520 84288 142536 84352
rect 142600 84288 142616 84352
rect 142680 84288 142696 84352
rect 142760 84288 142768 84352
rect 142448 84287 142768 84288
rect 173168 84352 173488 84353
rect 173168 84288 173176 84352
rect 173240 84288 173256 84352
rect 173320 84288 173336 84352
rect 173400 84288 173416 84352
rect 173480 84288 173488 84352
rect 173168 84287 173488 84288
rect 4208 83808 4528 83809
rect 4208 83744 4216 83808
rect 4280 83744 4296 83808
rect 4360 83744 4376 83808
rect 4440 83744 4456 83808
rect 4520 83744 4528 83808
rect 4208 83743 4528 83744
rect 34928 83808 35248 83809
rect 34928 83744 34936 83808
rect 35000 83744 35016 83808
rect 35080 83744 35096 83808
rect 35160 83744 35176 83808
rect 35240 83744 35248 83808
rect 34928 83743 35248 83744
rect 65648 83808 65968 83809
rect 65648 83744 65656 83808
rect 65720 83744 65736 83808
rect 65800 83744 65816 83808
rect 65880 83744 65896 83808
rect 65960 83744 65968 83808
rect 65648 83743 65968 83744
rect 96368 83808 96688 83809
rect 96368 83744 96376 83808
rect 96440 83744 96456 83808
rect 96520 83744 96536 83808
rect 96600 83744 96616 83808
rect 96680 83744 96688 83808
rect 96368 83743 96688 83744
rect 127088 83808 127408 83809
rect 127088 83744 127096 83808
rect 127160 83744 127176 83808
rect 127240 83744 127256 83808
rect 127320 83744 127336 83808
rect 127400 83744 127408 83808
rect 127088 83743 127408 83744
rect 157808 83808 158128 83809
rect 157808 83744 157816 83808
rect 157880 83744 157896 83808
rect 157960 83744 157976 83808
rect 158040 83744 158056 83808
rect 158120 83744 158128 83808
rect 157808 83743 158128 83744
rect 19568 83264 19888 83265
rect 19568 83200 19576 83264
rect 19640 83200 19656 83264
rect 19720 83200 19736 83264
rect 19800 83200 19816 83264
rect 19880 83200 19888 83264
rect 19568 83199 19888 83200
rect 50288 83264 50608 83265
rect 50288 83200 50296 83264
rect 50360 83200 50376 83264
rect 50440 83200 50456 83264
rect 50520 83200 50536 83264
rect 50600 83200 50608 83264
rect 50288 83199 50608 83200
rect 81008 83264 81328 83265
rect 81008 83200 81016 83264
rect 81080 83200 81096 83264
rect 81160 83200 81176 83264
rect 81240 83200 81256 83264
rect 81320 83200 81328 83264
rect 81008 83199 81328 83200
rect 111728 83264 112048 83265
rect 111728 83200 111736 83264
rect 111800 83200 111816 83264
rect 111880 83200 111896 83264
rect 111960 83200 111976 83264
rect 112040 83200 112048 83264
rect 111728 83199 112048 83200
rect 142448 83264 142768 83265
rect 142448 83200 142456 83264
rect 142520 83200 142536 83264
rect 142600 83200 142616 83264
rect 142680 83200 142696 83264
rect 142760 83200 142768 83264
rect 142448 83199 142768 83200
rect 173168 83264 173488 83265
rect 173168 83200 173176 83264
rect 173240 83200 173256 83264
rect 173320 83200 173336 83264
rect 173400 83200 173416 83264
rect 173480 83200 173488 83264
rect 173168 83199 173488 83200
rect 4208 82720 4528 82721
rect 4208 82656 4216 82720
rect 4280 82656 4296 82720
rect 4360 82656 4376 82720
rect 4440 82656 4456 82720
rect 4520 82656 4528 82720
rect 4208 82655 4528 82656
rect 34928 82720 35248 82721
rect 34928 82656 34936 82720
rect 35000 82656 35016 82720
rect 35080 82656 35096 82720
rect 35160 82656 35176 82720
rect 35240 82656 35248 82720
rect 34928 82655 35248 82656
rect 65648 82720 65968 82721
rect 65648 82656 65656 82720
rect 65720 82656 65736 82720
rect 65800 82656 65816 82720
rect 65880 82656 65896 82720
rect 65960 82656 65968 82720
rect 65648 82655 65968 82656
rect 96368 82720 96688 82721
rect 96368 82656 96376 82720
rect 96440 82656 96456 82720
rect 96520 82656 96536 82720
rect 96600 82656 96616 82720
rect 96680 82656 96688 82720
rect 96368 82655 96688 82656
rect 127088 82720 127408 82721
rect 127088 82656 127096 82720
rect 127160 82656 127176 82720
rect 127240 82656 127256 82720
rect 127320 82656 127336 82720
rect 127400 82656 127408 82720
rect 127088 82655 127408 82656
rect 157808 82720 158128 82721
rect 157808 82656 157816 82720
rect 157880 82656 157896 82720
rect 157960 82656 157976 82720
rect 158040 82656 158056 82720
rect 158120 82656 158128 82720
rect 157808 82655 158128 82656
rect 19568 82176 19888 82177
rect 19568 82112 19576 82176
rect 19640 82112 19656 82176
rect 19720 82112 19736 82176
rect 19800 82112 19816 82176
rect 19880 82112 19888 82176
rect 19568 82111 19888 82112
rect 50288 82176 50608 82177
rect 50288 82112 50296 82176
rect 50360 82112 50376 82176
rect 50440 82112 50456 82176
rect 50520 82112 50536 82176
rect 50600 82112 50608 82176
rect 50288 82111 50608 82112
rect 81008 82176 81328 82177
rect 81008 82112 81016 82176
rect 81080 82112 81096 82176
rect 81160 82112 81176 82176
rect 81240 82112 81256 82176
rect 81320 82112 81328 82176
rect 81008 82111 81328 82112
rect 111728 82176 112048 82177
rect 111728 82112 111736 82176
rect 111800 82112 111816 82176
rect 111880 82112 111896 82176
rect 111960 82112 111976 82176
rect 112040 82112 112048 82176
rect 111728 82111 112048 82112
rect 142448 82176 142768 82177
rect 142448 82112 142456 82176
rect 142520 82112 142536 82176
rect 142600 82112 142616 82176
rect 142680 82112 142696 82176
rect 142760 82112 142768 82176
rect 142448 82111 142768 82112
rect 173168 82176 173488 82177
rect 173168 82112 173176 82176
rect 173240 82112 173256 82176
rect 173320 82112 173336 82176
rect 173400 82112 173416 82176
rect 173480 82112 173488 82176
rect 173168 82111 173488 82112
rect 4208 81632 4528 81633
rect 4208 81568 4216 81632
rect 4280 81568 4296 81632
rect 4360 81568 4376 81632
rect 4440 81568 4456 81632
rect 4520 81568 4528 81632
rect 4208 81567 4528 81568
rect 34928 81632 35248 81633
rect 34928 81568 34936 81632
rect 35000 81568 35016 81632
rect 35080 81568 35096 81632
rect 35160 81568 35176 81632
rect 35240 81568 35248 81632
rect 34928 81567 35248 81568
rect 65648 81632 65968 81633
rect 65648 81568 65656 81632
rect 65720 81568 65736 81632
rect 65800 81568 65816 81632
rect 65880 81568 65896 81632
rect 65960 81568 65968 81632
rect 65648 81567 65968 81568
rect 96368 81632 96688 81633
rect 96368 81568 96376 81632
rect 96440 81568 96456 81632
rect 96520 81568 96536 81632
rect 96600 81568 96616 81632
rect 96680 81568 96688 81632
rect 96368 81567 96688 81568
rect 127088 81632 127408 81633
rect 127088 81568 127096 81632
rect 127160 81568 127176 81632
rect 127240 81568 127256 81632
rect 127320 81568 127336 81632
rect 127400 81568 127408 81632
rect 127088 81567 127408 81568
rect 157808 81632 158128 81633
rect 157808 81568 157816 81632
rect 157880 81568 157896 81632
rect 157960 81568 157976 81632
rect 158040 81568 158056 81632
rect 158120 81568 158128 81632
rect 157808 81567 158128 81568
rect 19568 81088 19888 81089
rect 19568 81024 19576 81088
rect 19640 81024 19656 81088
rect 19720 81024 19736 81088
rect 19800 81024 19816 81088
rect 19880 81024 19888 81088
rect 19568 81023 19888 81024
rect 50288 81088 50608 81089
rect 50288 81024 50296 81088
rect 50360 81024 50376 81088
rect 50440 81024 50456 81088
rect 50520 81024 50536 81088
rect 50600 81024 50608 81088
rect 50288 81023 50608 81024
rect 81008 81088 81328 81089
rect 81008 81024 81016 81088
rect 81080 81024 81096 81088
rect 81160 81024 81176 81088
rect 81240 81024 81256 81088
rect 81320 81024 81328 81088
rect 81008 81023 81328 81024
rect 111728 81088 112048 81089
rect 111728 81024 111736 81088
rect 111800 81024 111816 81088
rect 111880 81024 111896 81088
rect 111960 81024 111976 81088
rect 112040 81024 112048 81088
rect 111728 81023 112048 81024
rect 142448 81088 142768 81089
rect 142448 81024 142456 81088
rect 142520 81024 142536 81088
rect 142600 81024 142616 81088
rect 142680 81024 142696 81088
rect 142760 81024 142768 81088
rect 142448 81023 142768 81024
rect 173168 81088 173488 81089
rect 173168 81024 173176 81088
rect 173240 81024 173256 81088
rect 173320 81024 173336 81088
rect 173400 81024 173416 81088
rect 173480 81024 173488 81088
rect 173168 81023 173488 81024
rect 4208 80544 4528 80545
rect 4208 80480 4216 80544
rect 4280 80480 4296 80544
rect 4360 80480 4376 80544
rect 4440 80480 4456 80544
rect 4520 80480 4528 80544
rect 4208 80479 4528 80480
rect 34928 80544 35248 80545
rect 34928 80480 34936 80544
rect 35000 80480 35016 80544
rect 35080 80480 35096 80544
rect 35160 80480 35176 80544
rect 35240 80480 35248 80544
rect 34928 80479 35248 80480
rect 65648 80544 65968 80545
rect 65648 80480 65656 80544
rect 65720 80480 65736 80544
rect 65800 80480 65816 80544
rect 65880 80480 65896 80544
rect 65960 80480 65968 80544
rect 65648 80479 65968 80480
rect 96368 80544 96688 80545
rect 96368 80480 96376 80544
rect 96440 80480 96456 80544
rect 96520 80480 96536 80544
rect 96600 80480 96616 80544
rect 96680 80480 96688 80544
rect 96368 80479 96688 80480
rect 127088 80544 127408 80545
rect 127088 80480 127096 80544
rect 127160 80480 127176 80544
rect 127240 80480 127256 80544
rect 127320 80480 127336 80544
rect 127400 80480 127408 80544
rect 127088 80479 127408 80480
rect 157808 80544 158128 80545
rect 157808 80480 157816 80544
rect 157880 80480 157896 80544
rect 157960 80480 157976 80544
rect 158040 80480 158056 80544
rect 158120 80480 158128 80544
rect 157808 80479 158128 80480
rect 19568 80000 19888 80001
rect 19568 79936 19576 80000
rect 19640 79936 19656 80000
rect 19720 79936 19736 80000
rect 19800 79936 19816 80000
rect 19880 79936 19888 80000
rect 19568 79935 19888 79936
rect 50288 80000 50608 80001
rect 50288 79936 50296 80000
rect 50360 79936 50376 80000
rect 50440 79936 50456 80000
rect 50520 79936 50536 80000
rect 50600 79936 50608 80000
rect 50288 79935 50608 79936
rect 81008 80000 81328 80001
rect 81008 79936 81016 80000
rect 81080 79936 81096 80000
rect 81160 79936 81176 80000
rect 81240 79936 81256 80000
rect 81320 79936 81328 80000
rect 81008 79935 81328 79936
rect 111728 80000 112048 80001
rect 111728 79936 111736 80000
rect 111800 79936 111816 80000
rect 111880 79936 111896 80000
rect 111960 79936 111976 80000
rect 112040 79936 112048 80000
rect 111728 79935 112048 79936
rect 142448 80000 142768 80001
rect 142448 79936 142456 80000
rect 142520 79936 142536 80000
rect 142600 79936 142616 80000
rect 142680 79936 142696 80000
rect 142760 79936 142768 80000
rect 142448 79935 142768 79936
rect 173168 80000 173488 80001
rect 173168 79936 173176 80000
rect 173240 79936 173256 80000
rect 173320 79936 173336 80000
rect 173400 79936 173416 80000
rect 173480 79936 173488 80000
rect 173168 79935 173488 79936
rect 4208 79456 4528 79457
rect 4208 79392 4216 79456
rect 4280 79392 4296 79456
rect 4360 79392 4376 79456
rect 4440 79392 4456 79456
rect 4520 79392 4528 79456
rect 4208 79391 4528 79392
rect 34928 79456 35248 79457
rect 34928 79392 34936 79456
rect 35000 79392 35016 79456
rect 35080 79392 35096 79456
rect 35160 79392 35176 79456
rect 35240 79392 35248 79456
rect 34928 79391 35248 79392
rect 65648 79456 65968 79457
rect 65648 79392 65656 79456
rect 65720 79392 65736 79456
rect 65800 79392 65816 79456
rect 65880 79392 65896 79456
rect 65960 79392 65968 79456
rect 65648 79391 65968 79392
rect 96368 79456 96688 79457
rect 96368 79392 96376 79456
rect 96440 79392 96456 79456
rect 96520 79392 96536 79456
rect 96600 79392 96616 79456
rect 96680 79392 96688 79456
rect 96368 79391 96688 79392
rect 127088 79456 127408 79457
rect 127088 79392 127096 79456
rect 127160 79392 127176 79456
rect 127240 79392 127256 79456
rect 127320 79392 127336 79456
rect 127400 79392 127408 79456
rect 127088 79391 127408 79392
rect 157808 79456 158128 79457
rect 157808 79392 157816 79456
rect 157880 79392 157896 79456
rect 157960 79392 157976 79456
rect 158040 79392 158056 79456
rect 158120 79392 158128 79456
rect 157808 79391 158128 79392
rect 19568 78912 19888 78913
rect 19568 78848 19576 78912
rect 19640 78848 19656 78912
rect 19720 78848 19736 78912
rect 19800 78848 19816 78912
rect 19880 78848 19888 78912
rect 19568 78847 19888 78848
rect 50288 78912 50608 78913
rect 50288 78848 50296 78912
rect 50360 78848 50376 78912
rect 50440 78848 50456 78912
rect 50520 78848 50536 78912
rect 50600 78848 50608 78912
rect 50288 78847 50608 78848
rect 81008 78912 81328 78913
rect 81008 78848 81016 78912
rect 81080 78848 81096 78912
rect 81160 78848 81176 78912
rect 81240 78848 81256 78912
rect 81320 78848 81328 78912
rect 81008 78847 81328 78848
rect 111728 78912 112048 78913
rect 111728 78848 111736 78912
rect 111800 78848 111816 78912
rect 111880 78848 111896 78912
rect 111960 78848 111976 78912
rect 112040 78848 112048 78912
rect 111728 78847 112048 78848
rect 142448 78912 142768 78913
rect 142448 78848 142456 78912
rect 142520 78848 142536 78912
rect 142600 78848 142616 78912
rect 142680 78848 142696 78912
rect 142760 78848 142768 78912
rect 142448 78847 142768 78848
rect 173168 78912 173488 78913
rect 173168 78848 173176 78912
rect 173240 78848 173256 78912
rect 173320 78848 173336 78912
rect 173400 78848 173416 78912
rect 173480 78848 173488 78912
rect 173168 78847 173488 78848
rect 4208 78368 4528 78369
rect 4208 78304 4216 78368
rect 4280 78304 4296 78368
rect 4360 78304 4376 78368
rect 4440 78304 4456 78368
rect 4520 78304 4528 78368
rect 4208 78303 4528 78304
rect 34928 78368 35248 78369
rect 34928 78304 34936 78368
rect 35000 78304 35016 78368
rect 35080 78304 35096 78368
rect 35160 78304 35176 78368
rect 35240 78304 35248 78368
rect 34928 78303 35248 78304
rect 65648 78368 65968 78369
rect 65648 78304 65656 78368
rect 65720 78304 65736 78368
rect 65800 78304 65816 78368
rect 65880 78304 65896 78368
rect 65960 78304 65968 78368
rect 65648 78303 65968 78304
rect 96368 78368 96688 78369
rect 96368 78304 96376 78368
rect 96440 78304 96456 78368
rect 96520 78304 96536 78368
rect 96600 78304 96616 78368
rect 96680 78304 96688 78368
rect 96368 78303 96688 78304
rect 127088 78368 127408 78369
rect 127088 78304 127096 78368
rect 127160 78304 127176 78368
rect 127240 78304 127256 78368
rect 127320 78304 127336 78368
rect 127400 78304 127408 78368
rect 127088 78303 127408 78304
rect 157808 78368 158128 78369
rect 157808 78304 157816 78368
rect 157880 78304 157896 78368
rect 157960 78304 157976 78368
rect 158040 78304 158056 78368
rect 158120 78304 158128 78368
rect 157808 78303 158128 78304
rect 19568 77824 19888 77825
rect 19568 77760 19576 77824
rect 19640 77760 19656 77824
rect 19720 77760 19736 77824
rect 19800 77760 19816 77824
rect 19880 77760 19888 77824
rect 19568 77759 19888 77760
rect 50288 77824 50608 77825
rect 50288 77760 50296 77824
rect 50360 77760 50376 77824
rect 50440 77760 50456 77824
rect 50520 77760 50536 77824
rect 50600 77760 50608 77824
rect 50288 77759 50608 77760
rect 81008 77824 81328 77825
rect 81008 77760 81016 77824
rect 81080 77760 81096 77824
rect 81160 77760 81176 77824
rect 81240 77760 81256 77824
rect 81320 77760 81328 77824
rect 81008 77759 81328 77760
rect 111728 77824 112048 77825
rect 111728 77760 111736 77824
rect 111800 77760 111816 77824
rect 111880 77760 111896 77824
rect 111960 77760 111976 77824
rect 112040 77760 112048 77824
rect 111728 77759 112048 77760
rect 142448 77824 142768 77825
rect 142448 77760 142456 77824
rect 142520 77760 142536 77824
rect 142600 77760 142616 77824
rect 142680 77760 142696 77824
rect 142760 77760 142768 77824
rect 142448 77759 142768 77760
rect 173168 77824 173488 77825
rect 173168 77760 173176 77824
rect 173240 77760 173256 77824
rect 173320 77760 173336 77824
rect 173400 77760 173416 77824
rect 173480 77760 173488 77824
rect 173168 77759 173488 77760
rect 4208 77280 4528 77281
rect 4208 77216 4216 77280
rect 4280 77216 4296 77280
rect 4360 77216 4376 77280
rect 4440 77216 4456 77280
rect 4520 77216 4528 77280
rect 4208 77215 4528 77216
rect 34928 77280 35248 77281
rect 34928 77216 34936 77280
rect 35000 77216 35016 77280
rect 35080 77216 35096 77280
rect 35160 77216 35176 77280
rect 35240 77216 35248 77280
rect 34928 77215 35248 77216
rect 65648 77280 65968 77281
rect 65648 77216 65656 77280
rect 65720 77216 65736 77280
rect 65800 77216 65816 77280
rect 65880 77216 65896 77280
rect 65960 77216 65968 77280
rect 65648 77215 65968 77216
rect 96368 77280 96688 77281
rect 96368 77216 96376 77280
rect 96440 77216 96456 77280
rect 96520 77216 96536 77280
rect 96600 77216 96616 77280
rect 96680 77216 96688 77280
rect 96368 77215 96688 77216
rect 127088 77280 127408 77281
rect 127088 77216 127096 77280
rect 127160 77216 127176 77280
rect 127240 77216 127256 77280
rect 127320 77216 127336 77280
rect 127400 77216 127408 77280
rect 127088 77215 127408 77216
rect 157808 77280 158128 77281
rect 157808 77216 157816 77280
rect 157880 77216 157896 77280
rect 157960 77216 157976 77280
rect 158040 77216 158056 77280
rect 158120 77216 158128 77280
rect 157808 77215 158128 77216
rect 19568 76736 19888 76737
rect 19568 76672 19576 76736
rect 19640 76672 19656 76736
rect 19720 76672 19736 76736
rect 19800 76672 19816 76736
rect 19880 76672 19888 76736
rect 19568 76671 19888 76672
rect 50288 76736 50608 76737
rect 50288 76672 50296 76736
rect 50360 76672 50376 76736
rect 50440 76672 50456 76736
rect 50520 76672 50536 76736
rect 50600 76672 50608 76736
rect 50288 76671 50608 76672
rect 81008 76736 81328 76737
rect 81008 76672 81016 76736
rect 81080 76672 81096 76736
rect 81160 76672 81176 76736
rect 81240 76672 81256 76736
rect 81320 76672 81328 76736
rect 81008 76671 81328 76672
rect 111728 76736 112048 76737
rect 111728 76672 111736 76736
rect 111800 76672 111816 76736
rect 111880 76672 111896 76736
rect 111960 76672 111976 76736
rect 112040 76672 112048 76736
rect 111728 76671 112048 76672
rect 142448 76736 142768 76737
rect 142448 76672 142456 76736
rect 142520 76672 142536 76736
rect 142600 76672 142616 76736
rect 142680 76672 142696 76736
rect 142760 76672 142768 76736
rect 142448 76671 142768 76672
rect 173168 76736 173488 76737
rect 173168 76672 173176 76736
rect 173240 76672 173256 76736
rect 173320 76672 173336 76736
rect 173400 76672 173416 76736
rect 173480 76672 173488 76736
rect 173168 76671 173488 76672
rect 4208 76192 4528 76193
rect 4208 76128 4216 76192
rect 4280 76128 4296 76192
rect 4360 76128 4376 76192
rect 4440 76128 4456 76192
rect 4520 76128 4528 76192
rect 4208 76127 4528 76128
rect 34928 76192 35248 76193
rect 34928 76128 34936 76192
rect 35000 76128 35016 76192
rect 35080 76128 35096 76192
rect 35160 76128 35176 76192
rect 35240 76128 35248 76192
rect 34928 76127 35248 76128
rect 65648 76192 65968 76193
rect 65648 76128 65656 76192
rect 65720 76128 65736 76192
rect 65800 76128 65816 76192
rect 65880 76128 65896 76192
rect 65960 76128 65968 76192
rect 65648 76127 65968 76128
rect 96368 76192 96688 76193
rect 96368 76128 96376 76192
rect 96440 76128 96456 76192
rect 96520 76128 96536 76192
rect 96600 76128 96616 76192
rect 96680 76128 96688 76192
rect 96368 76127 96688 76128
rect 127088 76192 127408 76193
rect 127088 76128 127096 76192
rect 127160 76128 127176 76192
rect 127240 76128 127256 76192
rect 127320 76128 127336 76192
rect 127400 76128 127408 76192
rect 127088 76127 127408 76128
rect 157808 76192 158128 76193
rect 157808 76128 157816 76192
rect 157880 76128 157896 76192
rect 157960 76128 157976 76192
rect 158040 76128 158056 76192
rect 158120 76128 158128 76192
rect 157808 76127 158128 76128
rect 19568 75648 19888 75649
rect 19568 75584 19576 75648
rect 19640 75584 19656 75648
rect 19720 75584 19736 75648
rect 19800 75584 19816 75648
rect 19880 75584 19888 75648
rect 19568 75583 19888 75584
rect 50288 75648 50608 75649
rect 50288 75584 50296 75648
rect 50360 75584 50376 75648
rect 50440 75584 50456 75648
rect 50520 75584 50536 75648
rect 50600 75584 50608 75648
rect 50288 75583 50608 75584
rect 81008 75648 81328 75649
rect 81008 75584 81016 75648
rect 81080 75584 81096 75648
rect 81160 75584 81176 75648
rect 81240 75584 81256 75648
rect 81320 75584 81328 75648
rect 81008 75583 81328 75584
rect 111728 75648 112048 75649
rect 111728 75584 111736 75648
rect 111800 75584 111816 75648
rect 111880 75584 111896 75648
rect 111960 75584 111976 75648
rect 112040 75584 112048 75648
rect 111728 75583 112048 75584
rect 142448 75648 142768 75649
rect 142448 75584 142456 75648
rect 142520 75584 142536 75648
rect 142600 75584 142616 75648
rect 142680 75584 142696 75648
rect 142760 75584 142768 75648
rect 142448 75583 142768 75584
rect 173168 75648 173488 75649
rect 173168 75584 173176 75648
rect 173240 75584 173256 75648
rect 173320 75584 173336 75648
rect 173400 75584 173416 75648
rect 173480 75584 173488 75648
rect 173168 75583 173488 75584
rect 4208 75104 4528 75105
rect 4208 75040 4216 75104
rect 4280 75040 4296 75104
rect 4360 75040 4376 75104
rect 4440 75040 4456 75104
rect 4520 75040 4528 75104
rect 4208 75039 4528 75040
rect 34928 75104 35248 75105
rect 34928 75040 34936 75104
rect 35000 75040 35016 75104
rect 35080 75040 35096 75104
rect 35160 75040 35176 75104
rect 35240 75040 35248 75104
rect 34928 75039 35248 75040
rect 65648 75104 65968 75105
rect 65648 75040 65656 75104
rect 65720 75040 65736 75104
rect 65800 75040 65816 75104
rect 65880 75040 65896 75104
rect 65960 75040 65968 75104
rect 65648 75039 65968 75040
rect 96368 75104 96688 75105
rect 96368 75040 96376 75104
rect 96440 75040 96456 75104
rect 96520 75040 96536 75104
rect 96600 75040 96616 75104
rect 96680 75040 96688 75104
rect 96368 75039 96688 75040
rect 127088 75104 127408 75105
rect 127088 75040 127096 75104
rect 127160 75040 127176 75104
rect 127240 75040 127256 75104
rect 127320 75040 127336 75104
rect 127400 75040 127408 75104
rect 127088 75039 127408 75040
rect 157808 75104 158128 75105
rect 157808 75040 157816 75104
rect 157880 75040 157896 75104
rect 157960 75040 157976 75104
rect 158040 75040 158056 75104
rect 158120 75040 158128 75104
rect 157808 75039 158128 75040
rect 19568 74560 19888 74561
rect 19568 74496 19576 74560
rect 19640 74496 19656 74560
rect 19720 74496 19736 74560
rect 19800 74496 19816 74560
rect 19880 74496 19888 74560
rect 19568 74495 19888 74496
rect 50288 74560 50608 74561
rect 50288 74496 50296 74560
rect 50360 74496 50376 74560
rect 50440 74496 50456 74560
rect 50520 74496 50536 74560
rect 50600 74496 50608 74560
rect 50288 74495 50608 74496
rect 81008 74560 81328 74561
rect 81008 74496 81016 74560
rect 81080 74496 81096 74560
rect 81160 74496 81176 74560
rect 81240 74496 81256 74560
rect 81320 74496 81328 74560
rect 81008 74495 81328 74496
rect 111728 74560 112048 74561
rect 111728 74496 111736 74560
rect 111800 74496 111816 74560
rect 111880 74496 111896 74560
rect 111960 74496 111976 74560
rect 112040 74496 112048 74560
rect 111728 74495 112048 74496
rect 142448 74560 142768 74561
rect 142448 74496 142456 74560
rect 142520 74496 142536 74560
rect 142600 74496 142616 74560
rect 142680 74496 142696 74560
rect 142760 74496 142768 74560
rect 142448 74495 142768 74496
rect 173168 74560 173488 74561
rect 173168 74496 173176 74560
rect 173240 74496 173256 74560
rect 173320 74496 173336 74560
rect 173400 74496 173416 74560
rect 173480 74496 173488 74560
rect 173168 74495 173488 74496
rect 4208 74016 4528 74017
rect 4208 73952 4216 74016
rect 4280 73952 4296 74016
rect 4360 73952 4376 74016
rect 4440 73952 4456 74016
rect 4520 73952 4528 74016
rect 4208 73951 4528 73952
rect 34928 74016 35248 74017
rect 34928 73952 34936 74016
rect 35000 73952 35016 74016
rect 35080 73952 35096 74016
rect 35160 73952 35176 74016
rect 35240 73952 35248 74016
rect 34928 73951 35248 73952
rect 65648 74016 65968 74017
rect 65648 73952 65656 74016
rect 65720 73952 65736 74016
rect 65800 73952 65816 74016
rect 65880 73952 65896 74016
rect 65960 73952 65968 74016
rect 65648 73951 65968 73952
rect 96368 74016 96688 74017
rect 96368 73952 96376 74016
rect 96440 73952 96456 74016
rect 96520 73952 96536 74016
rect 96600 73952 96616 74016
rect 96680 73952 96688 74016
rect 96368 73951 96688 73952
rect 127088 74016 127408 74017
rect 127088 73952 127096 74016
rect 127160 73952 127176 74016
rect 127240 73952 127256 74016
rect 127320 73952 127336 74016
rect 127400 73952 127408 74016
rect 127088 73951 127408 73952
rect 157808 74016 158128 74017
rect 157808 73952 157816 74016
rect 157880 73952 157896 74016
rect 157960 73952 157976 74016
rect 158040 73952 158056 74016
rect 158120 73952 158128 74016
rect 157808 73951 158128 73952
rect 19568 73472 19888 73473
rect 19568 73408 19576 73472
rect 19640 73408 19656 73472
rect 19720 73408 19736 73472
rect 19800 73408 19816 73472
rect 19880 73408 19888 73472
rect 19568 73407 19888 73408
rect 50288 73472 50608 73473
rect 50288 73408 50296 73472
rect 50360 73408 50376 73472
rect 50440 73408 50456 73472
rect 50520 73408 50536 73472
rect 50600 73408 50608 73472
rect 50288 73407 50608 73408
rect 81008 73472 81328 73473
rect 81008 73408 81016 73472
rect 81080 73408 81096 73472
rect 81160 73408 81176 73472
rect 81240 73408 81256 73472
rect 81320 73408 81328 73472
rect 81008 73407 81328 73408
rect 111728 73472 112048 73473
rect 111728 73408 111736 73472
rect 111800 73408 111816 73472
rect 111880 73408 111896 73472
rect 111960 73408 111976 73472
rect 112040 73408 112048 73472
rect 111728 73407 112048 73408
rect 142448 73472 142768 73473
rect 142448 73408 142456 73472
rect 142520 73408 142536 73472
rect 142600 73408 142616 73472
rect 142680 73408 142696 73472
rect 142760 73408 142768 73472
rect 142448 73407 142768 73408
rect 173168 73472 173488 73473
rect 173168 73408 173176 73472
rect 173240 73408 173256 73472
rect 173320 73408 173336 73472
rect 173400 73408 173416 73472
rect 173480 73408 173488 73472
rect 173168 73407 173488 73408
rect 4208 72928 4528 72929
rect 4208 72864 4216 72928
rect 4280 72864 4296 72928
rect 4360 72864 4376 72928
rect 4440 72864 4456 72928
rect 4520 72864 4528 72928
rect 4208 72863 4528 72864
rect 34928 72928 35248 72929
rect 34928 72864 34936 72928
rect 35000 72864 35016 72928
rect 35080 72864 35096 72928
rect 35160 72864 35176 72928
rect 35240 72864 35248 72928
rect 34928 72863 35248 72864
rect 65648 72928 65968 72929
rect 65648 72864 65656 72928
rect 65720 72864 65736 72928
rect 65800 72864 65816 72928
rect 65880 72864 65896 72928
rect 65960 72864 65968 72928
rect 65648 72863 65968 72864
rect 96368 72928 96688 72929
rect 96368 72864 96376 72928
rect 96440 72864 96456 72928
rect 96520 72864 96536 72928
rect 96600 72864 96616 72928
rect 96680 72864 96688 72928
rect 96368 72863 96688 72864
rect 127088 72928 127408 72929
rect 127088 72864 127096 72928
rect 127160 72864 127176 72928
rect 127240 72864 127256 72928
rect 127320 72864 127336 72928
rect 127400 72864 127408 72928
rect 127088 72863 127408 72864
rect 157808 72928 158128 72929
rect 157808 72864 157816 72928
rect 157880 72864 157896 72928
rect 157960 72864 157976 72928
rect 158040 72864 158056 72928
rect 158120 72864 158128 72928
rect 157808 72863 158128 72864
rect 19568 72384 19888 72385
rect 19568 72320 19576 72384
rect 19640 72320 19656 72384
rect 19720 72320 19736 72384
rect 19800 72320 19816 72384
rect 19880 72320 19888 72384
rect 19568 72319 19888 72320
rect 50288 72384 50608 72385
rect 50288 72320 50296 72384
rect 50360 72320 50376 72384
rect 50440 72320 50456 72384
rect 50520 72320 50536 72384
rect 50600 72320 50608 72384
rect 50288 72319 50608 72320
rect 81008 72384 81328 72385
rect 81008 72320 81016 72384
rect 81080 72320 81096 72384
rect 81160 72320 81176 72384
rect 81240 72320 81256 72384
rect 81320 72320 81328 72384
rect 81008 72319 81328 72320
rect 111728 72384 112048 72385
rect 111728 72320 111736 72384
rect 111800 72320 111816 72384
rect 111880 72320 111896 72384
rect 111960 72320 111976 72384
rect 112040 72320 112048 72384
rect 111728 72319 112048 72320
rect 142448 72384 142768 72385
rect 142448 72320 142456 72384
rect 142520 72320 142536 72384
rect 142600 72320 142616 72384
rect 142680 72320 142696 72384
rect 142760 72320 142768 72384
rect 142448 72319 142768 72320
rect 173168 72384 173488 72385
rect 173168 72320 173176 72384
rect 173240 72320 173256 72384
rect 173320 72320 173336 72384
rect 173400 72320 173416 72384
rect 173480 72320 173488 72384
rect 173168 72319 173488 72320
rect 4208 71840 4528 71841
rect 4208 71776 4216 71840
rect 4280 71776 4296 71840
rect 4360 71776 4376 71840
rect 4440 71776 4456 71840
rect 4520 71776 4528 71840
rect 4208 71775 4528 71776
rect 34928 71840 35248 71841
rect 34928 71776 34936 71840
rect 35000 71776 35016 71840
rect 35080 71776 35096 71840
rect 35160 71776 35176 71840
rect 35240 71776 35248 71840
rect 34928 71775 35248 71776
rect 65648 71840 65968 71841
rect 65648 71776 65656 71840
rect 65720 71776 65736 71840
rect 65800 71776 65816 71840
rect 65880 71776 65896 71840
rect 65960 71776 65968 71840
rect 65648 71775 65968 71776
rect 96368 71840 96688 71841
rect 96368 71776 96376 71840
rect 96440 71776 96456 71840
rect 96520 71776 96536 71840
rect 96600 71776 96616 71840
rect 96680 71776 96688 71840
rect 96368 71775 96688 71776
rect 127088 71840 127408 71841
rect 127088 71776 127096 71840
rect 127160 71776 127176 71840
rect 127240 71776 127256 71840
rect 127320 71776 127336 71840
rect 127400 71776 127408 71840
rect 127088 71775 127408 71776
rect 157808 71840 158128 71841
rect 157808 71776 157816 71840
rect 157880 71776 157896 71840
rect 157960 71776 157976 71840
rect 158040 71776 158056 71840
rect 158120 71776 158128 71840
rect 157808 71775 158128 71776
rect 19568 71296 19888 71297
rect 19568 71232 19576 71296
rect 19640 71232 19656 71296
rect 19720 71232 19736 71296
rect 19800 71232 19816 71296
rect 19880 71232 19888 71296
rect 19568 71231 19888 71232
rect 50288 71296 50608 71297
rect 50288 71232 50296 71296
rect 50360 71232 50376 71296
rect 50440 71232 50456 71296
rect 50520 71232 50536 71296
rect 50600 71232 50608 71296
rect 50288 71231 50608 71232
rect 81008 71296 81328 71297
rect 81008 71232 81016 71296
rect 81080 71232 81096 71296
rect 81160 71232 81176 71296
rect 81240 71232 81256 71296
rect 81320 71232 81328 71296
rect 81008 71231 81328 71232
rect 111728 71296 112048 71297
rect 111728 71232 111736 71296
rect 111800 71232 111816 71296
rect 111880 71232 111896 71296
rect 111960 71232 111976 71296
rect 112040 71232 112048 71296
rect 111728 71231 112048 71232
rect 142448 71296 142768 71297
rect 142448 71232 142456 71296
rect 142520 71232 142536 71296
rect 142600 71232 142616 71296
rect 142680 71232 142696 71296
rect 142760 71232 142768 71296
rect 142448 71231 142768 71232
rect 173168 71296 173488 71297
rect 173168 71232 173176 71296
rect 173240 71232 173256 71296
rect 173320 71232 173336 71296
rect 173400 71232 173416 71296
rect 173480 71232 173488 71296
rect 173168 71231 173488 71232
rect 4208 70752 4528 70753
rect 4208 70688 4216 70752
rect 4280 70688 4296 70752
rect 4360 70688 4376 70752
rect 4440 70688 4456 70752
rect 4520 70688 4528 70752
rect 4208 70687 4528 70688
rect 34928 70752 35248 70753
rect 34928 70688 34936 70752
rect 35000 70688 35016 70752
rect 35080 70688 35096 70752
rect 35160 70688 35176 70752
rect 35240 70688 35248 70752
rect 34928 70687 35248 70688
rect 65648 70752 65968 70753
rect 65648 70688 65656 70752
rect 65720 70688 65736 70752
rect 65800 70688 65816 70752
rect 65880 70688 65896 70752
rect 65960 70688 65968 70752
rect 65648 70687 65968 70688
rect 96368 70752 96688 70753
rect 96368 70688 96376 70752
rect 96440 70688 96456 70752
rect 96520 70688 96536 70752
rect 96600 70688 96616 70752
rect 96680 70688 96688 70752
rect 96368 70687 96688 70688
rect 127088 70752 127408 70753
rect 127088 70688 127096 70752
rect 127160 70688 127176 70752
rect 127240 70688 127256 70752
rect 127320 70688 127336 70752
rect 127400 70688 127408 70752
rect 127088 70687 127408 70688
rect 157808 70752 158128 70753
rect 157808 70688 157816 70752
rect 157880 70688 157896 70752
rect 157960 70688 157976 70752
rect 158040 70688 158056 70752
rect 158120 70688 158128 70752
rect 157808 70687 158128 70688
rect 19568 70208 19888 70209
rect 19568 70144 19576 70208
rect 19640 70144 19656 70208
rect 19720 70144 19736 70208
rect 19800 70144 19816 70208
rect 19880 70144 19888 70208
rect 19568 70143 19888 70144
rect 50288 70208 50608 70209
rect 50288 70144 50296 70208
rect 50360 70144 50376 70208
rect 50440 70144 50456 70208
rect 50520 70144 50536 70208
rect 50600 70144 50608 70208
rect 50288 70143 50608 70144
rect 81008 70208 81328 70209
rect 81008 70144 81016 70208
rect 81080 70144 81096 70208
rect 81160 70144 81176 70208
rect 81240 70144 81256 70208
rect 81320 70144 81328 70208
rect 81008 70143 81328 70144
rect 111728 70208 112048 70209
rect 111728 70144 111736 70208
rect 111800 70144 111816 70208
rect 111880 70144 111896 70208
rect 111960 70144 111976 70208
rect 112040 70144 112048 70208
rect 111728 70143 112048 70144
rect 142448 70208 142768 70209
rect 142448 70144 142456 70208
rect 142520 70144 142536 70208
rect 142600 70144 142616 70208
rect 142680 70144 142696 70208
rect 142760 70144 142768 70208
rect 142448 70143 142768 70144
rect 173168 70208 173488 70209
rect 173168 70144 173176 70208
rect 173240 70144 173256 70208
rect 173320 70144 173336 70208
rect 173400 70144 173416 70208
rect 173480 70144 173488 70208
rect 173168 70143 173488 70144
rect 4208 69664 4528 69665
rect 4208 69600 4216 69664
rect 4280 69600 4296 69664
rect 4360 69600 4376 69664
rect 4440 69600 4456 69664
rect 4520 69600 4528 69664
rect 4208 69599 4528 69600
rect 34928 69664 35248 69665
rect 34928 69600 34936 69664
rect 35000 69600 35016 69664
rect 35080 69600 35096 69664
rect 35160 69600 35176 69664
rect 35240 69600 35248 69664
rect 34928 69599 35248 69600
rect 65648 69664 65968 69665
rect 65648 69600 65656 69664
rect 65720 69600 65736 69664
rect 65800 69600 65816 69664
rect 65880 69600 65896 69664
rect 65960 69600 65968 69664
rect 65648 69599 65968 69600
rect 96368 69664 96688 69665
rect 96368 69600 96376 69664
rect 96440 69600 96456 69664
rect 96520 69600 96536 69664
rect 96600 69600 96616 69664
rect 96680 69600 96688 69664
rect 96368 69599 96688 69600
rect 127088 69664 127408 69665
rect 127088 69600 127096 69664
rect 127160 69600 127176 69664
rect 127240 69600 127256 69664
rect 127320 69600 127336 69664
rect 127400 69600 127408 69664
rect 127088 69599 127408 69600
rect 157808 69664 158128 69665
rect 157808 69600 157816 69664
rect 157880 69600 157896 69664
rect 157960 69600 157976 69664
rect 158040 69600 158056 69664
rect 158120 69600 158128 69664
rect 157808 69599 158128 69600
rect 19568 69120 19888 69121
rect 19568 69056 19576 69120
rect 19640 69056 19656 69120
rect 19720 69056 19736 69120
rect 19800 69056 19816 69120
rect 19880 69056 19888 69120
rect 19568 69055 19888 69056
rect 50288 69120 50608 69121
rect 50288 69056 50296 69120
rect 50360 69056 50376 69120
rect 50440 69056 50456 69120
rect 50520 69056 50536 69120
rect 50600 69056 50608 69120
rect 50288 69055 50608 69056
rect 81008 69120 81328 69121
rect 81008 69056 81016 69120
rect 81080 69056 81096 69120
rect 81160 69056 81176 69120
rect 81240 69056 81256 69120
rect 81320 69056 81328 69120
rect 81008 69055 81328 69056
rect 111728 69120 112048 69121
rect 111728 69056 111736 69120
rect 111800 69056 111816 69120
rect 111880 69056 111896 69120
rect 111960 69056 111976 69120
rect 112040 69056 112048 69120
rect 111728 69055 112048 69056
rect 142448 69120 142768 69121
rect 142448 69056 142456 69120
rect 142520 69056 142536 69120
rect 142600 69056 142616 69120
rect 142680 69056 142696 69120
rect 142760 69056 142768 69120
rect 142448 69055 142768 69056
rect 173168 69120 173488 69121
rect 173168 69056 173176 69120
rect 173240 69056 173256 69120
rect 173320 69056 173336 69120
rect 173400 69056 173416 69120
rect 173480 69056 173488 69120
rect 173168 69055 173488 69056
rect 4208 68576 4528 68577
rect 4208 68512 4216 68576
rect 4280 68512 4296 68576
rect 4360 68512 4376 68576
rect 4440 68512 4456 68576
rect 4520 68512 4528 68576
rect 4208 68511 4528 68512
rect 34928 68576 35248 68577
rect 34928 68512 34936 68576
rect 35000 68512 35016 68576
rect 35080 68512 35096 68576
rect 35160 68512 35176 68576
rect 35240 68512 35248 68576
rect 34928 68511 35248 68512
rect 65648 68576 65968 68577
rect 65648 68512 65656 68576
rect 65720 68512 65736 68576
rect 65800 68512 65816 68576
rect 65880 68512 65896 68576
rect 65960 68512 65968 68576
rect 65648 68511 65968 68512
rect 96368 68576 96688 68577
rect 96368 68512 96376 68576
rect 96440 68512 96456 68576
rect 96520 68512 96536 68576
rect 96600 68512 96616 68576
rect 96680 68512 96688 68576
rect 96368 68511 96688 68512
rect 127088 68576 127408 68577
rect 127088 68512 127096 68576
rect 127160 68512 127176 68576
rect 127240 68512 127256 68576
rect 127320 68512 127336 68576
rect 127400 68512 127408 68576
rect 127088 68511 127408 68512
rect 157808 68576 158128 68577
rect 157808 68512 157816 68576
rect 157880 68512 157896 68576
rect 157960 68512 157976 68576
rect 158040 68512 158056 68576
rect 158120 68512 158128 68576
rect 157808 68511 158128 68512
rect 19568 68032 19888 68033
rect 19568 67968 19576 68032
rect 19640 67968 19656 68032
rect 19720 67968 19736 68032
rect 19800 67968 19816 68032
rect 19880 67968 19888 68032
rect 19568 67967 19888 67968
rect 50288 68032 50608 68033
rect 50288 67968 50296 68032
rect 50360 67968 50376 68032
rect 50440 67968 50456 68032
rect 50520 67968 50536 68032
rect 50600 67968 50608 68032
rect 50288 67967 50608 67968
rect 81008 68032 81328 68033
rect 81008 67968 81016 68032
rect 81080 67968 81096 68032
rect 81160 67968 81176 68032
rect 81240 67968 81256 68032
rect 81320 67968 81328 68032
rect 81008 67967 81328 67968
rect 111728 68032 112048 68033
rect 111728 67968 111736 68032
rect 111800 67968 111816 68032
rect 111880 67968 111896 68032
rect 111960 67968 111976 68032
rect 112040 67968 112048 68032
rect 111728 67967 112048 67968
rect 142448 68032 142768 68033
rect 142448 67968 142456 68032
rect 142520 67968 142536 68032
rect 142600 67968 142616 68032
rect 142680 67968 142696 68032
rect 142760 67968 142768 68032
rect 142448 67967 142768 67968
rect 173168 68032 173488 68033
rect 173168 67968 173176 68032
rect 173240 67968 173256 68032
rect 173320 67968 173336 68032
rect 173400 67968 173416 68032
rect 173480 67968 173488 68032
rect 173168 67967 173488 67968
rect 4208 67488 4528 67489
rect 4208 67424 4216 67488
rect 4280 67424 4296 67488
rect 4360 67424 4376 67488
rect 4440 67424 4456 67488
rect 4520 67424 4528 67488
rect 4208 67423 4528 67424
rect 34928 67488 35248 67489
rect 34928 67424 34936 67488
rect 35000 67424 35016 67488
rect 35080 67424 35096 67488
rect 35160 67424 35176 67488
rect 35240 67424 35248 67488
rect 34928 67423 35248 67424
rect 65648 67488 65968 67489
rect 65648 67424 65656 67488
rect 65720 67424 65736 67488
rect 65800 67424 65816 67488
rect 65880 67424 65896 67488
rect 65960 67424 65968 67488
rect 65648 67423 65968 67424
rect 96368 67488 96688 67489
rect 96368 67424 96376 67488
rect 96440 67424 96456 67488
rect 96520 67424 96536 67488
rect 96600 67424 96616 67488
rect 96680 67424 96688 67488
rect 96368 67423 96688 67424
rect 127088 67488 127408 67489
rect 127088 67424 127096 67488
rect 127160 67424 127176 67488
rect 127240 67424 127256 67488
rect 127320 67424 127336 67488
rect 127400 67424 127408 67488
rect 127088 67423 127408 67424
rect 157808 67488 158128 67489
rect 157808 67424 157816 67488
rect 157880 67424 157896 67488
rect 157960 67424 157976 67488
rect 158040 67424 158056 67488
rect 158120 67424 158128 67488
rect 157808 67423 158128 67424
rect 19568 66944 19888 66945
rect 19568 66880 19576 66944
rect 19640 66880 19656 66944
rect 19720 66880 19736 66944
rect 19800 66880 19816 66944
rect 19880 66880 19888 66944
rect 19568 66879 19888 66880
rect 50288 66944 50608 66945
rect 50288 66880 50296 66944
rect 50360 66880 50376 66944
rect 50440 66880 50456 66944
rect 50520 66880 50536 66944
rect 50600 66880 50608 66944
rect 50288 66879 50608 66880
rect 81008 66944 81328 66945
rect 81008 66880 81016 66944
rect 81080 66880 81096 66944
rect 81160 66880 81176 66944
rect 81240 66880 81256 66944
rect 81320 66880 81328 66944
rect 81008 66879 81328 66880
rect 111728 66944 112048 66945
rect 111728 66880 111736 66944
rect 111800 66880 111816 66944
rect 111880 66880 111896 66944
rect 111960 66880 111976 66944
rect 112040 66880 112048 66944
rect 111728 66879 112048 66880
rect 142448 66944 142768 66945
rect 142448 66880 142456 66944
rect 142520 66880 142536 66944
rect 142600 66880 142616 66944
rect 142680 66880 142696 66944
rect 142760 66880 142768 66944
rect 142448 66879 142768 66880
rect 173168 66944 173488 66945
rect 173168 66880 173176 66944
rect 173240 66880 173256 66944
rect 173320 66880 173336 66944
rect 173400 66880 173416 66944
rect 173480 66880 173488 66944
rect 173168 66879 173488 66880
rect 4208 66400 4528 66401
rect 4208 66336 4216 66400
rect 4280 66336 4296 66400
rect 4360 66336 4376 66400
rect 4440 66336 4456 66400
rect 4520 66336 4528 66400
rect 4208 66335 4528 66336
rect 34928 66400 35248 66401
rect 34928 66336 34936 66400
rect 35000 66336 35016 66400
rect 35080 66336 35096 66400
rect 35160 66336 35176 66400
rect 35240 66336 35248 66400
rect 34928 66335 35248 66336
rect 65648 66400 65968 66401
rect 65648 66336 65656 66400
rect 65720 66336 65736 66400
rect 65800 66336 65816 66400
rect 65880 66336 65896 66400
rect 65960 66336 65968 66400
rect 65648 66335 65968 66336
rect 96368 66400 96688 66401
rect 96368 66336 96376 66400
rect 96440 66336 96456 66400
rect 96520 66336 96536 66400
rect 96600 66336 96616 66400
rect 96680 66336 96688 66400
rect 96368 66335 96688 66336
rect 127088 66400 127408 66401
rect 127088 66336 127096 66400
rect 127160 66336 127176 66400
rect 127240 66336 127256 66400
rect 127320 66336 127336 66400
rect 127400 66336 127408 66400
rect 127088 66335 127408 66336
rect 157808 66400 158128 66401
rect 157808 66336 157816 66400
rect 157880 66336 157896 66400
rect 157960 66336 157976 66400
rect 158040 66336 158056 66400
rect 158120 66336 158128 66400
rect 157808 66335 158128 66336
rect 19568 65856 19888 65857
rect 19568 65792 19576 65856
rect 19640 65792 19656 65856
rect 19720 65792 19736 65856
rect 19800 65792 19816 65856
rect 19880 65792 19888 65856
rect 19568 65791 19888 65792
rect 50288 65856 50608 65857
rect 50288 65792 50296 65856
rect 50360 65792 50376 65856
rect 50440 65792 50456 65856
rect 50520 65792 50536 65856
rect 50600 65792 50608 65856
rect 50288 65791 50608 65792
rect 81008 65856 81328 65857
rect 81008 65792 81016 65856
rect 81080 65792 81096 65856
rect 81160 65792 81176 65856
rect 81240 65792 81256 65856
rect 81320 65792 81328 65856
rect 81008 65791 81328 65792
rect 111728 65856 112048 65857
rect 111728 65792 111736 65856
rect 111800 65792 111816 65856
rect 111880 65792 111896 65856
rect 111960 65792 111976 65856
rect 112040 65792 112048 65856
rect 111728 65791 112048 65792
rect 142448 65856 142768 65857
rect 142448 65792 142456 65856
rect 142520 65792 142536 65856
rect 142600 65792 142616 65856
rect 142680 65792 142696 65856
rect 142760 65792 142768 65856
rect 142448 65791 142768 65792
rect 173168 65856 173488 65857
rect 173168 65792 173176 65856
rect 173240 65792 173256 65856
rect 173320 65792 173336 65856
rect 173400 65792 173416 65856
rect 173480 65792 173488 65856
rect 173168 65791 173488 65792
rect 4208 65312 4528 65313
rect 4208 65248 4216 65312
rect 4280 65248 4296 65312
rect 4360 65248 4376 65312
rect 4440 65248 4456 65312
rect 4520 65248 4528 65312
rect 4208 65247 4528 65248
rect 34928 65312 35248 65313
rect 34928 65248 34936 65312
rect 35000 65248 35016 65312
rect 35080 65248 35096 65312
rect 35160 65248 35176 65312
rect 35240 65248 35248 65312
rect 34928 65247 35248 65248
rect 65648 65312 65968 65313
rect 65648 65248 65656 65312
rect 65720 65248 65736 65312
rect 65800 65248 65816 65312
rect 65880 65248 65896 65312
rect 65960 65248 65968 65312
rect 65648 65247 65968 65248
rect 96368 65312 96688 65313
rect 96368 65248 96376 65312
rect 96440 65248 96456 65312
rect 96520 65248 96536 65312
rect 96600 65248 96616 65312
rect 96680 65248 96688 65312
rect 96368 65247 96688 65248
rect 127088 65312 127408 65313
rect 127088 65248 127096 65312
rect 127160 65248 127176 65312
rect 127240 65248 127256 65312
rect 127320 65248 127336 65312
rect 127400 65248 127408 65312
rect 127088 65247 127408 65248
rect 157808 65312 158128 65313
rect 157808 65248 157816 65312
rect 157880 65248 157896 65312
rect 157960 65248 157976 65312
rect 158040 65248 158056 65312
rect 158120 65248 158128 65312
rect 157808 65247 158128 65248
rect 19568 64768 19888 64769
rect 19568 64704 19576 64768
rect 19640 64704 19656 64768
rect 19720 64704 19736 64768
rect 19800 64704 19816 64768
rect 19880 64704 19888 64768
rect 19568 64703 19888 64704
rect 50288 64768 50608 64769
rect 50288 64704 50296 64768
rect 50360 64704 50376 64768
rect 50440 64704 50456 64768
rect 50520 64704 50536 64768
rect 50600 64704 50608 64768
rect 50288 64703 50608 64704
rect 81008 64768 81328 64769
rect 81008 64704 81016 64768
rect 81080 64704 81096 64768
rect 81160 64704 81176 64768
rect 81240 64704 81256 64768
rect 81320 64704 81328 64768
rect 81008 64703 81328 64704
rect 111728 64768 112048 64769
rect 111728 64704 111736 64768
rect 111800 64704 111816 64768
rect 111880 64704 111896 64768
rect 111960 64704 111976 64768
rect 112040 64704 112048 64768
rect 111728 64703 112048 64704
rect 142448 64768 142768 64769
rect 142448 64704 142456 64768
rect 142520 64704 142536 64768
rect 142600 64704 142616 64768
rect 142680 64704 142696 64768
rect 142760 64704 142768 64768
rect 142448 64703 142768 64704
rect 173168 64768 173488 64769
rect 173168 64704 173176 64768
rect 173240 64704 173256 64768
rect 173320 64704 173336 64768
rect 173400 64704 173416 64768
rect 173480 64704 173488 64768
rect 173168 64703 173488 64704
rect 4208 64224 4528 64225
rect 4208 64160 4216 64224
rect 4280 64160 4296 64224
rect 4360 64160 4376 64224
rect 4440 64160 4456 64224
rect 4520 64160 4528 64224
rect 4208 64159 4528 64160
rect 34928 64224 35248 64225
rect 34928 64160 34936 64224
rect 35000 64160 35016 64224
rect 35080 64160 35096 64224
rect 35160 64160 35176 64224
rect 35240 64160 35248 64224
rect 34928 64159 35248 64160
rect 65648 64224 65968 64225
rect 65648 64160 65656 64224
rect 65720 64160 65736 64224
rect 65800 64160 65816 64224
rect 65880 64160 65896 64224
rect 65960 64160 65968 64224
rect 65648 64159 65968 64160
rect 96368 64224 96688 64225
rect 96368 64160 96376 64224
rect 96440 64160 96456 64224
rect 96520 64160 96536 64224
rect 96600 64160 96616 64224
rect 96680 64160 96688 64224
rect 96368 64159 96688 64160
rect 127088 64224 127408 64225
rect 127088 64160 127096 64224
rect 127160 64160 127176 64224
rect 127240 64160 127256 64224
rect 127320 64160 127336 64224
rect 127400 64160 127408 64224
rect 127088 64159 127408 64160
rect 157808 64224 158128 64225
rect 157808 64160 157816 64224
rect 157880 64160 157896 64224
rect 157960 64160 157976 64224
rect 158040 64160 158056 64224
rect 158120 64160 158128 64224
rect 157808 64159 158128 64160
rect 19568 63680 19888 63681
rect 19568 63616 19576 63680
rect 19640 63616 19656 63680
rect 19720 63616 19736 63680
rect 19800 63616 19816 63680
rect 19880 63616 19888 63680
rect 19568 63615 19888 63616
rect 50288 63680 50608 63681
rect 50288 63616 50296 63680
rect 50360 63616 50376 63680
rect 50440 63616 50456 63680
rect 50520 63616 50536 63680
rect 50600 63616 50608 63680
rect 50288 63615 50608 63616
rect 81008 63680 81328 63681
rect 81008 63616 81016 63680
rect 81080 63616 81096 63680
rect 81160 63616 81176 63680
rect 81240 63616 81256 63680
rect 81320 63616 81328 63680
rect 81008 63615 81328 63616
rect 111728 63680 112048 63681
rect 111728 63616 111736 63680
rect 111800 63616 111816 63680
rect 111880 63616 111896 63680
rect 111960 63616 111976 63680
rect 112040 63616 112048 63680
rect 111728 63615 112048 63616
rect 142448 63680 142768 63681
rect 142448 63616 142456 63680
rect 142520 63616 142536 63680
rect 142600 63616 142616 63680
rect 142680 63616 142696 63680
rect 142760 63616 142768 63680
rect 142448 63615 142768 63616
rect 173168 63680 173488 63681
rect 173168 63616 173176 63680
rect 173240 63616 173256 63680
rect 173320 63616 173336 63680
rect 173400 63616 173416 63680
rect 173480 63616 173488 63680
rect 173168 63615 173488 63616
rect 4208 63136 4528 63137
rect 4208 63072 4216 63136
rect 4280 63072 4296 63136
rect 4360 63072 4376 63136
rect 4440 63072 4456 63136
rect 4520 63072 4528 63136
rect 4208 63071 4528 63072
rect 34928 63136 35248 63137
rect 34928 63072 34936 63136
rect 35000 63072 35016 63136
rect 35080 63072 35096 63136
rect 35160 63072 35176 63136
rect 35240 63072 35248 63136
rect 34928 63071 35248 63072
rect 65648 63136 65968 63137
rect 65648 63072 65656 63136
rect 65720 63072 65736 63136
rect 65800 63072 65816 63136
rect 65880 63072 65896 63136
rect 65960 63072 65968 63136
rect 65648 63071 65968 63072
rect 96368 63136 96688 63137
rect 96368 63072 96376 63136
rect 96440 63072 96456 63136
rect 96520 63072 96536 63136
rect 96600 63072 96616 63136
rect 96680 63072 96688 63136
rect 96368 63071 96688 63072
rect 127088 63136 127408 63137
rect 127088 63072 127096 63136
rect 127160 63072 127176 63136
rect 127240 63072 127256 63136
rect 127320 63072 127336 63136
rect 127400 63072 127408 63136
rect 127088 63071 127408 63072
rect 157808 63136 158128 63137
rect 157808 63072 157816 63136
rect 157880 63072 157896 63136
rect 157960 63072 157976 63136
rect 158040 63072 158056 63136
rect 158120 63072 158128 63136
rect 157808 63071 158128 63072
rect 19568 62592 19888 62593
rect 19568 62528 19576 62592
rect 19640 62528 19656 62592
rect 19720 62528 19736 62592
rect 19800 62528 19816 62592
rect 19880 62528 19888 62592
rect 19568 62527 19888 62528
rect 50288 62592 50608 62593
rect 50288 62528 50296 62592
rect 50360 62528 50376 62592
rect 50440 62528 50456 62592
rect 50520 62528 50536 62592
rect 50600 62528 50608 62592
rect 50288 62527 50608 62528
rect 81008 62592 81328 62593
rect 81008 62528 81016 62592
rect 81080 62528 81096 62592
rect 81160 62528 81176 62592
rect 81240 62528 81256 62592
rect 81320 62528 81328 62592
rect 81008 62527 81328 62528
rect 111728 62592 112048 62593
rect 111728 62528 111736 62592
rect 111800 62528 111816 62592
rect 111880 62528 111896 62592
rect 111960 62528 111976 62592
rect 112040 62528 112048 62592
rect 111728 62527 112048 62528
rect 142448 62592 142768 62593
rect 142448 62528 142456 62592
rect 142520 62528 142536 62592
rect 142600 62528 142616 62592
rect 142680 62528 142696 62592
rect 142760 62528 142768 62592
rect 142448 62527 142768 62528
rect 173168 62592 173488 62593
rect 173168 62528 173176 62592
rect 173240 62528 173256 62592
rect 173320 62528 173336 62592
rect 173400 62528 173416 62592
rect 173480 62528 173488 62592
rect 173168 62527 173488 62528
rect 4208 62048 4528 62049
rect 4208 61984 4216 62048
rect 4280 61984 4296 62048
rect 4360 61984 4376 62048
rect 4440 61984 4456 62048
rect 4520 61984 4528 62048
rect 4208 61983 4528 61984
rect 34928 62048 35248 62049
rect 34928 61984 34936 62048
rect 35000 61984 35016 62048
rect 35080 61984 35096 62048
rect 35160 61984 35176 62048
rect 35240 61984 35248 62048
rect 34928 61983 35248 61984
rect 65648 62048 65968 62049
rect 65648 61984 65656 62048
rect 65720 61984 65736 62048
rect 65800 61984 65816 62048
rect 65880 61984 65896 62048
rect 65960 61984 65968 62048
rect 65648 61983 65968 61984
rect 96368 62048 96688 62049
rect 96368 61984 96376 62048
rect 96440 61984 96456 62048
rect 96520 61984 96536 62048
rect 96600 61984 96616 62048
rect 96680 61984 96688 62048
rect 96368 61983 96688 61984
rect 127088 62048 127408 62049
rect 127088 61984 127096 62048
rect 127160 61984 127176 62048
rect 127240 61984 127256 62048
rect 127320 61984 127336 62048
rect 127400 61984 127408 62048
rect 127088 61983 127408 61984
rect 157808 62048 158128 62049
rect 157808 61984 157816 62048
rect 157880 61984 157896 62048
rect 157960 61984 157976 62048
rect 158040 61984 158056 62048
rect 158120 61984 158128 62048
rect 157808 61983 158128 61984
rect 19568 61504 19888 61505
rect 19568 61440 19576 61504
rect 19640 61440 19656 61504
rect 19720 61440 19736 61504
rect 19800 61440 19816 61504
rect 19880 61440 19888 61504
rect 19568 61439 19888 61440
rect 50288 61504 50608 61505
rect 50288 61440 50296 61504
rect 50360 61440 50376 61504
rect 50440 61440 50456 61504
rect 50520 61440 50536 61504
rect 50600 61440 50608 61504
rect 50288 61439 50608 61440
rect 81008 61504 81328 61505
rect 81008 61440 81016 61504
rect 81080 61440 81096 61504
rect 81160 61440 81176 61504
rect 81240 61440 81256 61504
rect 81320 61440 81328 61504
rect 81008 61439 81328 61440
rect 111728 61504 112048 61505
rect 111728 61440 111736 61504
rect 111800 61440 111816 61504
rect 111880 61440 111896 61504
rect 111960 61440 111976 61504
rect 112040 61440 112048 61504
rect 111728 61439 112048 61440
rect 142448 61504 142768 61505
rect 142448 61440 142456 61504
rect 142520 61440 142536 61504
rect 142600 61440 142616 61504
rect 142680 61440 142696 61504
rect 142760 61440 142768 61504
rect 142448 61439 142768 61440
rect 173168 61504 173488 61505
rect 173168 61440 173176 61504
rect 173240 61440 173256 61504
rect 173320 61440 173336 61504
rect 173400 61440 173416 61504
rect 173480 61440 173488 61504
rect 173168 61439 173488 61440
rect 4208 60960 4528 60961
rect 4208 60896 4216 60960
rect 4280 60896 4296 60960
rect 4360 60896 4376 60960
rect 4440 60896 4456 60960
rect 4520 60896 4528 60960
rect 4208 60895 4528 60896
rect 34928 60960 35248 60961
rect 34928 60896 34936 60960
rect 35000 60896 35016 60960
rect 35080 60896 35096 60960
rect 35160 60896 35176 60960
rect 35240 60896 35248 60960
rect 34928 60895 35248 60896
rect 65648 60960 65968 60961
rect 65648 60896 65656 60960
rect 65720 60896 65736 60960
rect 65800 60896 65816 60960
rect 65880 60896 65896 60960
rect 65960 60896 65968 60960
rect 65648 60895 65968 60896
rect 96368 60960 96688 60961
rect 96368 60896 96376 60960
rect 96440 60896 96456 60960
rect 96520 60896 96536 60960
rect 96600 60896 96616 60960
rect 96680 60896 96688 60960
rect 96368 60895 96688 60896
rect 127088 60960 127408 60961
rect 127088 60896 127096 60960
rect 127160 60896 127176 60960
rect 127240 60896 127256 60960
rect 127320 60896 127336 60960
rect 127400 60896 127408 60960
rect 127088 60895 127408 60896
rect 157808 60960 158128 60961
rect 157808 60896 157816 60960
rect 157880 60896 157896 60960
rect 157960 60896 157976 60960
rect 158040 60896 158056 60960
rect 158120 60896 158128 60960
rect 157808 60895 158128 60896
rect 19568 60416 19888 60417
rect 19568 60352 19576 60416
rect 19640 60352 19656 60416
rect 19720 60352 19736 60416
rect 19800 60352 19816 60416
rect 19880 60352 19888 60416
rect 19568 60351 19888 60352
rect 50288 60416 50608 60417
rect 50288 60352 50296 60416
rect 50360 60352 50376 60416
rect 50440 60352 50456 60416
rect 50520 60352 50536 60416
rect 50600 60352 50608 60416
rect 50288 60351 50608 60352
rect 81008 60416 81328 60417
rect 81008 60352 81016 60416
rect 81080 60352 81096 60416
rect 81160 60352 81176 60416
rect 81240 60352 81256 60416
rect 81320 60352 81328 60416
rect 81008 60351 81328 60352
rect 111728 60416 112048 60417
rect 111728 60352 111736 60416
rect 111800 60352 111816 60416
rect 111880 60352 111896 60416
rect 111960 60352 111976 60416
rect 112040 60352 112048 60416
rect 111728 60351 112048 60352
rect 142448 60416 142768 60417
rect 142448 60352 142456 60416
rect 142520 60352 142536 60416
rect 142600 60352 142616 60416
rect 142680 60352 142696 60416
rect 142760 60352 142768 60416
rect 142448 60351 142768 60352
rect 173168 60416 173488 60417
rect 173168 60352 173176 60416
rect 173240 60352 173256 60416
rect 173320 60352 173336 60416
rect 173400 60352 173416 60416
rect 173480 60352 173488 60416
rect 173168 60351 173488 60352
rect 0 60074 800 60104
rect 2037 60074 2103 60077
rect 0 60072 2103 60074
rect 0 60016 2042 60072
rect 2098 60016 2103 60072
rect 0 60014 2103 60016
rect 0 59984 800 60014
rect 2037 60011 2103 60014
rect 178125 60074 178191 60077
rect 179200 60074 180000 60104
rect 178125 60072 180000 60074
rect 178125 60016 178130 60072
rect 178186 60016 180000 60072
rect 178125 60014 180000 60016
rect 178125 60011 178191 60014
rect 179200 59984 180000 60014
rect 4208 59872 4528 59873
rect 4208 59808 4216 59872
rect 4280 59808 4296 59872
rect 4360 59808 4376 59872
rect 4440 59808 4456 59872
rect 4520 59808 4528 59872
rect 4208 59807 4528 59808
rect 34928 59872 35248 59873
rect 34928 59808 34936 59872
rect 35000 59808 35016 59872
rect 35080 59808 35096 59872
rect 35160 59808 35176 59872
rect 35240 59808 35248 59872
rect 34928 59807 35248 59808
rect 65648 59872 65968 59873
rect 65648 59808 65656 59872
rect 65720 59808 65736 59872
rect 65800 59808 65816 59872
rect 65880 59808 65896 59872
rect 65960 59808 65968 59872
rect 65648 59807 65968 59808
rect 96368 59872 96688 59873
rect 96368 59808 96376 59872
rect 96440 59808 96456 59872
rect 96520 59808 96536 59872
rect 96600 59808 96616 59872
rect 96680 59808 96688 59872
rect 96368 59807 96688 59808
rect 127088 59872 127408 59873
rect 127088 59808 127096 59872
rect 127160 59808 127176 59872
rect 127240 59808 127256 59872
rect 127320 59808 127336 59872
rect 127400 59808 127408 59872
rect 127088 59807 127408 59808
rect 157808 59872 158128 59873
rect 157808 59808 157816 59872
rect 157880 59808 157896 59872
rect 157960 59808 157976 59872
rect 158040 59808 158056 59872
rect 158120 59808 158128 59872
rect 157808 59807 158128 59808
rect 19568 59328 19888 59329
rect 19568 59264 19576 59328
rect 19640 59264 19656 59328
rect 19720 59264 19736 59328
rect 19800 59264 19816 59328
rect 19880 59264 19888 59328
rect 19568 59263 19888 59264
rect 50288 59328 50608 59329
rect 50288 59264 50296 59328
rect 50360 59264 50376 59328
rect 50440 59264 50456 59328
rect 50520 59264 50536 59328
rect 50600 59264 50608 59328
rect 50288 59263 50608 59264
rect 81008 59328 81328 59329
rect 81008 59264 81016 59328
rect 81080 59264 81096 59328
rect 81160 59264 81176 59328
rect 81240 59264 81256 59328
rect 81320 59264 81328 59328
rect 81008 59263 81328 59264
rect 111728 59328 112048 59329
rect 111728 59264 111736 59328
rect 111800 59264 111816 59328
rect 111880 59264 111896 59328
rect 111960 59264 111976 59328
rect 112040 59264 112048 59328
rect 111728 59263 112048 59264
rect 142448 59328 142768 59329
rect 142448 59264 142456 59328
rect 142520 59264 142536 59328
rect 142600 59264 142616 59328
rect 142680 59264 142696 59328
rect 142760 59264 142768 59328
rect 142448 59263 142768 59264
rect 173168 59328 173488 59329
rect 173168 59264 173176 59328
rect 173240 59264 173256 59328
rect 173320 59264 173336 59328
rect 173400 59264 173416 59328
rect 173480 59264 173488 59328
rect 173168 59263 173488 59264
rect 4208 58784 4528 58785
rect 4208 58720 4216 58784
rect 4280 58720 4296 58784
rect 4360 58720 4376 58784
rect 4440 58720 4456 58784
rect 4520 58720 4528 58784
rect 4208 58719 4528 58720
rect 34928 58784 35248 58785
rect 34928 58720 34936 58784
rect 35000 58720 35016 58784
rect 35080 58720 35096 58784
rect 35160 58720 35176 58784
rect 35240 58720 35248 58784
rect 34928 58719 35248 58720
rect 65648 58784 65968 58785
rect 65648 58720 65656 58784
rect 65720 58720 65736 58784
rect 65800 58720 65816 58784
rect 65880 58720 65896 58784
rect 65960 58720 65968 58784
rect 65648 58719 65968 58720
rect 96368 58784 96688 58785
rect 96368 58720 96376 58784
rect 96440 58720 96456 58784
rect 96520 58720 96536 58784
rect 96600 58720 96616 58784
rect 96680 58720 96688 58784
rect 96368 58719 96688 58720
rect 127088 58784 127408 58785
rect 127088 58720 127096 58784
rect 127160 58720 127176 58784
rect 127240 58720 127256 58784
rect 127320 58720 127336 58784
rect 127400 58720 127408 58784
rect 127088 58719 127408 58720
rect 157808 58784 158128 58785
rect 157808 58720 157816 58784
rect 157880 58720 157896 58784
rect 157960 58720 157976 58784
rect 158040 58720 158056 58784
rect 158120 58720 158128 58784
rect 157808 58719 158128 58720
rect 19568 58240 19888 58241
rect 19568 58176 19576 58240
rect 19640 58176 19656 58240
rect 19720 58176 19736 58240
rect 19800 58176 19816 58240
rect 19880 58176 19888 58240
rect 19568 58175 19888 58176
rect 50288 58240 50608 58241
rect 50288 58176 50296 58240
rect 50360 58176 50376 58240
rect 50440 58176 50456 58240
rect 50520 58176 50536 58240
rect 50600 58176 50608 58240
rect 50288 58175 50608 58176
rect 81008 58240 81328 58241
rect 81008 58176 81016 58240
rect 81080 58176 81096 58240
rect 81160 58176 81176 58240
rect 81240 58176 81256 58240
rect 81320 58176 81328 58240
rect 81008 58175 81328 58176
rect 111728 58240 112048 58241
rect 111728 58176 111736 58240
rect 111800 58176 111816 58240
rect 111880 58176 111896 58240
rect 111960 58176 111976 58240
rect 112040 58176 112048 58240
rect 111728 58175 112048 58176
rect 142448 58240 142768 58241
rect 142448 58176 142456 58240
rect 142520 58176 142536 58240
rect 142600 58176 142616 58240
rect 142680 58176 142696 58240
rect 142760 58176 142768 58240
rect 142448 58175 142768 58176
rect 173168 58240 173488 58241
rect 173168 58176 173176 58240
rect 173240 58176 173256 58240
rect 173320 58176 173336 58240
rect 173400 58176 173416 58240
rect 173480 58176 173488 58240
rect 173168 58175 173488 58176
rect 4208 57696 4528 57697
rect 4208 57632 4216 57696
rect 4280 57632 4296 57696
rect 4360 57632 4376 57696
rect 4440 57632 4456 57696
rect 4520 57632 4528 57696
rect 4208 57631 4528 57632
rect 34928 57696 35248 57697
rect 34928 57632 34936 57696
rect 35000 57632 35016 57696
rect 35080 57632 35096 57696
rect 35160 57632 35176 57696
rect 35240 57632 35248 57696
rect 34928 57631 35248 57632
rect 65648 57696 65968 57697
rect 65648 57632 65656 57696
rect 65720 57632 65736 57696
rect 65800 57632 65816 57696
rect 65880 57632 65896 57696
rect 65960 57632 65968 57696
rect 65648 57631 65968 57632
rect 96368 57696 96688 57697
rect 96368 57632 96376 57696
rect 96440 57632 96456 57696
rect 96520 57632 96536 57696
rect 96600 57632 96616 57696
rect 96680 57632 96688 57696
rect 96368 57631 96688 57632
rect 127088 57696 127408 57697
rect 127088 57632 127096 57696
rect 127160 57632 127176 57696
rect 127240 57632 127256 57696
rect 127320 57632 127336 57696
rect 127400 57632 127408 57696
rect 127088 57631 127408 57632
rect 157808 57696 158128 57697
rect 157808 57632 157816 57696
rect 157880 57632 157896 57696
rect 157960 57632 157976 57696
rect 158040 57632 158056 57696
rect 158120 57632 158128 57696
rect 157808 57631 158128 57632
rect 19568 57152 19888 57153
rect 19568 57088 19576 57152
rect 19640 57088 19656 57152
rect 19720 57088 19736 57152
rect 19800 57088 19816 57152
rect 19880 57088 19888 57152
rect 19568 57087 19888 57088
rect 50288 57152 50608 57153
rect 50288 57088 50296 57152
rect 50360 57088 50376 57152
rect 50440 57088 50456 57152
rect 50520 57088 50536 57152
rect 50600 57088 50608 57152
rect 50288 57087 50608 57088
rect 81008 57152 81328 57153
rect 81008 57088 81016 57152
rect 81080 57088 81096 57152
rect 81160 57088 81176 57152
rect 81240 57088 81256 57152
rect 81320 57088 81328 57152
rect 81008 57087 81328 57088
rect 111728 57152 112048 57153
rect 111728 57088 111736 57152
rect 111800 57088 111816 57152
rect 111880 57088 111896 57152
rect 111960 57088 111976 57152
rect 112040 57088 112048 57152
rect 111728 57087 112048 57088
rect 142448 57152 142768 57153
rect 142448 57088 142456 57152
rect 142520 57088 142536 57152
rect 142600 57088 142616 57152
rect 142680 57088 142696 57152
rect 142760 57088 142768 57152
rect 142448 57087 142768 57088
rect 173168 57152 173488 57153
rect 173168 57088 173176 57152
rect 173240 57088 173256 57152
rect 173320 57088 173336 57152
rect 173400 57088 173416 57152
rect 173480 57088 173488 57152
rect 173168 57087 173488 57088
rect 4208 56608 4528 56609
rect 4208 56544 4216 56608
rect 4280 56544 4296 56608
rect 4360 56544 4376 56608
rect 4440 56544 4456 56608
rect 4520 56544 4528 56608
rect 4208 56543 4528 56544
rect 34928 56608 35248 56609
rect 34928 56544 34936 56608
rect 35000 56544 35016 56608
rect 35080 56544 35096 56608
rect 35160 56544 35176 56608
rect 35240 56544 35248 56608
rect 34928 56543 35248 56544
rect 65648 56608 65968 56609
rect 65648 56544 65656 56608
rect 65720 56544 65736 56608
rect 65800 56544 65816 56608
rect 65880 56544 65896 56608
rect 65960 56544 65968 56608
rect 65648 56543 65968 56544
rect 96368 56608 96688 56609
rect 96368 56544 96376 56608
rect 96440 56544 96456 56608
rect 96520 56544 96536 56608
rect 96600 56544 96616 56608
rect 96680 56544 96688 56608
rect 96368 56543 96688 56544
rect 127088 56608 127408 56609
rect 127088 56544 127096 56608
rect 127160 56544 127176 56608
rect 127240 56544 127256 56608
rect 127320 56544 127336 56608
rect 127400 56544 127408 56608
rect 127088 56543 127408 56544
rect 157808 56608 158128 56609
rect 157808 56544 157816 56608
rect 157880 56544 157896 56608
rect 157960 56544 157976 56608
rect 158040 56544 158056 56608
rect 158120 56544 158128 56608
rect 157808 56543 158128 56544
rect 19568 56064 19888 56065
rect 19568 56000 19576 56064
rect 19640 56000 19656 56064
rect 19720 56000 19736 56064
rect 19800 56000 19816 56064
rect 19880 56000 19888 56064
rect 19568 55999 19888 56000
rect 50288 56064 50608 56065
rect 50288 56000 50296 56064
rect 50360 56000 50376 56064
rect 50440 56000 50456 56064
rect 50520 56000 50536 56064
rect 50600 56000 50608 56064
rect 50288 55999 50608 56000
rect 81008 56064 81328 56065
rect 81008 56000 81016 56064
rect 81080 56000 81096 56064
rect 81160 56000 81176 56064
rect 81240 56000 81256 56064
rect 81320 56000 81328 56064
rect 81008 55999 81328 56000
rect 111728 56064 112048 56065
rect 111728 56000 111736 56064
rect 111800 56000 111816 56064
rect 111880 56000 111896 56064
rect 111960 56000 111976 56064
rect 112040 56000 112048 56064
rect 111728 55999 112048 56000
rect 142448 56064 142768 56065
rect 142448 56000 142456 56064
rect 142520 56000 142536 56064
rect 142600 56000 142616 56064
rect 142680 56000 142696 56064
rect 142760 56000 142768 56064
rect 142448 55999 142768 56000
rect 173168 56064 173488 56065
rect 173168 56000 173176 56064
rect 173240 56000 173256 56064
rect 173320 56000 173336 56064
rect 173400 56000 173416 56064
rect 173480 56000 173488 56064
rect 173168 55999 173488 56000
rect 4208 55520 4528 55521
rect 4208 55456 4216 55520
rect 4280 55456 4296 55520
rect 4360 55456 4376 55520
rect 4440 55456 4456 55520
rect 4520 55456 4528 55520
rect 4208 55455 4528 55456
rect 34928 55520 35248 55521
rect 34928 55456 34936 55520
rect 35000 55456 35016 55520
rect 35080 55456 35096 55520
rect 35160 55456 35176 55520
rect 35240 55456 35248 55520
rect 34928 55455 35248 55456
rect 65648 55520 65968 55521
rect 65648 55456 65656 55520
rect 65720 55456 65736 55520
rect 65800 55456 65816 55520
rect 65880 55456 65896 55520
rect 65960 55456 65968 55520
rect 65648 55455 65968 55456
rect 96368 55520 96688 55521
rect 96368 55456 96376 55520
rect 96440 55456 96456 55520
rect 96520 55456 96536 55520
rect 96600 55456 96616 55520
rect 96680 55456 96688 55520
rect 96368 55455 96688 55456
rect 127088 55520 127408 55521
rect 127088 55456 127096 55520
rect 127160 55456 127176 55520
rect 127240 55456 127256 55520
rect 127320 55456 127336 55520
rect 127400 55456 127408 55520
rect 127088 55455 127408 55456
rect 157808 55520 158128 55521
rect 157808 55456 157816 55520
rect 157880 55456 157896 55520
rect 157960 55456 157976 55520
rect 158040 55456 158056 55520
rect 158120 55456 158128 55520
rect 157808 55455 158128 55456
rect 19568 54976 19888 54977
rect 19568 54912 19576 54976
rect 19640 54912 19656 54976
rect 19720 54912 19736 54976
rect 19800 54912 19816 54976
rect 19880 54912 19888 54976
rect 19568 54911 19888 54912
rect 50288 54976 50608 54977
rect 50288 54912 50296 54976
rect 50360 54912 50376 54976
rect 50440 54912 50456 54976
rect 50520 54912 50536 54976
rect 50600 54912 50608 54976
rect 50288 54911 50608 54912
rect 81008 54976 81328 54977
rect 81008 54912 81016 54976
rect 81080 54912 81096 54976
rect 81160 54912 81176 54976
rect 81240 54912 81256 54976
rect 81320 54912 81328 54976
rect 81008 54911 81328 54912
rect 111728 54976 112048 54977
rect 111728 54912 111736 54976
rect 111800 54912 111816 54976
rect 111880 54912 111896 54976
rect 111960 54912 111976 54976
rect 112040 54912 112048 54976
rect 111728 54911 112048 54912
rect 142448 54976 142768 54977
rect 142448 54912 142456 54976
rect 142520 54912 142536 54976
rect 142600 54912 142616 54976
rect 142680 54912 142696 54976
rect 142760 54912 142768 54976
rect 142448 54911 142768 54912
rect 173168 54976 173488 54977
rect 173168 54912 173176 54976
rect 173240 54912 173256 54976
rect 173320 54912 173336 54976
rect 173400 54912 173416 54976
rect 173480 54912 173488 54976
rect 173168 54911 173488 54912
rect 4208 54432 4528 54433
rect 4208 54368 4216 54432
rect 4280 54368 4296 54432
rect 4360 54368 4376 54432
rect 4440 54368 4456 54432
rect 4520 54368 4528 54432
rect 4208 54367 4528 54368
rect 34928 54432 35248 54433
rect 34928 54368 34936 54432
rect 35000 54368 35016 54432
rect 35080 54368 35096 54432
rect 35160 54368 35176 54432
rect 35240 54368 35248 54432
rect 34928 54367 35248 54368
rect 65648 54432 65968 54433
rect 65648 54368 65656 54432
rect 65720 54368 65736 54432
rect 65800 54368 65816 54432
rect 65880 54368 65896 54432
rect 65960 54368 65968 54432
rect 65648 54367 65968 54368
rect 96368 54432 96688 54433
rect 96368 54368 96376 54432
rect 96440 54368 96456 54432
rect 96520 54368 96536 54432
rect 96600 54368 96616 54432
rect 96680 54368 96688 54432
rect 96368 54367 96688 54368
rect 127088 54432 127408 54433
rect 127088 54368 127096 54432
rect 127160 54368 127176 54432
rect 127240 54368 127256 54432
rect 127320 54368 127336 54432
rect 127400 54368 127408 54432
rect 127088 54367 127408 54368
rect 157808 54432 158128 54433
rect 157808 54368 157816 54432
rect 157880 54368 157896 54432
rect 157960 54368 157976 54432
rect 158040 54368 158056 54432
rect 158120 54368 158128 54432
rect 157808 54367 158128 54368
rect 19568 53888 19888 53889
rect 19568 53824 19576 53888
rect 19640 53824 19656 53888
rect 19720 53824 19736 53888
rect 19800 53824 19816 53888
rect 19880 53824 19888 53888
rect 19568 53823 19888 53824
rect 50288 53888 50608 53889
rect 50288 53824 50296 53888
rect 50360 53824 50376 53888
rect 50440 53824 50456 53888
rect 50520 53824 50536 53888
rect 50600 53824 50608 53888
rect 50288 53823 50608 53824
rect 81008 53888 81328 53889
rect 81008 53824 81016 53888
rect 81080 53824 81096 53888
rect 81160 53824 81176 53888
rect 81240 53824 81256 53888
rect 81320 53824 81328 53888
rect 81008 53823 81328 53824
rect 111728 53888 112048 53889
rect 111728 53824 111736 53888
rect 111800 53824 111816 53888
rect 111880 53824 111896 53888
rect 111960 53824 111976 53888
rect 112040 53824 112048 53888
rect 111728 53823 112048 53824
rect 142448 53888 142768 53889
rect 142448 53824 142456 53888
rect 142520 53824 142536 53888
rect 142600 53824 142616 53888
rect 142680 53824 142696 53888
rect 142760 53824 142768 53888
rect 142448 53823 142768 53824
rect 173168 53888 173488 53889
rect 173168 53824 173176 53888
rect 173240 53824 173256 53888
rect 173320 53824 173336 53888
rect 173400 53824 173416 53888
rect 173480 53824 173488 53888
rect 173168 53823 173488 53824
rect 4208 53344 4528 53345
rect 4208 53280 4216 53344
rect 4280 53280 4296 53344
rect 4360 53280 4376 53344
rect 4440 53280 4456 53344
rect 4520 53280 4528 53344
rect 4208 53279 4528 53280
rect 34928 53344 35248 53345
rect 34928 53280 34936 53344
rect 35000 53280 35016 53344
rect 35080 53280 35096 53344
rect 35160 53280 35176 53344
rect 35240 53280 35248 53344
rect 34928 53279 35248 53280
rect 65648 53344 65968 53345
rect 65648 53280 65656 53344
rect 65720 53280 65736 53344
rect 65800 53280 65816 53344
rect 65880 53280 65896 53344
rect 65960 53280 65968 53344
rect 65648 53279 65968 53280
rect 96368 53344 96688 53345
rect 96368 53280 96376 53344
rect 96440 53280 96456 53344
rect 96520 53280 96536 53344
rect 96600 53280 96616 53344
rect 96680 53280 96688 53344
rect 96368 53279 96688 53280
rect 127088 53344 127408 53345
rect 127088 53280 127096 53344
rect 127160 53280 127176 53344
rect 127240 53280 127256 53344
rect 127320 53280 127336 53344
rect 127400 53280 127408 53344
rect 127088 53279 127408 53280
rect 157808 53344 158128 53345
rect 157808 53280 157816 53344
rect 157880 53280 157896 53344
rect 157960 53280 157976 53344
rect 158040 53280 158056 53344
rect 158120 53280 158128 53344
rect 157808 53279 158128 53280
rect 19568 52800 19888 52801
rect 19568 52736 19576 52800
rect 19640 52736 19656 52800
rect 19720 52736 19736 52800
rect 19800 52736 19816 52800
rect 19880 52736 19888 52800
rect 19568 52735 19888 52736
rect 50288 52800 50608 52801
rect 50288 52736 50296 52800
rect 50360 52736 50376 52800
rect 50440 52736 50456 52800
rect 50520 52736 50536 52800
rect 50600 52736 50608 52800
rect 50288 52735 50608 52736
rect 81008 52800 81328 52801
rect 81008 52736 81016 52800
rect 81080 52736 81096 52800
rect 81160 52736 81176 52800
rect 81240 52736 81256 52800
rect 81320 52736 81328 52800
rect 81008 52735 81328 52736
rect 111728 52800 112048 52801
rect 111728 52736 111736 52800
rect 111800 52736 111816 52800
rect 111880 52736 111896 52800
rect 111960 52736 111976 52800
rect 112040 52736 112048 52800
rect 111728 52735 112048 52736
rect 142448 52800 142768 52801
rect 142448 52736 142456 52800
rect 142520 52736 142536 52800
rect 142600 52736 142616 52800
rect 142680 52736 142696 52800
rect 142760 52736 142768 52800
rect 142448 52735 142768 52736
rect 173168 52800 173488 52801
rect 173168 52736 173176 52800
rect 173240 52736 173256 52800
rect 173320 52736 173336 52800
rect 173400 52736 173416 52800
rect 173480 52736 173488 52800
rect 173168 52735 173488 52736
rect 4208 52256 4528 52257
rect 4208 52192 4216 52256
rect 4280 52192 4296 52256
rect 4360 52192 4376 52256
rect 4440 52192 4456 52256
rect 4520 52192 4528 52256
rect 4208 52191 4528 52192
rect 34928 52256 35248 52257
rect 34928 52192 34936 52256
rect 35000 52192 35016 52256
rect 35080 52192 35096 52256
rect 35160 52192 35176 52256
rect 35240 52192 35248 52256
rect 34928 52191 35248 52192
rect 65648 52256 65968 52257
rect 65648 52192 65656 52256
rect 65720 52192 65736 52256
rect 65800 52192 65816 52256
rect 65880 52192 65896 52256
rect 65960 52192 65968 52256
rect 65648 52191 65968 52192
rect 96368 52256 96688 52257
rect 96368 52192 96376 52256
rect 96440 52192 96456 52256
rect 96520 52192 96536 52256
rect 96600 52192 96616 52256
rect 96680 52192 96688 52256
rect 96368 52191 96688 52192
rect 127088 52256 127408 52257
rect 127088 52192 127096 52256
rect 127160 52192 127176 52256
rect 127240 52192 127256 52256
rect 127320 52192 127336 52256
rect 127400 52192 127408 52256
rect 127088 52191 127408 52192
rect 157808 52256 158128 52257
rect 157808 52192 157816 52256
rect 157880 52192 157896 52256
rect 157960 52192 157976 52256
rect 158040 52192 158056 52256
rect 158120 52192 158128 52256
rect 157808 52191 158128 52192
rect 19568 51712 19888 51713
rect 19568 51648 19576 51712
rect 19640 51648 19656 51712
rect 19720 51648 19736 51712
rect 19800 51648 19816 51712
rect 19880 51648 19888 51712
rect 19568 51647 19888 51648
rect 50288 51712 50608 51713
rect 50288 51648 50296 51712
rect 50360 51648 50376 51712
rect 50440 51648 50456 51712
rect 50520 51648 50536 51712
rect 50600 51648 50608 51712
rect 50288 51647 50608 51648
rect 81008 51712 81328 51713
rect 81008 51648 81016 51712
rect 81080 51648 81096 51712
rect 81160 51648 81176 51712
rect 81240 51648 81256 51712
rect 81320 51648 81328 51712
rect 81008 51647 81328 51648
rect 111728 51712 112048 51713
rect 111728 51648 111736 51712
rect 111800 51648 111816 51712
rect 111880 51648 111896 51712
rect 111960 51648 111976 51712
rect 112040 51648 112048 51712
rect 111728 51647 112048 51648
rect 142448 51712 142768 51713
rect 142448 51648 142456 51712
rect 142520 51648 142536 51712
rect 142600 51648 142616 51712
rect 142680 51648 142696 51712
rect 142760 51648 142768 51712
rect 142448 51647 142768 51648
rect 173168 51712 173488 51713
rect 173168 51648 173176 51712
rect 173240 51648 173256 51712
rect 173320 51648 173336 51712
rect 173400 51648 173416 51712
rect 173480 51648 173488 51712
rect 173168 51647 173488 51648
rect 4208 51168 4528 51169
rect 4208 51104 4216 51168
rect 4280 51104 4296 51168
rect 4360 51104 4376 51168
rect 4440 51104 4456 51168
rect 4520 51104 4528 51168
rect 4208 51103 4528 51104
rect 34928 51168 35248 51169
rect 34928 51104 34936 51168
rect 35000 51104 35016 51168
rect 35080 51104 35096 51168
rect 35160 51104 35176 51168
rect 35240 51104 35248 51168
rect 34928 51103 35248 51104
rect 65648 51168 65968 51169
rect 65648 51104 65656 51168
rect 65720 51104 65736 51168
rect 65800 51104 65816 51168
rect 65880 51104 65896 51168
rect 65960 51104 65968 51168
rect 65648 51103 65968 51104
rect 96368 51168 96688 51169
rect 96368 51104 96376 51168
rect 96440 51104 96456 51168
rect 96520 51104 96536 51168
rect 96600 51104 96616 51168
rect 96680 51104 96688 51168
rect 96368 51103 96688 51104
rect 127088 51168 127408 51169
rect 127088 51104 127096 51168
rect 127160 51104 127176 51168
rect 127240 51104 127256 51168
rect 127320 51104 127336 51168
rect 127400 51104 127408 51168
rect 127088 51103 127408 51104
rect 157808 51168 158128 51169
rect 157808 51104 157816 51168
rect 157880 51104 157896 51168
rect 157960 51104 157976 51168
rect 158040 51104 158056 51168
rect 158120 51104 158128 51168
rect 157808 51103 158128 51104
rect 19568 50624 19888 50625
rect 19568 50560 19576 50624
rect 19640 50560 19656 50624
rect 19720 50560 19736 50624
rect 19800 50560 19816 50624
rect 19880 50560 19888 50624
rect 19568 50559 19888 50560
rect 50288 50624 50608 50625
rect 50288 50560 50296 50624
rect 50360 50560 50376 50624
rect 50440 50560 50456 50624
rect 50520 50560 50536 50624
rect 50600 50560 50608 50624
rect 50288 50559 50608 50560
rect 81008 50624 81328 50625
rect 81008 50560 81016 50624
rect 81080 50560 81096 50624
rect 81160 50560 81176 50624
rect 81240 50560 81256 50624
rect 81320 50560 81328 50624
rect 81008 50559 81328 50560
rect 111728 50624 112048 50625
rect 111728 50560 111736 50624
rect 111800 50560 111816 50624
rect 111880 50560 111896 50624
rect 111960 50560 111976 50624
rect 112040 50560 112048 50624
rect 111728 50559 112048 50560
rect 142448 50624 142768 50625
rect 142448 50560 142456 50624
rect 142520 50560 142536 50624
rect 142600 50560 142616 50624
rect 142680 50560 142696 50624
rect 142760 50560 142768 50624
rect 142448 50559 142768 50560
rect 173168 50624 173488 50625
rect 173168 50560 173176 50624
rect 173240 50560 173256 50624
rect 173320 50560 173336 50624
rect 173400 50560 173416 50624
rect 173480 50560 173488 50624
rect 173168 50559 173488 50560
rect 4208 50080 4528 50081
rect 4208 50016 4216 50080
rect 4280 50016 4296 50080
rect 4360 50016 4376 50080
rect 4440 50016 4456 50080
rect 4520 50016 4528 50080
rect 4208 50015 4528 50016
rect 34928 50080 35248 50081
rect 34928 50016 34936 50080
rect 35000 50016 35016 50080
rect 35080 50016 35096 50080
rect 35160 50016 35176 50080
rect 35240 50016 35248 50080
rect 34928 50015 35248 50016
rect 65648 50080 65968 50081
rect 65648 50016 65656 50080
rect 65720 50016 65736 50080
rect 65800 50016 65816 50080
rect 65880 50016 65896 50080
rect 65960 50016 65968 50080
rect 65648 50015 65968 50016
rect 96368 50080 96688 50081
rect 96368 50016 96376 50080
rect 96440 50016 96456 50080
rect 96520 50016 96536 50080
rect 96600 50016 96616 50080
rect 96680 50016 96688 50080
rect 96368 50015 96688 50016
rect 127088 50080 127408 50081
rect 127088 50016 127096 50080
rect 127160 50016 127176 50080
rect 127240 50016 127256 50080
rect 127320 50016 127336 50080
rect 127400 50016 127408 50080
rect 127088 50015 127408 50016
rect 157808 50080 158128 50081
rect 157808 50016 157816 50080
rect 157880 50016 157896 50080
rect 157960 50016 157976 50080
rect 158040 50016 158056 50080
rect 158120 50016 158128 50080
rect 157808 50015 158128 50016
rect 19568 49536 19888 49537
rect 19568 49472 19576 49536
rect 19640 49472 19656 49536
rect 19720 49472 19736 49536
rect 19800 49472 19816 49536
rect 19880 49472 19888 49536
rect 19568 49471 19888 49472
rect 50288 49536 50608 49537
rect 50288 49472 50296 49536
rect 50360 49472 50376 49536
rect 50440 49472 50456 49536
rect 50520 49472 50536 49536
rect 50600 49472 50608 49536
rect 50288 49471 50608 49472
rect 81008 49536 81328 49537
rect 81008 49472 81016 49536
rect 81080 49472 81096 49536
rect 81160 49472 81176 49536
rect 81240 49472 81256 49536
rect 81320 49472 81328 49536
rect 81008 49471 81328 49472
rect 111728 49536 112048 49537
rect 111728 49472 111736 49536
rect 111800 49472 111816 49536
rect 111880 49472 111896 49536
rect 111960 49472 111976 49536
rect 112040 49472 112048 49536
rect 111728 49471 112048 49472
rect 142448 49536 142768 49537
rect 142448 49472 142456 49536
rect 142520 49472 142536 49536
rect 142600 49472 142616 49536
rect 142680 49472 142696 49536
rect 142760 49472 142768 49536
rect 142448 49471 142768 49472
rect 173168 49536 173488 49537
rect 173168 49472 173176 49536
rect 173240 49472 173256 49536
rect 173320 49472 173336 49536
rect 173400 49472 173416 49536
rect 173480 49472 173488 49536
rect 173168 49471 173488 49472
rect 4208 48992 4528 48993
rect 4208 48928 4216 48992
rect 4280 48928 4296 48992
rect 4360 48928 4376 48992
rect 4440 48928 4456 48992
rect 4520 48928 4528 48992
rect 4208 48927 4528 48928
rect 34928 48992 35248 48993
rect 34928 48928 34936 48992
rect 35000 48928 35016 48992
rect 35080 48928 35096 48992
rect 35160 48928 35176 48992
rect 35240 48928 35248 48992
rect 34928 48927 35248 48928
rect 65648 48992 65968 48993
rect 65648 48928 65656 48992
rect 65720 48928 65736 48992
rect 65800 48928 65816 48992
rect 65880 48928 65896 48992
rect 65960 48928 65968 48992
rect 65648 48927 65968 48928
rect 96368 48992 96688 48993
rect 96368 48928 96376 48992
rect 96440 48928 96456 48992
rect 96520 48928 96536 48992
rect 96600 48928 96616 48992
rect 96680 48928 96688 48992
rect 96368 48927 96688 48928
rect 127088 48992 127408 48993
rect 127088 48928 127096 48992
rect 127160 48928 127176 48992
rect 127240 48928 127256 48992
rect 127320 48928 127336 48992
rect 127400 48928 127408 48992
rect 127088 48927 127408 48928
rect 157808 48992 158128 48993
rect 157808 48928 157816 48992
rect 157880 48928 157896 48992
rect 157960 48928 157976 48992
rect 158040 48928 158056 48992
rect 158120 48928 158128 48992
rect 157808 48927 158128 48928
rect 19568 48448 19888 48449
rect 19568 48384 19576 48448
rect 19640 48384 19656 48448
rect 19720 48384 19736 48448
rect 19800 48384 19816 48448
rect 19880 48384 19888 48448
rect 19568 48383 19888 48384
rect 50288 48448 50608 48449
rect 50288 48384 50296 48448
rect 50360 48384 50376 48448
rect 50440 48384 50456 48448
rect 50520 48384 50536 48448
rect 50600 48384 50608 48448
rect 50288 48383 50608 48384
rect 81008 48448 81328 48449
rect 81008 48384 81016 48448
rect 81080 48384 81096 48448
rect 81160 48384 81176 48448
rect 81240 48384 81256 48448
rect 81320 48384 81328 48448
rect 81008 48383 81328 48384
rect 111728 48448 112048 48449
rect 111728 48384 111736 48448
rect 111800 48384 111816 48448
rect 111880 48384 111896 48448
rect 111960 48384 111976 48448
rect 112040 48384 112048 48448
rect 111728 48383 112048 48384
rect 142448 48448 142768 48449
rect 142448 48384 142456 48448
rect 142520 48384 142536 48448
rect 142600 48384 142616 48448
rect 142680 48384 142696 48448
rect 142760 48384 142768 48448
rect 142448 48383 142768 48384
rect 173168 48448 173488 48449
rect 173168 48384 173176 48448
rect 173240 48384 173256 48448
rect 173320 48384 173336 48448
rect 173400 48384 173416 48448
rect 173480 48384 173488 48448
rect 173168 48383 173488 48384
rect 4208 47904 4528 47905
rect 4208 47840 4216 47904
rect 4280 47840 4296 47904
rect 4360 47840 4376 47904
rect 4440 47840 4456 47904
rect 4520 47840 4528 47904
rect 4208 47839 4528 47840
rect 34928 47904 35248 47905
rect 34928 47840 34936 47904
rect 35000 47840 35016 47904
rect 35080 47840 35096 47904
rect 35160 47840 35176 47904
rect 35240 47840 35248 47904
rect 34928 47839 35248 47840
rect 65648 47904 65968 47905
rect 65648 47840 65656 47904
rect 65720 47840 65736 47904
rect 65800 47840 65816 47904
rect 65880 47840 65896 47904
rect 65960 47840 65968 47904
rect 65648 47839 65968 47840
rect 96368 47904 96688 47905
rect 96368 47840 96376 47904
rect 96440 47840 96456 47904
rect 96520 47840 96536 47904
rect 96600 47840 96616 47904
rect 96680 47840 96688 47904
rect 96368 47839 96688 47840
rect 127088 47904 127408 47905
rect 127088 47840 127096 47904
rect 127160 47840 127176 47904
rect 127240 47840 127256 47904
rect 127320 47840 127336 47904
rect 127400 47840 127408 47904
rect 127088 47839 127408 47840
rect 157808 47904 158128 47905
rect 157808 47840 157816 47904
rect 157880 47840 157896 47904
rect 157960 47840 157976 47904
rect 158040 47840 158056 47904
rect 158120 47840 158128 47904
rect 157808 47839 158128 47840
rect 19568 47360 19888 47361
rect 19568 47296 19576 47360
rect 19640 47296 19656 47360
rect 19720 47296 19736 47360
rect 19800 47296 19816 47360
rect 19880 47296 19888 47360
rect 19568 47295 19888 47296
rect 50288 47360 50608 47361
rect 50288 47296 50296 47360
rect 50360 47296 50376 47360
rect 50440 47296 50456 47360
rect 50520 47296 50536 47360
rect 50600 47296 50608 47360
rect 50288 47295 50608 47296
rect 81008 47360 81328 47361
rect 81008 47296 81016 47360
rect 81080 47296 81096 47360
rect 81160 47296 81176 47360
rect 81240 47296 81256 47360
rect 81320 47296 81328 47360
rect 81008 47295 81328 47296
rect 111728 47360 112048 47361
rect 111728 47296 111736 47360
rect 111800 47296 111816 47360
rect 111880 47296 111896 47360
rect 111960 47296 111976 47360
rect 112040 47296 112048 47360
rect 111728 47295 112048 47296
rect 142448 47360 142768 47361
rect 142448 47296 142456 47360
rect 142520 47296 142536 47360
rect 142600 47296 142616 47360
rect 142680 47296 142696 47360
rect 142760 47296 142768 47360
rect 142448 47295 142768 47296
rect 173168 47360 173488 47361
rect 173168 47296 173176 47360
rect 173240 47296 173256 47360
rect 173320 47296 173336 47360
rect 173400 47296 173416 47360
rect 173480 47296 173488 47360
rect 173168 47295 173488 47296
rect 4208 46816 4528 46817
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 46751 4528 46752
rect 34928 46816 35248 46817
rect 34928 46752 34936 46816
rect 35000 46752 35016 46816
rect 35080 46752 35096 46816
rect 35160 46752 35176 46816
rect 35240 46752 35248 46816
rect 34928 46751 35248 46752
rect 65648 46816 65968 46817
rect 65648 46752 65656 46816
rect 65720 46752 65736 46816
rect 65800 46752 65816 46816
rect 65880 46752 65896 46816
rect 65960 46752 65968 46816
rect 65648 46751 65968 46752
rect 96368 46816 96688 46817
rect 96368 46752 96376 46816
rect 96440 46752 96456 46816
rect 96520 46752 96536 46816
rect 96600 46752 96616 46816
rect 96680 46752 96688 46816
rect 96368 46751 96688 46752
rect 127088 46816 127408 46817
rect 127088 46752 127096 46816
rect 127160 46752 127176 46816
rect 127240 46752 127256 46816
rect 127320 46752 127336 46816
rect 127400 46752 127408 46816
rect 127088 46751 127408 46752
rect 157808 46816 158128 46817
rect 157808 46752 157816 46816
rect 157880 46752 157896 46816
rect 157960 46752 157976 46816
rect 158040 46752 158056 46816
rect 158120 46752 158128 46816
rect 157808 46751 158128 46752
rect 19568 46272 19888 46273
rect 19568 46208 19576 46272
rect 19640 46208 19656 46272
rect 19720 46208 19736 46272
rect 19800 46208 19816 46272
rect 19880 46208 19888 46272
rect 19568 46207 19888 46208
rect 50288 46272 50608 46273
rect 50288 46208 50296 46272
rect 50360 46208 50376 46272
rect 50440 46208 50456 46272
rect 50520 46208 50536 46272
rect 50600 46208 50608 46272
rect 50288 46207 50608 46208
rect 81008 46272 81328 46273
rect 81008 46208 81016 46272
rect 81080 46208 81096 46272
rect 81160 46208 81176 46272
rect 81240 46208 81256 46272
rect 81320 46208 81328 46272
rect 81008 46207 81328 46208
rect 111728 46272 112048 46273
rect 111728 46208 111736 46272
rect 111800 46208 111816 46272
rect 111880 46208 111896 46272
rect 111960 46208 111976 46272
rect 112040 46208 112048 46272
rect 111728 46207 112048 46208
rect 142448 46272 142768 46273
rect 142448 46208 142456 46272
rect 142520 46208 142536 46272
rect 142600 46208 142616 46272
rect 142680 46208 142696 46272
rect 142760 46208 142768 46272
rect 142448 46207 142768 46208
rect 173168 46272 173488 46273
rect 173168 46208 173176 46272
rect 173240 46208 173256 46272
rect 173320 46208 173336 46272
rect 173400 46208 173416 46272
rect 173480 46208 173488 46272
rect 173168 46207 173488 46208
rect 4208 45728 4528 45729
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 45663 4528 45664
rect 34928 45728 35248 45729
rect 34928 45664 34936 45728
rect 35000 45664 35016 45728
rect 35080 45664 35096 45728
rect 35160 45664 35176 45728
rect 35240 45664 35248 45728
rect 34928 45663 35248 45664
rect 65648 45728 65968 45729
rect 65648 45664 65656 45728
rect 65720 45664 65736 45728
rect 65800 45664 65816 45728
rect 65880 45664 65896 45728
rect 65960 45664 65968 45728
rect 65648 45663 65968 45664
rect 96368 45728 96688 45729
rect 96368 45664 96376 45728
rect 96440 45664 96456 45728
rect 96520 45664 96536 45728
rect 96600 45664 96616 45728
rect 96680 45664 96688 45728
rect 96368 45663 96688 45664
rect 127088 45728 127408 45729
rect 127088 45664 127096 45728
rect 127160 45664 127176 45728
rect 127240 45664 127256 45728
rect 127320 45664 127336 45728
rect 127400 45664 127408 45728
rect 127088 45663 127408 45664
rect 157808 45728 158128 45729
rect 157808 45664 157816 45728
rect 157880 45664 157896 45728
rect 157960 45664 157976 45728
rect 158040 45664 158056 45728
rect 158120 45664 158128 45728
rect 157808 45663 158128 45664
rect 19568 45184 19888 45185
rect 19568 45120 19576 45184
rect 19640 45120 19656 45184
rect 19720 45120 19736 45184
rect 19800 45120 19816 45184
rect 19880 45120 19888 45184
rect 19568 45119 19888 45120
rect 50288 45184 50608 45185
rect 50288 45120 50296 45184
rect 50360 45120 50376 45184
rect 50440 45120 50456 45184
rect 50520 45120 50536 45184
rect 50600 45120 50608 45184
rect 50288 45119 50608 45120
rect 81008 45184 81328 45185
rect 81008 45120 81016 45184
rect 81080 45120 81096 45184
rect 81160 45120 81176 45184
rect 81240 45120 81256 45184
rect 81320 45120 81328 45184
rect 81008 45119 81328 45120
rect 111728 45184 112048 45185
rect 111728 45120 111736 45184
rect 111800 45120 111816 45184
rect 111880 45120 111896 45184
rect 111960 45120 111976 45184
rect 112040 45120 112048 45184
rect 111728 45119 112048 45120
rect 142448 45184 142768 45185
rect 142448 45120 142456 45184
rect 142520 45120 142536 45184
rect 142600 45120 142616 45184
rect 142680 45120 142696 45184
rect 142760 45120 142768 45184
rect 142448 45119 142768 45120
rect 173168 45184 173488 45185
rect 173168 45120 173176 45184
rect 173240 45120 173256 45184
rect 173320 45120 173336 45184
rect 173400 45120 173416 45184
rect 173480 45120 173488 45184
rect 173168 45119 173488 45120
rect 4208 44640 4528 44641
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 44575 4528 44576
rect 34928 44640 35248 44641
rect 34928 44576 34936 44640
rect 35000 44576 35016 44640
rect 35080 44576 35096 44640
rect 35160 44576 35176 44640
rect 35240 44576 35248 44640
rect 34928 44575 35248 44576
rect 65648 44640 65968 44641
rect 65648 44576 65656 44640
rect 65720 44576 65736 44640
rect 65800 44576 65816 44640
rect 65880 44576 65896 44640
rect 65960 44576 65968 44640
rect 65648 44575 65968 44576
rect 96368 44640 96688 44641
rect 96368 44576 96376 44640
rect 96440 44576 96456 44640
rect 96520 44576 96536 44640
rect 96600 44576 96616 44640
rect 96680 44576 96688 44640
rect 96368 44575 96688 44576
rect 127088 44640 127408 44641
rect 127088 44576 127096 44640
rect 127160 44576 127176 44640
rect 127240 44576 127256 44640
rect 127320 44576 127336 44640
rect 127400 44576 127408 44640
rect 127088 44575 127408 44576
rect 157808 44640 158128 44641
rect 157808 44576 157816 44640
rect 157880 44576 157896 44640
rect 157960 44576 157976 44640
rect 158040 44576 158056 44640
rect 158120 44576 158128 44640
rect 157808 44575 158128 44576
rect 19568 44096 19888 44097
rect 19568 44032 19576 44096
rect 19640 44032 19656 44096
rect 19720 44032 19736 44096
rect 19800 44032 19816 44096
rect 19880 44032 19888 44096
rect 19568 44031 19888 44032
rect 50288 44096 50608 44097
rect 50288 44032 50296 44096
rect 50360 44032 50376 44096
rect 50440 44032 50456 44096
rect 50520 44032 50536 44096
rect 50600 44032 50608 44096
rect 50288 44031 50608 44032
rect 81008 44096 81328 44097
rect 81008 44032 81016 44096
rect 81080 44032 81096 44096
rect 81160 44032 81176 44096
rect 81240 44032 81256 44096
rect 81320 44032 81328 44096
rect 81008 44031 81328 44032
rect 111728 44096 112048 44097
rect 111728 44032 111736 44096
rect 111800 44032 111816 44096
rect 111880 44032 111896 44096
rect 111960 44032 111976 44096
rect 112040 44032 112048 44096
rect 111728 44031 112048 44032
rect 142448 44096 142768 44097
rect 142448 44032 142456 44096
rect 142520 44032 142536 44096
rect 142600 44032 142616 44096
rect 142680 44032 142696 44096
rect 142760 44032 142768 44096
rect 142448 44031 142768 44032
rect 173168 44096 173488 44097
rect 173168 44032 173176 44096
rect 173240 44032 173256 44096
rect 173320 44032 173336 44096
rect 173400 44032 173416 44096
rect 173480 44032 173488 44096
rect 173168 44031 173488 44032
rect 4208 43552 4528 43553
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 43487 4528 43488
rect 34928 43552 35248 43553
rect 34928 43488 34936 43552
rect 35000 43488 35016 43552
rect 35080 43488 35096 43552
rect 35160 43488 35176 43552
rect 35240 43488 35248 43552
rect 34928 43487 35248 43488
rect 65648 43552 65968 43553
rect 65648 43488 65656 43552
rect 65720 43488 65736 43552
rect 65800 43488 65816 43552
rect 65880 43488 65896 43552
rect 65960 43488 65968 43552
rect 65648 43487 65968 43488
rect 96368 43552 96688 43553
rect 96368 43488 96376 43552
rect 96440 43488 96456 43552
rect 96520 43488 96536 43552
rect 96600 43488 96616 43552
rect 96680 43488 96688 43552
rect 96368 43487 96688 43488
rect 127088 43552 127408 43553
rect 127088 43488 127096 43552
rect 127160 43488 127176 43552
rect 127240 43488 127256 43552
rect 127320 43488 127336 43552
rect 127400 43488 127408 43552
rect 127088 43487 127408 43488
rect 157808 43552 158128 43553
rect 157808 43488 157816 43552
rect 157880 43488 157896 43552
rect 157960 43488 157976 43552
rect 158040 43488 158056 43552
rect 158120 43488 158128 43552
rect 157808 43487 158128 43488
rect 19568 43008 19888 43009
rect 19568 42944 19576 43008
rect 19640 42944 19656 43008
rect 19720 42944 19736 43008
rect 19800 42944 19816 43008
rect 19880 42944 19888 43008
rect 19568 42943 19888 42944
rect 50288 43008 50608 43009
rect 50288 42944 50296 43008
rect 50360 42944 50376 43008
rect 50440 42944 50456 43008
rect 50520 42944 50536 43008
rect 50600 42944 50608 43008
rect 50288 42943 50608 42944
rect 81008 43008 81328 43009
rect 81008 42944 81016 43008
rect 81080 42944 81096 43008
rect 81160 42944 81176 43008
rect 81240 42944 81256 43008
rect 81320 42944 81328 43008
rect 81008 42943 81328 42944
rect 111728 43008 112048 43009
rect 111728 42944 111736 43008
rect 111800 42944 111816 43008
rect 111880 42944 111896 43008
rect 111960 42944 111976 43008
rect 112040 42944 112048 43008
rect 111728 42943 112048 42944
rect 142448 43008 142768 43009
rect 142448 42944 142456 43008
rect 142520 42944 142536 43008
rect 142600 42944 142616 43008
rect 142680 42944 142696 43008
rect 142760 42944 142768 43008
rect 142448 42943 142768 42944
rect 173168 43008 173488 43009
rect 173168 42944 173176 43008
rect 173240 42944 173256 43008
rect 173320 42944 173336 43008
rect 173400 42944 173416 43008
rect 173480 42944 173488 43008
rect 173168 42943 173488 42944
rect 4208 42464 4528 42465
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 42399 4528 42400
rect 34928 42464 35248 42465
rect 34928 42400 34936 42464
rect 35000 42400 35016 42464
rect 35080 42400 35096 42464
rect 35160 42400 35176 42464
rect 35240 42400 35248 42464
rect 34928 42399 35248 42400
rect 65648 42464 65968 42465
rect 65648 42400 65656 42464
rect 65720 42400 65736 42464
rect 65800 42400 65816 42464
rect 65880 42400 65896 42464
rect 65960 42400 65968 42464
rect 65648 42399 65968 42400
rect 96368 42464 96688 42465
rect 96368 42400 96376 42464
rect 96440 42400 96456 42464
rect 96520 42400 96536 42464
rect 96600 42400 96616 42464
rect 96680 42400 96688 42464
rect 96368 42399 96688 42400
rect 127088 42464 127408 42465
rect 127088 42400 127096 42464
rect 127160 42400 127176 42464
rect 127240 42400 127256 42464
rect 127320 42400 127336 42464
rect 127400 42400 127408 42464
rect 127088 42399 127408 42400
rect 157808 42464 158128 42465
rect 157808 42400 157816 42464
rect 157880 42400 157896 42464
rect 157960 42400 157976 42464
rect 158040 42400 158056 42464
rect 158120 42400 158128 42464
rect 157808 42399 158128 42400
rect 19568 41920 19888 41921
rect 19568 41856 19576 41920
rect 19640 41856 19656 41920
rect 19720 41856 19736 41920
rect 19800 41856 19816 41920
rect 19880 41856 19888 41920
rect 19568 41855 19888 41856
rect 50288 41920 50608 41921
rect 50288 41856 50296 41920
rect 50360 41856 50376 41920
rect 50440 41856 50456 41920
rect 50520 41856 50536 41920
rect 50600 41856 50608 41920
rect 50288 41855 50608 41856
rect 81008 41920 81328 41921
rect 81008 41856 81016 41920
rect 81080 41856 81096 41920
rect 81160 41856 81176 41920
rect 81240 41856 81256 41920
rect 81320 41856 81328 41920
rect 81008 41855 81328 41856
rect 111728 41920 112048 41921
rect 111728 41856 111736 41920
rect 111800 41856 111816 41920
rect 111880 41856 111896 41920
rect 111960 41856 111976 41920
rect 112040 41856 112048 41920
rect 111728 41855 112048 41856
rect 142448 41920 142768 41921
rect 142448 41856 142456 41920
rect 142520 41856 142536 41920
rect 142600 41856 142616 41920
rect 142680 41856 142696 41920
rect 142760 41856 142768 41920
rect 142448 41855 142768 41856
rect 173168 41920 173488 41921
rect 173168 41856 173176 41920
rect 173240 41856 173256 41920
rect 173320 41856 173336 41920
rect 173400 41856 173416 41920
rect 173480 41856 173488 41920
rect 173168 41855 173488 41856
rect 4208 41376 4528 41377
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 41311 4528 41312
rect 34928 41376 35248 41377
rect 34928 41312 34936 41376
rect 35000 41312 35016 41376
rect 35080 41312 35096 41376
rect 35160 41312 35176 41376
rect 35240 41312 35248 41376
rect 34928 41311 35248 41312
rect 65648 41376 65968 41377
rect 65648 41312 65656 41376
rect 65720 41312 65736 41376
rect 65800 41312 65816 41376
rect 65880 41312 65896 41376
rect 65960 41312 65968 41376
rect 65648 41311 65968 41312
rect 96368 41376 96688 41377
rect 96368 41312 96376 41376
rect 96440 41312 96456 41376
rect 96520 41312 96536 41376
rect 96600 41312 96616 41376
rect 96680 41312 96688 41376
rect 96368 41311 96688 41312
rect 127088 41376 127408 41377
rect 127088 41312 127096 41376
rect 127160 41312 127176 41376
rect 127240 41312 127256 41376
rect 127320 41312 127336 41376
rect 127400 41312 127408 41376
rect 127088 41311 127408 41312
rect 157808 41376 158128 41377
rect 157808 41312 157816 41376
rect 157880 41312 157896 41376
rect 157960 41312 157976 41376
rect 158040 41312 158056 41376
rect 158120 41312 158128 41376
rect 157808 41311 158128 41312
rect 19568 40832 19888 40833
rect 19568 40768 19576 40832
rect 19640 40768 19656 40832
rect 19720 40768 19736 40832
rect 19800 40768 19816 40832
rect 19880 40768 19888 40832
rect 19568 40767 19888 40768
rect 50288 40832 50608 40833
rect 50288 40768 50296 40832
rect 50360 40768 50376 40832
rect 50440 40768 50456 40832
rect 50520 40768 50536 40832
rect 50600 40768 50608 40832
rect 50288 40767 50608 40768
rect 81008 40832 81328 40833
rect 81008 40768 81016 40832
rect 81080 40768 81096 40832
rect 81160 40768 81176 40832
rect 81240 40768 81256 40832
rect 81320 40768 81328 40832
rect 81008 40767 81328 40768
rect 111728 40832 112048 40833
rect 111728 40768 111736 40832
rect 111800 40768 111816 40832
rect 111880 40768 111896 40832
rect 111960 40768 111976 40832
rect 112040 40768 112048 40832
rect 111728 40767 112048 40768
rect 142448 40832 142768 40833
rect 142448 40768 142456 40832
rect 142520 40768 142536 40832
rect 142600 40768 142616 40832
rect 142680 40768 142696 40832
rect 142760 40768 142768 40832
rect 142448 40767 142768 40768
rect 173168 40832 173488 40833
rect 173168 40768 173176 40832
rect 173240 40768 173256 40832
rect 173320 40768 173336 40832
rect 173400 40768 173416 40832
rect 173480 40768 173488 40832
rect 173168 40767 173488 40768
rect 4208 40288 4528 40289
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 40223 4528 40224
rect 34928 40288 35248 40289
rect 34928 40224 34936 40288
rect 35000 40224 35016 40288
rect 35080 40224 35096 40288
rect 35160 40224 35176 40288
rect 35240 40224 35248 40288
rect 34928 40223 35248 40224
rect 65648 40288 65968 40289
rect 65648 40224 65656 40288
rect 65720 40224 65736 40288
rect 65800 40224 65816 40288
rect 65880 40224 65896 40288
rect 65960 40224 65968 40288
rect 65648 40223 65968 40224
rect 96368 40288 96688 40289
rect 96368 40224 96376 40288
rect 96440 40224 96456 40288
rect 96520 40224 96536 40288
rect 96600 40224 96616 40288
rect 96680 40224 96688 40288
rect 96368 40223 96688 40224
rect 127088 40288 127408 40289
rect 127088 40224 127096 40288
rect 127160 40224 127176 40288
rect 127240 40224 127256 40288
rect 127320 40224 127336 40288
rect 127400 40224 127408 40288
rect 127088 40223 127408 40224
rect 157808 40288 158128 40289
rect 157808 40224 157816 40288
rect 157880 40224 157896 40288
rect 157960 40224 157976 40288
rect 158040 40224 158056 40288
rect 158120 40224 158128 40288
rect 157808 40223 158128 40224
rect 19568 39744 19888 39745
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 19568 39679 19888 39680
rect 50288 39744 50608 39745
rect 50288 39680 50296 39744
rect 50360 39680 50376 39744
rect 50440 39680 50456 39744
rect 50520 39680 50536 39744
rect 50600 39680 50608 39744
rect 50288 39679 50608 39680
rect 81008 39744 81328 39745
rect 81008 39680 81016 39744
rect 81080 39680 81096 39744
rect 81160 39680 81176 39744
rect 81240 39680 81256 39744
rect 81320 39680 81328 39744
rect 81008 39679 81328 39680
rect 111728 39744 112048 39745
rect 111728 39680 111736 39744
rect 111800 39680 111816 39744
rect 111880 39680 111896 39744
rect 111960 39680 111976 39744
rect 112040 39680 112048 39744
rect 111728 39679 112048 39680
rect 142448 39744 142768 39745
rect 142448 39680 142456 39744
rect 142520 39680 142536 39744
rect 142600 39680 142616 39744
rect 142680 39680 142696 39744
rect 142760 39680 142768 39744
rect 142448 39679 142768 39680
rect 173168 39744 173488 39745
rect 173168 39680 173176 39744
rect 173240 39680 173256 39744
rect 173320 39680 173336 39744
rect 173400 39680 173416 39744
rect 173480 39680 173488 39744
rect 173168 39679 173488 39680
rect 4208 39200 4528 39201
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 39135 4528 39136
rect 34928 39200 35248 39201
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 39135 35248 39136
rect 65648 39200 65968 39201
rect 65648 39136 65656 39200
rect 65720 39136 65736 39200
rect 65800 39136 65816 39200
rect 65880 39136 65896 39200
rect 65960 39136 65968 39200
rect 65648 39135 65968 39136
rect 96368 39200 96688 39201
rect 96368 39136 96376 39200
rect 96440 39136 96456 39200
rect 96520 39136 96536 39200
rect 96600 39136 96616 39200
rect 96680 39136 96688 39200
rect 96368 39135 96688 39136
rect 127088 39200 127408 39201
rect 127088 39136 127096 39200
rect 127160 39136 127176 39200
rect 127240 39136 127256 39200
rect 127320 39136 127336 39200
rect 127400 39136 127408 39200
rect 127088 39135 127408 39136
rect 157808 39200 158128 39201
rect 157808 39136 157816 39200
rect 157880 39136 157896 39200
rect 157960 39136 157976 39200
rect 158040 39136 158056 39200
rect 158120 39136 158128 39200
rect 157808 39135 158128 39136
rect 19568 38656 19888 38657
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 38591 19888 38592
rect 50288 38656 50608 38657
rect 50288 38592 50296 38656
rect 50360 38592 50376 38656
rect 50440 38592 50456 38656
rect 50520 38592 50536 38656
rect 50600 38592 50608 38656
rect 50288 38591 50608 38592
rect 81008 38656 81328 38657
rect 81008 38592 81016 38656
rect 81080 38592 81096 38656
rect 81160 38592 81176 38656
rect 81240 38592 81256 38656
rect 81320 38592 81328 38656
rect 81008 38591 81328 38592
rect 111728 38656 112048 38657
rect 111728 38592 111736 38656
rect 111800 38592 111816 38656
rect 111880 38592 111896 38656
rect 111960 38592 111976 38656
rect 112040 38592 112048 38656
rect 111728 38591 112048 38592
rect 142448 38656 142768 38657
rect 142448 38592 142456 38656
rect 142520 38592 142536 38656
rect 142600 38592 142616 38656
rect 142680 38592 142696 38656
rect 142760 38592 142768 38656
rect 142448 38591 142768 38592
rect 173168 38656 173488 38657
rect 173168 38592 173176 38656
rect 173240 38592 173256 38656
rect 173320 38592 173336 38656
rect 173400 38592 173416 38656
rect 173480 38592 173488 38656
rect 173168 38591 173488 38592
rect 4208 38112 4528 38113
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 38047 4528 38048
rect 34928 38112 35248 38113
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 38047 35248 38048
rect 65648 38112 65968 38113
rect 65648 38048 65656 38112
rect 65720 38048 65736 38112
rect 65800 38048 65816 38112
rect 65880 38048 65896 38112
rect 65960 38048 65968 38112
rect 65648 38047 65968 38048
rect 96368 38112 96688 38113
rect 96368 38048 96376 38112
rect 96440 38048 96456 38112
rect 96520 38048 96536 38112
rect 96600 38048 96616 38112
rect 96680 38048 96688 38112
rect 96368 38047 96688 38048
rect 127088 38112 127408 38113
rect 127088 38048 127096 38112
rect 127160 38048 127176 38112
rect 127240 38048 127256 38112
rect 127320 38048 127336 38112
rect 127400 38048 127408 38112
rect 127088 38047 127408 38048
rect 157808 38112 158128 38113
rect 157808 38048 157816 38112
rect 157880 38048 157896 38112
rect 157960 38048 157976 38112
rect 158040 38048 158056 38112
rect 158120 38048 158128 38112
rect 157808 38047 158128 38048
rect 19568 37568 19888 37569
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 37503 19888 37504
rect 50288 37568 50608 37569
rect 50288 37504 50296 37568
rect 50360 37504 50376 37568
rect 50440 37504 50456 37568
rect 50520 37504 50536 37568
rect 50600 37504 50608 37568
rect 50288 37503 50608 37504
rect 81008 37568 81328 37569
rect 81008 37504 81016 37568
rect 81080 37504 81096 37568
rect 81160 37504 81176 37568
rect 81240 37504 81256 37568
rect 81320 37504 81328 37568
rect 81008 37503 81328 37504
rect 111728 37568 112048 37569
rect 111728 37504 111736 37568
rect 111800 37504 111816 37568
rect 111880 37504 111896 37568
rect 111960 37504 111976 37568
rect 112040 37504 112048 37568
rect 111728 37503 112048 37504
rect 142448 37568 142768 37569
rect 142448 37504 142456 37568
rect 142520 37504 142536 37568
rect 142600 37504 142616 37568
rect 142680 37504 142696 37568
rect 142760 37504 142768 37568
rect 142448 37503 142768 37504
rect 173168 37568 173488 37569
rect 173168 37504 173176 37568
rect 173240 37504 173256 37568
rect 173320 37504 173336 37568
rect 173400 37504 173416 37568
rect 173480 37504 173488 37568
rect 173168 37503 173488 37504
rect 4208 37024 4528 37025
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 34928 37024 35248 37025
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 36959 35248 36960
rect 65648 37024 65968 37025
rect 65648 36960 65656 37024
rect 65720 36960 65736 37024
rect 65800 36960 65816 37024
rect 65880 36960 65896 37024
rect 65960 36960 65968 37024
rect 65648 36959 65968 36960
rect 96368 37024 96688 37025
rect 96368 36960 96376 37024
rect 96440 36960 96456 37024
rect 96520 36960 96536 37024
rect 96600 36960 96616 37024
rect 96680 36960 96688 37024
rect 96368 36959 96688 36960
rect 127088 37024 127408 37025
rect 127088 36960 127096 37024
rect 127160 36960 127176 37024
rect 127240 36960 127256 37024
rect 127320 36960 127336 37024
rect 127400 36960 127408 37024
rect 127088 36959 127408 36960
rect 157808 37024 158128 37025
rect 157808 36960 157816 37024
rect 157880 36960 157896 37024
rect 157960 36960 157976 37024
rect 158040 36960 158056 37024
rect 158120 36960 158128 37024
rect 157808 36959 158128 36960
rect 19568 36480 19888 36481
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 36415 19888 36416
rect 50288 36480 50608 36481
rect 50288 36416 50296 36480
rect 50360 36416 50376 36480
rect 50440 36416 50456 36480
rect 50520 36416 50536 36480
rect 50600 36416 50608 36480
rect 50288 36415 50608 36416
rect 81008 36480 81328 36481
rect 81008 36416 81016 36480
rect 81080 36416 81096 36480
rect 81160 36416 81176 36480
rect 81240 36416 81256 36480
rect 81320 36416 81328 36480
rect 81008 36415 81328 36416
rect 111728 36480 112048 36481
rect 111728 36416 111736 36480
rect 111800 36416 111816 36480
rect 111880 36416 111896 36480
rect 111960 36416 111976 36480
rect 112040 36416 112048 36480
rect 111728 36415 112048 36416
rect 142448 36480 142768 36481
rect 142448 36416 142456 36480
rect 142520 36416 142536 36480
rect 142600 36416 142616 36480
rect 142680 36416 142696 36480
rect 142760 36416 142768 36480
rect 142448 36415 142768 36416
rect 173168 36480 173488 36481
rect 173168 36416 173176 36480
rect 173240 36416 173256 36480
rect 173320 36416 173336 36480
rect 173400 36416 173416 36480
rect 173480 36416 173488 36480
rect 173168 36415 173488 36416
rect 4208 35936 4528 35937
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 34928 35936 35248 35937
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 35871 35248 35872
rect 65648 35936 65968 35937
rect 65648 35872 65656 35936
rect 65720 35872 65736 35936
rect 65800 35872 65816 35936
rect 65880 35872 65896 35936
rect 65960 35872 65968 35936
rect 65648 35871 65968 35872
rect 96368 35936 96688 35937
rect 96368 35872 96376 35936
rect 96440 35872 96456 35936
rect 96520 35872 96536 35936
rect 96600 35872 96616 35936
rect 96680 35872 96688 35936
rect 96368 35871 96688 35872
rect 127088 35936 127408 35937
rect 127088 35872 127096 35936
rect 127160 35872 127176 35936
rect 127240 35872 127256 35936
rect 127320 35872 127336 35936
rect 127400 35872 127408 35936
rect 127088 35871 127408 35872
rect 157808 35936 158128 35937
rect 157808 35872 157816 35936
rect 157880 35872 157896 35936
rect 157960 35872 157976 35936
rect 158040 35872 158056 35936
rect 158120 35872 158128 35936
rect 157808 35871 158128 35872
rect 19568 35392 19888 35393
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 35327 19888 35328
rect 50288 35392 50608 35393
rect 50288 35328 50296 35392
rect 50360 35328 50376 35392
rect 50440 35328 50456 35392
rect 50520 35328 50536 35392
rect 50600 35328 50608 35392
rect 50288 35327 50608 35328
rect 81008 35392 81328 35393
rect 81008 35328 81016 35392
rect 81080 35328 81096 35392
rect 81160 35328 81176 35392
rect 81240 35328 81256 35392
rect 81320 35328 81328 35392
rect 81008 35327 81328 35328
rect 111728 35392 112048 35393
rect 111728 35328 111736 35392
rect 111800 35328 111816 35392
rect 111880 35328 111896 35392
rect 111960 35328 111976 35392
rect 112040 35328 112048 35392
rect 111728 35327 112048 35328
rect 142448 35392 142768 35393
rect 142448 35328 142456 35392
rect 142520 35328 142536 35392
rect 142600 35328 142616 35392
rect 142680 35328 142696 35392
rect 142760 35328 142768 35392
rect 142448 35327 142768 35328
rect 173168 35392 173488 35393
rect 173168 35328 173176 35392
rect 173240 35328 173256 35392
rect 173320 35328 173336 35392
rect 173400 35328 173416 35392
rect 173480 35328 173488 35392
rect 173168 35327 173488 35328
rect 4208 34848 4528 34849
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 34928 34848 35248 34849
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 34783 35248 34784
rect 65648 34848 65968 34849
rect 65648 34784 65656 34848
rect 65720 34784 65736 34848
rect 65800 34784 65816 34848
rect 65880 34784 65896 34848
rect 65960 34784 65968 34848
rect 65648 34783 65968 34784
rect 96368 34848 96688 34849
rect 96368 34784 96376 34848
rect 96440 34784 96456 34848
rect 96520 34784 96536 34848
rect 96600 34784 96616 34848
rect 96680 34784 96688 34848
rect 96368 34783 96688 34784
rect 127088 34848 127408 34849
rect 127088 34784 127096 34848
rect 127160 34784 127176 34848
rect 127240 34784 127256 34848
rect 127320 34784 127336 34848
rect 127400 34784 127408 34848
rect 127088 34783 127408 34784
rect 157808 34848 158128 34849
rect 157808 34784 157816 34848
rect 157880 34784 157896 34848
rect 157960 34784 157976 34848
rect 158040 34784 158056 34848
rect 158120 34784 158128 34848
rect 157808 34783 158128 34784
rect 19568 34304 19888 34305
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 34239 19888 34240
rect 50288 34304 50608 34305
rect 50288 34240 50296 34304
rect 50360 34240 50376 34304
rect 50440 34240 50456 34304
rect 50520 34240 50536 34304
rect 50600 34240 50608 34304
rect 50288 34239 50608 34240
rect 81008 34304 81328 34305
rect 81008 34240 81016 34304
rect 81080 34240 81096 34304
rect 81160 34240 81176 34304
rect 81240 34240 81256 34304
rect 81320 34240 81328 34304
rect 81008 34239 81328 34240
rect 111728 34304 112048 34305
rect 111728 34240 111736 34304
rect 111800 34240 111816 34304
rect 111880 34240 111896 34304
rect 111960 34240 111976 34304
rect 112040 34240 112048 34304
rect 111728 34239 112048 34240
rect 142448 34304 142768 34305
rect 142448 34240 142456 34304
rect 142520 34240 142536 34304
rect 142600 34240 142616 34304
rect 142680 34240 142696 34304
rect 142760 34240 142768 34304
rect 142448 34239 142768 34240
rect 173168 34304 173488 34305
rect 173168 34240 173176 34304
rect 173240 34240 173256 34304
rect 173320 34240 173336 34304
rect 173400 34240 173416 34304
rect 173480 34240 173488 34304
rect 173168 34239 173488 34240
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 34928 33760 35248 33761
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 33695 35248 33696
rect 65648 33760 65968 33761
rect 65648 33696 65656 33760
rect 65720 33696 65736 33760
rect 65800 33696 65816 33760
rect 65880 33696 65896 33760
rect 65960 33696 65968 33760
rect 65648 33695 65968 33696
rect 96368 33760 96688 33761
rect 96368 33696 96376 33760
rect 96440 33696 96456 33760
rect 96520 33696 96536 33760
rect 96600 33696 96616 33760
rect 96680 33696 96688 33760
rect 96368 33695 96688 33696
rect 127088 33760 127408 33761
rect 127088 33696 127096 33760
rect 127160 33696 127176 33760
rect 127240 33696 127256 33760
rect 127320 33696 127336 33760
rect 127400 33696 127408 33760
rect 127088 33695 127408 33696
rect 157808 33760 158128 33761
rect 157808 33696 157816 33760
rect 157880 33696 157896 33760
rect 157960 33696 157976 33760
rect 158040 33696 158056 33760
rect 158120 33696 158128 33760
rect 157808 33695 158128 33696
rect 19568 33216 19888 33217
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 33151 19888 33152
rect 50288 33216 50608 33217
rect 50288 33152 50296 33216
rect 50360 33152 50376 33216
rect 50440 33152 50456 33216
rect 50520 33152 50536 33216
rect 50600 33152 50608 33216
rect 50288 33151 50608 33152
rect 81008 33216 81328 33217
rect 81008 33152 81016 33216
rect 81080 33152 81096 33216
rect 81160 33152 81176 33216
rect 81240 33152 81256 33216
rect 81320 33152 81328 33216
rect 81008 33151 81328 33152
rect 111728 33216 112048 33217
rect 111728 33152 111736 33216
rect 111800 33152 111816 33216
rect 111880 33152 111896 33216
rect 111960 33152 111976 33216
rect 112040 33152 112048 33216
rect 111728 33151 112048 33152
rect 142448 33216 142768 33217
rect 142448 33152 142456 33216
rect 142520 33152 142536 33216
rect 142600 33152 142616 33216
rect 142680 33152 142696 33216
rect 142760 33152 142768 33216
rect 142448 33151 142768 33152
rect 173168 33216 173488 33217
rect 173168 33152 173176 33216
rect 173240 33152 173256 33216
rect 173320 33152 173336 33216
rect 173400 33152 173416 33216
rect 173480 33152 173488 33216
rect 173168 33151 173488 33152
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 34928 32672 35248 32673
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 32607 35248 32608
rect 65648 32672 65968 32673
rect 65648 32608 65656 32672
rect 65720 32608 65736 32672
rect 65800 32608 65816 32672
rect 65880 32608 65896 32672
rect 65960 32608 65968 32672
rect 65648 32607 65968 32608
rect 96368 32672 96688 32673
rect 96368 32608 96376 32672
rect 96440 32608 96456 32672
rect 96520 32608 96536 32672
rect 96600 32608 96616 32672
rect 96680 32608 96688 32672
rect 96368 32607 96688 32608
rect 127088 32672 127408 32673
rect 127088 32608 127096 32672
rect 127160 32608 127176 32672
rect 127240 32608 127256 32672
rect 127320 32608 127336 32672
rect 127400 32608 127408 32672
rect 127088 32607 127408 32608
rect 157808 32672 158128 32673
rect 157808 32608 157816 32672
rect 157880 32608 157896 32672
rect 157960 32608 157976 32672
rect 158040 32608 158056 32672
rect 158120 32608 158128 32672
rect 157808 32607 158128 32608
rect 19568 32128 19888 32129
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 32063 19888 32064
rect 50288 32128 50608 32129
rect 50288 32064 50296 32128
rect 50360 32064 50376 32128
rect 50440 32064 50456 32128
rect 50520 32064 50536 32128
rect 50600 32064 50608 32128
rect 50288 32063 50608 32064
rect 81008 32128 81328 32129
rect 81008 32064 81016 32128
rect 81080 32064 81096 32128
rect 81160 32064 81176 32128
rect 81240 32064 81256 32128
rect 81320 32064 81328 32128
rect 81008 32063 81328 32064
rect 111728 32128 112048 32129
rect 111728 32064 111736 32128
rect 111800 32064 111816 32128
rect 111880 32064 111896 32128
rect 111960 32064 111976 32128
rect 112040 32064 112048 32128
rect 111728 32063 112048 32064
rect 142448 32128 142768 32129
rect 142448 32064 142456 32128
rect 142520 32064 142536 32128
rect 142600 32064 142616 32128
rect 142680 32064 142696 32128
rect 142760 32064 142768 32128
rect 142448 32063 142768 32064
rect 173168 32128 173488 32129
rect 173168 32064 173176 32128
rect 173240 32064 173256 32128
rect 173320 32064 173336 32128
rect 173400 32064 173416 32128
rect 173480 32064 173488 32128
rect 173168 32063 173488 32064
rect 4208 31584 4528 31585
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 34928 31584 35248 31585
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 31519 35248 31520
rect 65648 31584 65968 31585
rect 65648 31520 65656 31584
rect 65720 31520 65736 31584
rect 65800 31520 65816 31584
rect 65880 31520 65896 31584
rect 65960 31520 65968 31584
rect 65648 31519 65968 31520
rect 96368 31584 96688 31585
rect 96368 31520 96376 31584
rect 96440 31520 96456 31584
rect 96520 31520 96536 31584
rect 96600 31520 96616 31584
rect 96680 31520 96688 31584
rect 96368 31519 96688 31520
rect 127088 31584 127408 31585
rect 127088 31520 127096 31584
rect 127160 31520 127176 31584
rect 127240 31520 127256 31584
rect 127320 31520 127336 31584
rect 127400 31520 127408 31584
rect 127088 31519 127408 31520
rect 157808 31584 158128 31585
rect 157808 31520 157816 31584
rect 157880 31520 157896 31584
rect 157960 31520 157976 31584
rect 158040 31520 158056 31584
rect 158120 31520 158128 31584
rect 157808 31519 158128 31520
rect 19568 31040 19888 31041
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 30975 19888 30976
rect 50288 31040 50608 31041
rect 50288 30976 50296 31040
rect 50360 30976 50376 31040
rect 50440 30976 50456 31040
rect 50520 30976 50536 31040
rect 50600 30976 50608 31040
rect 50288 30975 50608 30976
rect 81008 31040 81328 31041
rect 81008 30976 81016 31040
rect 81080 30976 81096 31040
rect 81160 30976 81176 31040
rect 81240 30976 81256 31040
rect 81320 30976 81328 31040
rect 81008 30975 81328 30976
rect 111728 31040 112048 31041
rect 111728 30976 111736 31040
rect 111800 30976 111816 31040
rect 111880 30976 111896 31040
rect 111960 30976 111976 31040
rect 112040 30976 112048 31040
rect 111728 30975 112048 30976
rect 142448 31040 142768 31041
rect 142448 30976 142456 31040
rect 142520 30976 142536 31040
rect 142600 30976 142616 31040
rect 142680 30976 142696 31040
rect 142760 30976 142768 31040
rect 142448 30975 142768 30976
rect 173168 31040 173488 31041
rect 173168 30976 173176 31040
rect 173240 30976 173256 31040
rect 173320 30976 173336 31040
rect 173400 30976 173416 31040
rect 173480 30976 173488 31040
rect 173168 30975 173488 30976
rect 4208 30496 4528 30497
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 34928 30496 35248 30497
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 30431 35248 30432
rect 65648 30496 65968 30497
rect 65648 30432 65656 30496
rect 65720 30432 65736 30496
rect 65800 30432 65816 30496
rect 65880 30432 65896 30496
rect 65960 30432 65968 30496
rect 65648 30431 65968 30432
rect 96368 30496 96688 30497
rect 96368 30432 96376 30496
rect 96440 30432 96456 30496
rect 96520 30432 96536 30496
rect 96600 30432 96616 30496
rect 96680 30432 96688 30496
rect 96368 30431 96688 30432
rect 127088 30496 127408 30497
rect 127088 30432 127096 30496
rect 127160 30432 127176 30496
rect 127240 30432 127256 30496
rect 127320 30432 127336 30496
rect 127400 30432 127408 30496
rect 127088 30431 127408 30432
rect 157808 30496 158128 30497
rect 157808 30432 157816 30496
rect 157880 30432 157896 30496
rect 157960 30432 157976 30496
rect 158040 30432 158056 30496
rect 158120 30432 158128 30496
rect 157808 30431 158128 30432
rect 19568 29952 19888 29953
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 29887 19888 29888
rect 50288 29952 50608 29953
rect 50288 29888 50296 29952
rect 50360 29888 50376 29952
rect 50440 29888 50456 29952
rect 50520 29888 50536 29952
rect 50600 29888 50608 29952
rect 50288 29887 50608 29888
rect 81008 29952 81328 29953
rect 81008 29888 81016 29952
rect 81080 29888 81096 29952
rect 81160 29888 81176 29952
rect 81240 29888 81256 29952
rect 81320 29888 81328 29952
rect 81008 29887 81328 29888
rect 111728 29952 112048 29953
rect 111728 29888 111736 29952
rect 111800 29888 111816 29952
rect 111880 29888 111896 29952
rect 111960 29888 111976 29952
rect 112040 29888 112048 29952
rect 111728 29887 112048 29888
rect 142448 29952 142768 29953
rect 142448 29888 142456 29952
rect 142520 29888 142536 29952
rect 142600 29888 142616 29952
rect 142680 29888 142696 29952
rect 142760 29888 142768 29952
rect 142448 29887 142768 29888
rect 173168 29952 173488 29953
rect 173168 29888 173176 29952
rect 173240 29888 173256 29952
rect 173320 29888 173336 29952
rect 173400 29888 173416 29952
rect 173480 29888 173488 29952
rect 173168 29887 173488 29888
rect 4208 29408 4528 29409
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 34928 29408 35248 29409
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 29343 35248 29344
rect 65648 29408 65968 29409
rect 65648 29344 65656 29408
rect 65720 29344 65736 29408
rect 65800 29344 65816 29408
rect 65880 29344 65896 29408
rect 65960 29344 65968 29408
rect 65648 29343 65968 29344
rect 96368 29408 96688 29409
rect 96368 29344 96376 29408
rect 96440 29344 96456 29408
rect 96520 29344 96536 29408
rect 96600 29344 96616 29408
rect 96680 29344 96688 29408
rect 96368 29343 96688 29344
rect 127088 29408 127408 29409
rect 127088 29344 127096 29408
rect 127160 29344 127176 29408
rect 127240 29344 127256 29408
rect 127320 29344 127336 29408
rect 127400 29344 127408 29408
rect 127088 29343 127408 29344
rect 157808 29408 158128 29409
rect 157808 29344 157816 29408
rect 157880 29344 157896 29408
rect 157960 29344 157976 29408
rect 158040 29344 158056 29408
rect 158120 29344 158128 29408
rect 157808 29343 158128 29344
rect 19568 28864 19888 28865
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 28799 19888 28800
rect 50288 28864 50608 28865
rect 50288 28800 50296 28864
rect 50360 28800 50376 28864
rect 50440 28800 50456 28864
rect 50520 28800 50536 28864
rect 50600 28800 50608 28864
rect 50288 28799 50608 28800
rect 81008 28864 81328 28865
rect 81008 28800 81016 28864
rect 81080 28800 81096 28864
rect 81160 28800 81176 28864
rect 81240 28800 81256 28864
rect 81320 28800 81328 28864
rect 81008 28799 81328 28800
rect 111728 28864 112048 28865
rect 111728 28800 111736 28864
rect 111800 28800 111816 28864
rect 111880 28800 111896 28864
rect 111960 28800 111976 28864
rect 112040 28800 112048 28864
rect 111728 28799 112048 28800
rect 142448 28864 142768 28865
rect 142448 28800 142456 28864
rect 142520 28800 142536 28864
rect 142600 28800 142616 28864
rect 142680 28800 142696 28864
rect 142760 28800 142768 28864
rect 142448 28799 142768 28800
rect 173168 28864 173488 28865
rect 173168 28800 173176 28864
rect 173240 28800 173256 28864
rect 173320 28800 173336 28864
rect 173400 28800 173416 28864
rect 173480 28800 173488 28864
rect 173168 28799 173488 28800
rect 4208 28320 4528 28321
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 34928 28320 35248 28321
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 28255 35248 28256
rect 65648 28320 65968 28321
rect 65648 28256 65656 28320
rect 65720 28256 65736 28320
rect 65800 28256 65816 28320
rect 65880 28256 65896 28320
rect 65960 28256 65968 28320
rect 65648 28255 65968 28256
rect 96368 28320 96688 28321
rect 96368 28256 96376 28320
rect 96440 28256 96456 28320
rect 96520 28256 96536 28320
rect 96600 28256 96616 28320
rect 96680 28256 96688 28320
rect 96368 28255 96688 28256
rect 127088 28320 127408 28321
rect 127088 28256 127096 28320
rect 127160 28256 127176 28320
rect 127240 28256 127256 28320
rect 127320 28256 127336 28320
rect 127400 28256 127408 28320
rect 127088 28255 127408 28256
rect 157808 28320 158128 28321
rect 157808 28256 157816 28320
rect 157880 28256 157896 28320
rect 157960 28256 157976 28320
rect 158040 28256 158056 28320
rect 158120 28256 158128 28320
rect 157808 28255 158128 28256
rect 19568 27776 19888 27777
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 27711 19888 27712
rect 50288 27776 50608 27777
rect 50288 27712 50296 27776
rect 50360 27712 50376 27776
rect 50440 27712 50456 27776
rect 50520 27712 50536 27776
rect 50600 27712 50608 27776
rect 50288 27711 50608 27712
rect 81008 27776 81328 27777
rect 81008 27712 81016 27776
rect 81080 27712 81096 27776
rect 81160 27712 81176 27776
rect 81240 27712 81256 27776
rect 81320 27712 81328 27776
rect 81008 27711 81328 27712
rect 111728 27776 112048 27777
rect 111728 27712 111736 27776
rect 111800 27712 111816 27776
rect 111880 27712 111896 27776
rect 111960 27712 111976 27776
rect 112040 27712 112048 27776
rect 111728 27711 112048 27712
rect 142448 27776 142768 27777
rect 142448 27712 142456 27776
rect 142520 27712 142536 27776
rect 142600 27712 142616 27776
rect 142680 27712 142696 27776
rect 142760 27712 142768 27776
rect 142448 27711 142768 27712
rect 173168 27776 173488 27777
rect 173168 27712 173176 27776
rect 173240 27712 173256 27776
rect 173320 27712 173336 27776
rect 173400 27712 173416 27776
rect 173480 27712 173488 27776
rect 173168 27711 173488 27712
rect 4208 27232 4528 27233
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 34928 27232 35248 27233
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 27167 35248 27168
rect 65648 27232 65968 27233
rect 65648 27168 65656 27232
rect 65720 27168 65736 27232
rect 65800 27168 65816 27232
rect 65880 27168 65896 27232
rect 65960 27168 65968 27232
rect 65648 27167 65968 27168
rect 96368 27232 96688 27233
rect 96368 27168 96376 27232
rect 96440 27168 96456 27232
rect 96520 27168 96536 27232
rect 96600 27168 96616 27232
rect 96680 27168 96688 27232
rect 96368 27167 96688 27168
rect 127088 27232 127408 27233
rect 127088 27168 127096 27232
rect 127160 27168 127176 27232
rect 127240 27168 127256 27232
rect 127320 27168 127336 27232
rect 127400 27168 127408 27232
rect 127088 27167 127408 27168
rect 157808 27232 158128 27233
rect 157808 27168 157816 27232
rect 157880 27168 157896 27232
rect 157960 27168 157976 27232
rect 158040 27168 158056 27232
rect 158120 27168 158128 27232
rect 157808 27167 158128 27168
rect 19568 26688 19888 26689
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 26623 19888 26624
rect 50288 26688 50608 26689
rect 50288 26624 50296 26688
rect 50360 26624 50376 26688
rect 50440 26624 50456 26688
rect 50520 26624 50536 26688
rect 50600 26624 50608 26688
rect 50288 26623 50608 26624
rect 81008 26688 81328 26689
rect 81008 26624 81016 26688
rect 81080 26624 81096 26688
rect 81160 26624 81176 26688
rect 81240 26624 81256 26688
rect 81320 26624 81328 26688
rect 81008 26623 81328 26624
rect 111728 26688 112048 26689
rect 111728 26624 111736 26688
rect 111800 26624 111816 26688
rect 111880 26624 111896 26688
rect 111960 26624 111976 26688
rect 112040 26624 112048 26688
rect 111728 26623 112048 26624
rect 142448 26688 142768 26689
rect 142448 26624 142456 26688
rect 142520 26624 142536 26688
rect 142600 26624 142616 26688
rect 142680 26624 142696 26688
rect 142760 26624 142768 26688
rect 142448 26623 142768 26624
rect 173168 26688 173488 26689
rect 173168 26624 173176 26688
rect 173240 26624 173256 26688
rect 173320 26624 173336 26688
rect 173400 26624 173416 26688
rect 173480 26624 173488 26688
rect 173168 26623 173488 26624
rect 4208 26144 4528 26145
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 34928 26144 35248 26145
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 26079 35248 26080
rect 65648 26144 65968 26145
rect 65648 26080 65656 26144
rect 65720 26080 65736 26144
rect 65800 26080 65816 26144
rect 65880 26080 65896 26144
rect 65960 26080 65968 26144
rect 65648 26079 65968 26080
rect 96368 26144 96688 26145
rect 96368 26080 96376 26144
rect 96440 26080 96456 26144
rect 96520 26080 96536 26144
rect 96600 26080 96616 26144
rect 96680 26080 96688 26144
rect 96368 26079 96688 26080
rect 127088 26144 127408 26145
rect 127088 26080 127096 26144
rect 127160 26080 127176 26144
rect 127240 26080 127256 26144
rect 127320 26080 127336 26144
rect 127400 26080 127408 26144
rect 127088 26079 127408 26080
rect 157808 26144 158128 26145
rect 157808 26080 157816 26144
rect 157880 26080 157896 26144
rect 157960 26080 157976 26144
rect 158040 26080 158056 26144
rect 158120 26080 158128 26144
rect 157808 26079 158128 26080
rect 19568 25600 19888 25601
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 25535 19888 25536
rect 50288 25600 50608 25601
rect 50288 25536 50296 25600
rect 50360 25536 50376 25600
rect 50440 25536 50456 25600
rect 50520 25536 50536 25600
rect 50600 25536 50608 25600
rect 50288 25535 50608 25536
rect 81008 25600 81328 25601
rect 81008 25536 81016 25600
rect 81080 25536 81096 25600
rect 81160 25536 81176 25600
rect 81240 25536 81256 25600
rect 81320 25536 81328 25600
rect 81008 25535 81328 25536
rect 111728 25600 112048 25601
rect 111728 25536 111736 25600
rect 111800 25536 111816 25600
rect 111880 25536 111896 25600
rect 111960 25536 111976 25600
rect 112040 25536 112048 25600
rect 111728 25535 112048 25536
rect 142448 25600 142768 25601
rect 142448 25536 142456 25600
rect 142520 25536 142536 25600
rect 142600 25536 142616 25600
rect 142680 25536 142696 25600
rect 142760 25536 142768 25600
rect 142448 25535 142768 25536
rect 173168 25600 173488 25601
rect 173168 25536 173176 25600
rect 173240 25536 173256 25600
rect 173320 25536 173336 25600
rect 173400 25536 173416 25600
rect 173480 25536 173488 25600
rect 173168 25535 173488 25536
rect 4208 25056 4528 25057
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 34928 25056 35248 25057
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 24991 35248 24992
rect 65648 25056 65968 25057
rect 65648 24992 65656 25056
rect 65720 24992 65736 25056
rect 65800 24992 65816 25056
rect 65880 24992 65896 25056
rect 65960 24992 65968 25056
rect 65648 24991 65968 24992
rect 96368 25056 96688 25057
rect 96368 24992 96376 25056
rect 96440 24992 96456 25056
rect 96520 24992 96536 25056
rect 96600 24992 96616 25056
rect 96680 24992 96688 25056
rect 96368 24991 96688 24992
rect 127088 25056 127408 25057
rect 127088 24992 127096 25056
rect 127160 24992 127176 25056
rect 127240 24992 127256 25056
rect 127320 24992 127336 25056
rect 127400 24992 127408 25056
rect 127088 24991 127408 24992
rect 157808 25056 158128 25057
rect 157808 24992 157816 25056
rect 157880 24992 157896 25056
rect 157960 24992 157976 25056
rect 158040 24992 158056 25056
rect 158120 24992 158128 25056
rect 157808 24991 158128 24992
rect 19568 24512 19888 24513
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 24447 19888 24448
rect 50288 24512 50608 24513
rect 50288 24448 50296 24512
rect 50360 24448 50376 24512
rect 50440 24448 50456 24512
rect 50520 24448 50536 24512
rect 50600 24448 50608 24512
rect 50288 24447 50608 24448
rect 81008 24512 81328 24513
rect 81008 24448 81016 24512
rect 81080 24448 81096 24512
rect 81160 24448 81176 24512
rect 81240 24448 81256 24512
rect 81320 24448 81328 24512
rect 81008 24447 81328 24448
rect 111728 24512 112048 24513
rect 111728 24448 111736 24512
rect 111800 24448 111816 24512
rect 111880 24448 111896 24512
rect 111960 24448 111976 24512
rect 112040 24448 112048 24512
rect 111728 24447 112048 24448
rect 142448 24512 142768 24513
rect 142448 24448 142456 24512
rect 142520 24448 142536 24512
rect 142600 24448 142616 24512
rect 142680 24448 142696 24512
rect 142760 24448 142768 24512
rect 142448 24447 142768 24448
rect 173168 24512 173488 24513
rect 173168 24448 173176 24512
rect 173240 24448 173256 24512
rect 173320 24448 173336 24512
rect 173400 24448 173416 24512
rect 173480 24448 173488 24512
rect 173168 24447 173488 24448
rect 4208 23968 4528 23969
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 34928 23968 35248 23969
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 23903 35248 23904
rect 65648 23968 65968 23969
rect 65648 23904 65656 23968
rect 65720 23904 65736 23968
rect 65800 23904 65816 23968
rect 65880 23904 65896 23968
rect 65960 23904 65968 23968
rect 65648 23903 65968 23904
rect 96368 23968 96688 23969
rect 96368 23904 96376 23968
rect 96440 23904 96456 23968
rect 96520 23904 96536 23968
rect 96600 23904 96616 23968
rect 96680 23904 96688 23968
rect 96368 23903 96688 23904
rect 127088 23968 127408 23969
rect 127088 23904 127096 23968
rect 127160 23904 127176 23968
rect 127240 23904 127256 23968
rect 127320 23904 127336 23968
rect 127400 23904 127408 23968
rect 127088 23903 127408 23904
rect 157808 23968 158128 23969
rect 157808 23904 157816 23968
rect 157880 23904 157896 23968
rect 157960 23904 157976 23968
rect 158040 23904 158056 23968
rect 158120 23904 158128 23968
rect 157808 23903 158128 23904
rect 19568 23424 19888 23425
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 23359 19888 23360
rect 50288 23424 50608 23425
rect 50288 23360 50296 23424
rect 50360 23360 50376 23424
rect 50440 23360 50456 23424
rect 50520 23360 50536 23424
rect 50600 23360 50608 23424
rect 50288 23359 50608 23360
rect 81008 23424 81328 23425
rect 81008 23360 81016 23424
rect 81080 23360 81096 23424
rect 81160 23360 81176 23424
rect 81240 23360 81256 23424
rect 81320 23360 81328 23424
rect 81008 23359 81328 23360
rect 111728 23424 112048 23425
rect 111728 23360 111736 23424
rect 111800 23360 111816 23424
rect 111880 23360 111896 23424
rect 111960 23360 111976 23424
rect 112040 23360 112048 23424
rect 111728 23359 112048 23360
rect 142448 23424 142768 23425
rect 142448 23360 142456 23424
rect 142520 23360 142536 23424
rect 142600 23360 142616 23424
rect 142680 23360 142696 23424
rect 142760 23360 142768 23424
rect 142448 23359 142768 23360
rect 173168 23424 173488 23425
rect 173168 23360 173176 23424
rect 173240 23360 173256 23424
rect 173320 23360 173336 23424
rect 173400 23360 173416 23424
rect 173480 23360 173488 23424
rect 173168 23359 173488 23360
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 34928 22880 35248 22881
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 22815 35248 22816
rect 65648 22880 65968 22881
rect 65648 22816 65656 22880
rect 65720 22816 65736 22880
rect 65800 22816 65816 22880
rect 65880 22816 65896 22880
rect 65960 22816 65968 22880
rect 65648 22815 65968 22816
rect 96368 22880 96688 22881
rect 96368 22816 96376 22880
rect 96440 22816 96456 22880
rect 96520 22816 96536 22880
rect 96600 22816 96616 22880
rect 96680 22816 96688 22880
rect 96368 22815 96688 22816
rect 127088 22880 127408 22881
rect 127088 22816 127096 22880
rect 127160 22816 127176 22880
rect 127240 22816 127256 22880
rect 127320 22816 127336 22880
rect 127400 22816 127408 22880
rect 127088 22815 127408 22816
rect 157808 22880 158128 22881
rect 157808 22816 157816 22880
rect 157880 22816 157896 22880
rect 157960 22816 157976 22880
rect 158040 22816 158056 22880
rect 158120 22816 158128 22880
rect 157808 22815 158128 22816
rect 19568 22336 19888 22337
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 22271 19888 22272
rect 50288 22336 50608 22337
rect 50288 22272 50296 22336
rect 50360 22272 50376 22336
rect 50440 22272 50456 22336
rect 50520 22272 50536 22336
rect 50600 22272 50608 22336
rect 50288 22271 50608 22272
rect 81008 22336 81328 22337
rect 81008 22272 81016 22336
rect 81080 22272 81096 22336
rect 81160 22272 81176 22336
rect 81240 22272 81256 22336
rect 81320 22272 81328 22336
rect 81008 22271 81328 22272
rect 111728 22336 112048 22337
rect 111728 22272 111736 22336
rect 111800 22272 111816 22336
rect 111880 22272 111896 22336
rect 111960 22272 111976 22336
rect 112040 22272 112048 22336
rect 111728 22271 112048 22272
rect 142448 22336 142768 22337
rect 142448 22272 142456 22336
rect 142520 22272 142536 22336
rect 142600 22272 142616 22336
rect 142680 22272 142696 22336
rect 142760 22272 142768 22336
rect 142448 22271 142768 22272
rect 173168 22336 173488 22337
rect 173168 22272 173176 22336
rect 173240 22272 173256 22336
rect 173320 22272 173336 22336
rect 173400 22272 173416 22336
rect 173480 22272 173488 22336
rect 173168 22271 173488 22272
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 34928 21792 35248 21793
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 21727 35248 21728
rect 65648 21792 65968 21793
rect 65648 21728 65656 21792
rect 65720 21728 65736 21792
rect 65800 21728 65816 21792
rect 65880 21728 65896 21792
rect 65960 21728 65968 21792
rect 65648 21727 65968 21728
rect 96368 21792 96688 21793
rect 96368 21728 96376 21792
rect 96440 21728 96456 21792
rect 96520 21728 96536 21792
rect 96600 21728 96616 21792
rect 96680 21728 96688 21792
rect 96368 21727 96688 21728
rect 127088 21792 127408 21793
rect 127088 21728 127096 21792
rect 127160 21728 127176 21792
rect 127240 21728 127256 21792
rect 127320 21728 127336 21792
rect 127400 21728 127408 21792
rect 127088 21727 127408 21728
rect 157808 21792 158128 21793
rect 157808 21728 157816 21792
rect 157880 21728 157896 21792
rect 157960 21728 157976 21792
rect 158040 21728 158056 21792
rect 158120 21728 158128 21792
rect 157808 21727 158128 21728
rect 19568 21248 19888 21249
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 21183 19888 21184
rect 50288 21248 50608 21249
rect 50288 21184 50296 21248
rect 50360 21184 50376 21248
rect 50440 21184 50456 21248
rect 50520 21184 50536 21248
rect 50600 21184 50608 21248
rect 50288 21183 50608 21184
rect 81008 21248 81328 21249
rect 81008 21184 81016 21248
rect 81080 21184 81096 21248
rect 81160 21184 81176 21248
rect 81240 21184 81256 21248
rect 81320 21184 81328 21248
rect 81008 21183 81328 21184
rect 111728 21248 112048 21249
rect 111728 21184 111736 21248
rect 111800 21184 111816 21248
rect 111880 21184 111896 21248
rect 111960 21184 111976 21248
rect 112040 21184 112048 21248
rect 111728 21183 112048 21184
rect 142448 21248 142768 21249
rect 142448 21184 142456 21248
rect 142520 21184 142536 21248
rect 142600 21184 142616 21248
rect 142680 21184 142696 21248
rect 142760 21184 142768 21248
rect 142448 21183 142768 21184
rect 173168 21248 173488 21249
rect 173168 21184 173176 21248
rect 173240 21184 173256 21248
rect 173320 21184 173336 21248
rect 173400 21184 173416 21248
rect 173480 21184 173488 21248
rect 173168 21183 173488 21184
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 34928 20704 35248 20705
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 20639 35248 20640
rect 65648 20704 65968 20705
rect 65648 20640 65656 20704
rect 65720 20640 65736 20704
rect 65800 20640 65816 20704
rect 65880 20640 65896 20704
rect 65960 20640 65968 20704
rect 65648 20639 65968 20640
rect 96368 20704 96688 20705
rect 96368 20640 96376 20704
rect 96440 20640 96456 20704
rect 96520 20640 96536 20704
rect 96600 20640 96616 20704
rect 96680 20640 96688 20704
rect 96368 20639 96688 20640
rect 127088 20704 127408 20705
rect 127088 20640 127096 20704
rect 127160 20640 127176 20704
rect 127240 20640 127256 20704
rect 127320 20640 127336 20704
rect 127400 20640 127408 20704
rect 127088 20639 127408 20640
rect 157808 20704 158128 20705
rect 157808 20640 157816 20704
rect 157880 20640 157896 20704
rect 157960 20640 157976 20704
rect 158040 20640 158056 20704
rect 158120 20640 158128 20704
rect 157808 20639 158128 20640
rect 19568 20160 19888 20161
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 20095 19888 20096
rect 50288 20160 50608 20161
rect 50288 20096 50296 20160
rect 50360 20096 50376 20160
rect 50440 20096 50456 20160
rect 50520 20096 50536 20160
rect 50600 20096 50608 20160
rect 50288 20095 50608 20096
rect 81008 20160 81328 20161
rect 81008 20096 81016 20160
rect 81080 20096 81096 20160
rect 81160 20096 81176 20160
rect 81240 20096 81256 20160
rect 81320 20096 81328 20160
rect 81008 20095 81328 20096
rect 111728 20160 112048 20161
rect 111728 20096 111736 20160
rect 111800 20096 111816 20160
rect 111880 20096 111896 20160
rect 111960 20096 111976 20160
rect 112040 20096 112048 20160
rect 111728 20095 112048 20096
rect 142448 20160 142768 20161
rect 142448 20096 142456 20160
rect 142520 20096 142536 20160
rect 142600 20096 142616 20160
rect 142680 20096 142696 20160
rect 142760 20096 142768 20160
rect 142448 20095 142768 20096
rect 173168 20160 173488 20161
rect 173168 20096 173176 20160
rect 173240 20096 173256 20160
rect 173320 20096 173336 20160
rect 173400 20096 173416 20160
rect 173480 20096 173488 20160
rect 173168 20095 173488 20096
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 34928 19616 35248 19617
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 19551 35248 19552
rect 65648 19616 65968 19617
rect 65648 19552 65656 19616
rect 65720 19552 65736 19616
rect 65800 19552 65816 19616
rect 65880 19552 65896 19616
rect 65960 19552 65968 19616
rect 65648 19551 65968 19552
rect 96368 19616 96688 19617
rect 96368 19552 96376 19616
rect 96440 19552 96456 19616
rect 96520 19552 96536 19616
rect 96600 19552 96616 19616
rect 96680 19552 96688 19616
rect 96368 19551 96688 19552
rect 127088 19616 127408 19617
rect 127088 19552 127096 19616
rect 127160 19552 127176 19616
rect 127240 19552 127256 19616
rect 127320 19552 127336 19616
rect 127400 19552 127408 19616
rect 127088 19551 127408 19552
rect 157808 19616 158128 19617
rect 157808 19552 157816 19616
rect 157880 19552 157896 19616
rect 157960 19552 157976 19616
rect 158040 19552 158056 19616
rect 158120 19552 158128 19616
rect 157808 19551 158128 19552
rect 19568 19072 19888 19073
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 19007 19888 19008
rect 50288 19072 50608 19073
rect 50288 19008 50296 19072
rect 50360 19008 50376 19072
rect 50440 19008 50456 19072
rect 50520 19008 50536 19072
rect 50600 19008 50608 19072
rect 50288 19007 50608 19008
rect 81008 19072 81328 19073
rect 81008 19008 81016 19072
rect 81080 19008 81096 19072
rect 81160 19008 81176 19072
rect 81240 19008 81256 19072
rect 81320 19008 81328 19072
rect 81008 19007 81328 19008
rect 111728 19072 112048 19073
rect 111728 19008 111736 19072
rect 111800 19008 111816 19072
rect 111880 19008 111896 19072
rect 111960 19008 111976 19072
rect 112040 19008 112048 19072
rect 111728 19007 112048 19008
rect 142448 19072 142768 19073
rect 142448 19008 142456 19072
rect 142520 19008 142536 19072
rect 142600 19008 142616 19072
rect 142680 19008 142696 19072
rect 142760 19008 142768 19072
rect 142448 19007 142768 19008
rect 173168 19072 173488 19073
rect 173168 19008 173176 19072
rect 173240 19008 173256 19072
rect 173320 19008 173336 19072
rect 173400 19008 173416 19072
rect 173480 19008 173488 19072
rect 173168 19007 173488 19008
rect 4208 18528 4528 18529
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 34928 18528 35248 18529
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 18463 35248 18464
rect 65648 18528 65968 18529
rect 65648 18464 65656 18528
rect 65720 18464 65736 18528
rect 65800 18464 65816 18528
rect 65880 18464 65896 18528
rect 65960 18464 65968 18528
rect 65648 18463 65968 18464
rect 96368 18528 96688 18529
rect 96368 18464 96376 18528
rect 96440 18464 96456 18528
rect 96520 18464 96536 18528
rect 96600 18464 96616 18528
rect 96680 18464 96688 18528
rect 96368 18463 96688 18464
rect 127088 18528 127408 18529
rect 127088 18464 127096 18528
rect 127160 18464 127176 18528
rect 127240 18464 127256 18528
rect 127320 18464 127336 18528
rect 127400 18464 127408 18528
rect 127088 18463 127408 18464
rect 157808 18528 158128 18529
rect 157808 18464 157816 18528
rect 157880 18464 157896 18528
rect 157960 18464 157976 18528
rect 158040 18464 158056 18528
rect 158120 18464 158128 18528
rect 157808 18463 158128 18464
rect 19568 17984 19888 17985
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 17919 19888 17920
rect 50288 17984 50608 17985
rect 50288 17920 50296 17984
rect 50360 17920 50376 17984
rect 50440 17920 50456 17984
rect 50520 17920 50536 17984
rect 50600 17920 50608 17984
rect 50288 17919 50608 17920
rect 81008 17984 81328 17985
rect 81008 17920 81016 17984
rect 81080 17920 81096 17984
rect 81160 17920 81176 17984
rect 81240 17920 81256 17984
rect 81320 17920 81328 17984
rect 81008 17919 81328 17920
rect 111728 17984 112048 17985
rect 111728 17920 111736 17984
rect 111800 17920 111816 17984
rect 111880 17920 111896 17984
rect 111960 17920 111976 17984
rect 112040 17920 112048 17984
rect 111728 17919 112048 17920
rect 142448 17984 142768 17985
rect 142448 17920 142456 17984
rect 142520 17920 142536 17984
rect 142600 17920 142616 17984
rect 142680 17920 142696 17984
rect 142760 17920 142768 17984
rect 142448 17919 142768 17920
rect 173168 17984 173488 17985
rect 173168 17920 173176 17984
rect 173240 17920 173256 17984
rect 173320 17920 173336 17984
rect 173400 17920 173416 17984
rect 173480 17920 173488 17984
rect 173168 17919 173488 17920
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 34928 17440 35248 17441
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 17375 35248 17376
rect 65648 17440 65968 17441
rect 65648 17376 65656 17440
rect 65720 17376 65736 17440
rect 65800 17376 65816 17440
rect 65880 17376 65896 17440
rect 65960 17376 65968 17440
rect 65648 17375 65968 17376
rect 96368 17440 96688 17441
rect 96368 17376 96376 17440
rect 96440 17376 96456 17440
rect 96520 17376 96536 17440
rect 96600 17376 96616 17440
rect 96680 17376 96688 17440
rect 96368 17375 96688 17376
rect 127088 17440 127408 17441
rect 127088 17376 127096 17440
rect 127160 17376 127176 17440
rect 127240 17376 127256 17440
rect 127320 17376 127336 17440
rect 127400 17376 127408 17440
rect 127088 17375 127408 17376
rect 157808 17440 158128 17441
rect 157808 17376 157816 17440
rect 157880 17376 157896 17440
rect 157960 17376 157976 17440
rect 158040 17376 158056 17440
rect 158120 17376 158128 17440
rect 157808 17375 158128 17376
rect 19568 16896 19888 16897
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 16831 19888 16832
rect 50288 16896 50608 16897
rect 50288 16832 50296 16896
rect 50360 16832 50376 16896
rect 50440 16832 50456 16896
rect 50520 16832 50536 16896
rect 50600 16832 50608 16896
rect 50288 16831 50608 16832
rect 81008 16896 81328 16897
rect 81008 16832 81016 16896
rect 81080 16832 81096 16896
rect 81160 16832 81176 16896
rect 81240 16832 81256 16896
rect 81320 16832 81328 16896
rect 81008 16831 81328 16832
rect 111728 16896 112048 16897
rect 111728 16832 111736 16896
rect 111800 16832 111816 16896
rect 111880 16832 111896 16896
rect 111960 16832 111976 16896
rect 112040 16832 112048 16896
rect 111728 16831 112048 16832
rect 142448 16896 142768 16897
rect 142448 16832 142456 16896
rect 142520 16832 142536 16896
rect 142600 16832 142616 16896
rect 142680 16832 142696 16896
rect 142760 16832 142768 16896
rect 142448 16831 142768 16832
rect 173168 16896 173488 16897
rect 173168 16832 173176 16896
rect 173240 16832 173256 16896
rect 173320 16832 173336 16896
rect 173400 16832 173416 16896
rect 173480 16832 173488 16896
rect 173168 16831 173488 16832
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 34928 16352 35248 16353
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 16287 35248 16288
rect 65648 16352 65968 16353
rect 65648 16288 65656 16352
rect 65720 16288 65736 16352
rect 65800 16288 65816 16352
rect 65880 16288 65896 16352
rect 65960 16288 65968 16352
rect 65648 16287 65968 16288
rect 96368 16352 96688 16353
rect 96368 16288 96376 16352
rect 96440 16288 96456 16352
rect 96520 16288 96536 16352
rect 96600 16288 96616 16352
rect 96680 16288 96688 16352
rect 96368 16287 96688 16288
rect 127088 16352 127408 16353
rect 127088 16288 127096 16352
rect 127160 16288 127176 16352
rect 127240 16288 127256 16352
rect 127320 16288 127336 16352
rect 127400 16288 127408 16352
rect 127088 16287 127408 16288
rect 157808 16352 158128 16353
rect 157808 16288 157816 16352
rect 157880 16288 157896 16352
rect 157960 16288 157976 16352
rect 158040 16288 158056 16352
rect 158120 16288 158128 16352
rect 157808 16287 158128 16288
rect 19568 15808 19888 15809
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 15743 19888 15744
rect 50288 15808 50608 15809
rect 50288 15744 50296 15808
rect 50360 15744 50376 15808
rect 50440 15744 50456 15808
rect 50520 15744 50536 15808
rect 50600 15744 50608 15808
rect 50288 15743 50608 15744
rect 81008 15808 81328 15809
rect 81008 15744 81016 15808
rect 81080 15744 81096 15808
rect 81160 15744 81176 15808
rect 81240 15744 81256 15808
rect 81320 15744 81328 15808
rect 81008 15743 81328 15744
rect 111728 15808 112048 15809
rect 111728 15744 111736 15808
rect 111800 15744 111816 15808
rect 111880 15744 111896 15808
rect 111960 15744 111976 15808
rect 112040 15744 112048 15808
rect 111728 15743 112048 15744
rect 142448 15808 142768 15809
rect 142448 15744 142456 15808
rect 142520 15744 142536 15808
rect 142600 15744 142616 15808
rect 142680 15744 142696 15808
rect 142760 15744 142768 15808
rect 142448 15743 142768 15744
rect 173168 15808 173488 15809
rect 173168 15744 173176 15808
rect 173240 15744 173256 15808
rect 173320 15744 173336 15808
rect 173400 15744 173416 15808
rect 173480 15744 173488 15808
rect 173168 15743 173488 15744
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 34928 15264 35248 15265
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 15199 35248 15200
rect 65648 15264 65968 15265
rect 65648 15200 65656 15264
rect 65720 15200 65736 15264
rect 65800 15200 65816 15264
rect 65880 15200 65896 15264
rect 65960 15200 65968 15264
rect 65648 15199 65968 15200
rect 96368 15264 96688 15265
rect 96368 15200 96376 15264
rect 96440 15200 96456 15264
rect 96520 15200 96536 15264
rect 96600 15200 96616 15264
rect 96680 15200 96688 15264
rect 96368 15199 96688 15200
rect 127088 15264 127408 15265
rect 127088 15200 127096 15264
rect 127160 15200 127176 15264
rect 127240 15200 127256 15264
rect 127320 15200 127336 15264
rect 127400 15200 127408 15264
rect 127088 15199 127408 15200
rect 157808 15264 158128 15265
rect 157808 15200 157816 15264
rect 157880 15200 157896 15264
rect 157960 15200 157976 15264
rect 158040 15200 158056 15264
rect 158120 15200 158128 15264
rect 157808 15199 158128 15200
rect 19568 14720 19888 14721
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 14655 19888 14656
rect 50288 14720 50608 14721
rect 50288 14656 50296 14720
rect 50360 14656 50376 14720
rect 50440 14656 50456 14720
rect 50520 14656 50536 14720
rect 50600 14656 50608 14720
rect 50288 14655 50608 14656
rect 81008 14720 81328 14721
rect 81008 14656 81016 14720
rect 81080 14656 81096 14720
rect 81160 14656 81176 14720
rect 81240 14656 81256 14720
rect 81320 14656 81328 14720
rect 81008 14655 81328 14656
rect 111728 14720 112048 14721
rect 111728 14656 111736 14720
rect 111800 14656 111816 14720
rect 111880 14656 111896 14720
rect 111960 14656 111976 14720
rect 112040 14656 112048 14720
rect 111728 14655 112048 14656
rect 142448 14720 142768 14721
rect 142448 14656 142456 14720
rect 142520 14656 142536 14720
rect 142600 14656 142616 14720
rect 142680 14656 142696 14720
rect 142760 14656 142768 14720
rect 142448 14655 142768 14656
rect 173168 14720 173488 14721
rect 173168 14656 173176 14720
rect 173240 14656 173256 14720
rect 173320 14656 173336 14720
rect 173400 14656 173416 14720
rect 173480 14656 173488 14720
rect 173168 14655 173488 14656
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 34928 14176 35248 14177
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 14111 35248 14112
rect 65648 14176 65968 14177
rect 65648 14112 65656 14176
rect 65720 14112 65736 14176
rect 65800 14112 65816 14176
rect 65880 14112 65896 14176
rect 65960 14112 65968 14176
rect 65648 14111 65968 14112
rect 96368 14176 96688 14177
rect 96368 14112 96376 14176
rect 96440 14112 96456 14176
rect 96520 14112 96536 14176
rect 96600 14112 96616 14176
rect 96680 14112 96688 14176
rect 96368 14111 96688 14112
rect 127088 14176 127408 14177
rect 127088 14112 127096 14176
rect 127160 14112 127176 14176
rect 127240 14112 127256 14176
rect 127320 14112 127336 14176
rect 127400 14112 127408 14176
rect 127088 14111 127408 14112
rect 157808 14176 158128 14177
rect 157808 14112 157816 14176
rect 157880 14112 157896 14176
rect 157960 14112 157976 14176
rect 158040 14112 158056 14176
rect 158120 14112 158128 14176
rect 157808 14111 158128 14112
rect 19568 13632 19888 13633
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 13567 19888 13568
rect 50288 13632 50608 13633
rect 50288 13568 50296 13632
rect 50360 13568 50376 13632
rect 50440 13568 50456 13632
rect 50520 13568 50536 13632
rect 50600 13568 50608 13632
rect 50288 13567 50608 13568
rect 81008 13632 81328 13633
rect 81008 13568 81016 13632
rect 81080 13568 81096 13632
rect 81160 13568 81176 13632
rect 81240 13568 81256 13632
rect 81320 13568 81328 13632
rect 81008 13567 81328 13568
rect 111728 13632 112048 13633
rect 111728 13568 111736 13632
rect 111800 13568 111816 13632
rect 111880 13568 111896 13632
rect 111960 13568 111976 13632
rect 112040 13568 112048 13632
rect 111728 13567 112048 13568
rect 142448 13632 142768 13633
rect 142448 13568 142456 13632
rect 142520 13568 142536 13632
rect 142600 13568 142616 13632
rect 142680 13568 142696 13632
rect 142760 13568 142768 13632
rect 142448 13567 142768 13568
rect 173168 13632 173488 13633
rect 173168 13568 173176 13632
rect 173240 13568 173256 13632
rect 173320 13568 173336 13632
rect 173400 13568 173416 13632
rect 173480 13568 173488 13632
rect 173168 13567 173488 13568
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 34928 13088 35248 13089
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 13023 35248 13024
rect 65648 13088 65968 13089
rect 65648 13024 65656 13088
rect 65720 13024 65736 13088
rect 65800 13024 65816 13088
rect 65880 13024 65896 13088
rect 65960 13024 65968 13088
rect 65648 13023 65968 13024
rect 96368 13088 96688 13089
rect 96368 13024 96376 13088
rect 96440 13024 96456 13088
rect 96520 13024 96536 13088
rect 96600 13024 96616 13088
rect 96680 13024 96688 13088
rect 96368 13023 96688 13024
rect 127088 13088 127408 13089
rect 127088 13024 127096 13088
rect 127160 13024 127176 13088
rect 127240 13024 127256 13088
rect 127320 13024 127336 13088
rect 127400 13024 127408 13088
rect 127088 13023 127408 13024
rect 157808 13088 158128 13089
rect 157808 13024 157816 13088
rect 157880 13024 157896 13088
rect 157960 13024 157976 13088
rect 158040 13024 158056 13088
rect 158120 13024 158128 13088
rect 157808 13023 158128 13024
rect 19568 12544 19888 12545
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 12479 19888 12480
rect 50288 12544 50608 12545
rect 50288 12480 50296 12544
rect 50360 12480 50376 12544
rect 50440 12480 50456 12544
rect 50520 12480 50536 12544
rect 50600 12480 50608 12544
rect 50288 12479 50608 12480
rect 81008 12544 81328 12545
rect 81008 12480 81016 12544
rect 81080 12480 81096 12544
rect 81160 12480 81176 12544
rect 81240 12480 81256 12544
rect 81320 12480 81328 12544
rect 81008 12479 81328 12480
rect 111728 12544 112048 12545
rect 111728 12480 111736 12544
rect 111800 12480 111816 12544
rect 111880 12480 111896 12544
rect 111960 12480 111976 12544
rect 112040 12480 112048 12544
rect 111728 12479 112048 12480
rect 142448 12544 142768 12545
rect 142448 12480 142456 12544
rect 142520 12480 142536 12544
rect 142600 12480 142616 12544
rect 142680 12480 142696 12544
rect 142760 12480 142768 12544
rect 142448 12479 142768 12480
rect 173168 12544 173488 12545
rect 173168 12480 173176 12544
rect 173240 12480 173256 12544
rect 173320 12480 173336 12544
rect 173400 12480 173416 12544
rect 173480 12480 173488 12544
rect 173168 12479 173488 12480
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 34928 12000 35248 12001
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 11935 35248 11936
rect 65648 12000 65968 12001
rect 65648 11936 65656 12000
rect 65720 11936 65736 12000
rect 65800 11936 65816 12000
rect 65880 11936 65896 12000
rect 65960 11936 65968 12000
rect 65648 11935 65968 11936
rect 96368 12000 96688 12001
rect 96368 11936 96376 12000
rect 96440 11936 96456 12000
rect 96520 11936 96536 12000
rect 96600 11936 96616 12000
rect 96680 11936 96688 12000
rect 96368 11935 96688 11936
rect 127088 12000 127408 12001
rect 127088 11936 127096 12000
rect 127160 11936 127176 12000
rect 127240 11936 127256 12000
rect 127320 11936 127336 12000
rect 127400 11936 127408 12000
rect 127088 11935 127408 11936
rect 157808 12000 158128 12001
rect 157808 11936 157816 12000
rect 157880 11936 157896 12000
rect 157960 11936 157976 12000
rect 158040 11936 158056 12000
rect 158120 11936 158128 12000
rect 157808 11935 158128 11936
rect 19568 11456 19888 11457
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 11391 19888 11392
rect 50288 11456 50608 11457
rect 50288 11392 50296 11456
rect 50360 11392 50376 11456
rect 50440 11392 50456 11456
rect 50520 11392 50536 11456
rect 50600 11392 50608 11456
rect 50288 11391 50608 11392
rect 81008 11456 81328 11457
rect 81008 11392 81016 11456
rect 81080 11392 81096 11456
rect 81160 11392 81176 11456
rect 81240 11392 81256 11456
rect 81320 11392 81328 11456
rect 81008 11391 81328 11392
rect 111728 11456 112048 11457
rect 111728 11392 111736 11456
rect 111800 11392 111816 11456
rect 111880 11392 111896 11456
rect 111960 11392 111976 11456
rect 112040 11392 112048 11456
rect 111728 11391 112048 11392
rect 142448 11456 142768 11457
rect 142448 11392 142456 11456
rect 142520 11392 142536 11456
rect 142600 11392 142616 11456
rect 142680 11392 142696 11456
rect 142760 11392 142768 11456
rect 142448 11391 142768 11392
rect 173168 11456 173488 11457
rect 173168 11392 173176 11456
rect 173240 11392 173256 11456
rect 173320 11392 173336 11456
rect 173400 11392 173416 11456
rect 173480 11392 173488 11456
rect 173168 11391 173488 11392
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 34928 10912 35248 10913
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 10847 35248 10848
rect 65648 10912 65968 10913
rect 65648 10848 65656 10912
rect 65720 10848 65736 10912
rect 65800 10848 65816 10912
rect 65880 10848 65896 10912
rect 65960 10848 65968 10912
rect 65648 10847 65968 10848
rect 96368 10912 96688 10913
rect 96368 10848 96376 10912
rect 96440 10848 96456 10912
rect 96520 10848 96536 10912
rect 96600 10848 96616 10912
rect 96680 10848 96688 10912
rect 96368 10847 96688 10848
rect 127088 10912 127408 10913
rect 127088 10848 127096 10912
rect 127160 10848 127176 10912
rect 127240 10848 127256 10912
rect 127320 10848 127336 10912
rect 127400 10848 127408 10912
rect 127088 10847 127408 10848
rect 157808 10912 158128 10913
rect 157808 10848 157816 10912
rect 157880 10848 157896 10912
rect 157960 10848 157976 10912
rect 158040 10848 158056 10912
rect 158120 10848 158128 10912
rect 157808 10847 158128 10848
rect 19568 10368 19888 10369
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 10303 19888 10304
rect 50288 10368 50608 10369
rect 50288 10304 50296 10368
rect 50360 10304 50376 10368
rect 50440 10304 50456 10368
rect 50520 10304 50536 10368
rect 50600 10304 50608 10368
rect 50288 10303 50608 10304
rect 81008 10368 81328 10369
rect 81008 10304 81016 10368
rect 81080 10304 81096 10368
rect 81160 10304 81176 10368
rect 81240 10304 81256 10368
rect 81320 10304 81328 10368
rect 81008 10303 81328 10304
rect 111728 10368 112048 10369
rect 111728 10304 111736 10368
rect 111800 10304 111816 10368
rect 111880 10304 111896 10368
rect 111960 10304 111976 10368
rect 112040 10304 112048 10368
rect 111728 10303 112048 10304
rect 142448 10368 142768 10369
rect 142448 10304 142456 10368
rect 142520 10304 142536 10368
rect 142600 10304 142616 10368
rect 142680 10304 142696 10368
rect 142760 10304 142768 10368
rect 142448 10303 142768 10304
rect 173168 10368 173488 10369
rect 173168 10304 173176 10368
rect 173240 10304 173256 10368
rect 173320 10304 173336 10368
rect 173400 10304 173416 10368
rect 173480 10304 173488 10368
rect 173168 10303 173488 10304
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 34928 9824 35248 9825
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 9759 35248 9760
rect 65648 9824 65968 9825
rect 65648 9760 65656 9824
rect 65720 9760 65736 9824
rect 65800 9760 65816 9824
rect 65880 9760 65896 9824
rect 65960 9760 65968 9824
rect 65648 9759 65968 9760
rect 96368 9824 96688 9825
rect 96368 9760 96376 9824
rect 96440 9760 96456 9824
rect 96520 9760 96536 9824
rect 96600 9760 96616 9824
rect 96680 9760 96688 9824
rect 96368 9759 96688 9760
rect 127088 9824 127408 9825
rect 127088 9760 127096 9824
rect 127160 9760 127176 9824
rect 127240 9760 127256 9824
rect 127320 9760 127336 9824
rect 127400 9760 127408 9824
rect 127088 9759 127408 9760
rect 157808 9824 158128 9825
rect 157808 9760 157816 9824
rect 157880 9760 157896 9824
rect 157960 9760 157976 9824
rect 158040 9760 158056 9824
rect 158120 9760 158128 9824
rect 157808 9759 158128 9760
rect 19568 9280 19888 9281
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 9215 19888 9216
rect 50288 9280 50608 9281
rect 50288 9216 50296 9280
rect 50360 9216 50376 9280
rect 50440 9216 50456 9280
rect 50520 9216 50536 9280
rect 50600 9216 50608 9280
rect 50288 9215 50608 9216
rect 81008 9280 81328 9281
rect 81008 9216 81016 9280
rect 81080 9216 81096 9280
rect 81160 9216 81176 9280
rect 81240 9216 81256 9280
rect 81320 9216 81328 9280
rect 81008 9215 81328 9216
rect 111728 9280 112048 9281
rect 111728 9216 111736 9280
rect 111800 9216 111816 9280
rect 111880 9216 111896 9280
rect 111960 9216 111976 9280
rect 112040 9216 112048 9280
rect 111728 9215 112048 9216
rect 142448 9280 142768 9281
rect 142448 9216 142456 9280
rect 142520 9216 142536 9280
rect 142600 9216 142616 9280
rect 142680 9216 142696 9280
rect 142760 9216 142768 9280
rect 142448 9215 142768 9216
rect 173168 9280 173488 9281
rect 173168 9216 173176 9280
rect 173240 9216 173256 9280
rect 173320 9216 173336 9280
rect 173400 9216 173416 9280
rect 173480 9216 173488 9280
rect 173168 9215 173488 9216
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 34928 8736 35248 8737
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 8671 35248 8672
rect 65648 8736 65968 8737
rect 65648 8672 65656 8736
rect 65720 8672 65736 8736
rect 65800 8672 65816 8736
rect 65880 8672 65896 8736
rect 65960 8672 65968 8736
rect 65648 8671 65968 8672
rect 96368 8736 96688 8737
rect 96368 8672 96376 8736
rect 96440 8672 96456 8736
rect 96520 8672 96536 8736
rect 96600 8672 96616 8736
rect 96680 8672 96688 8736
rect 96368 8671 96688 8672
rect 127088 8736 127408 8737
rect 127088 8672 127096 8736
rect 127160 8672 127176 8736
rect 127240 8672 127256 8736
rect 127320 8672 127336 8736
rect 127400 8672 127408 8736
rect 127088 8671 127408 8672
rect 157808 8736 158128 8737
rect 157808 8672 157816 8736
rect 157880 8672 157896 8736
rect 157960 8672 157976 8736
rect 158040 8672 158056 8736
rect 158120 8672 158128 8736
rect 157808 8671 158128 8672
rect 39113 8258 39179 8261
rect 46013 8258 46079 8261
rect 46381 8258 46447 8261
rect 47301 8258 47367 8261
rect 39113 8256 47367 8258
rect 39113 8200 39118 8256
rect 39174 8200 46018 8256
rect 46074 8200 46386 8256
rect 46442 8200 47306 8256
rect 47362 8200 47367 8256
rect 39113 8198 47367 8200
rect 39113 8195 39179 8198
rect 46013 8195 46079 8198
rect 46381 8195 46447 8198
rect 47301 8195 47367 8198
rect 19568 8192 19888 8193
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 8127 19888 8128
rect 50288 8192 50608 8193
rect 50288 8128 50296 8192
rect 50360 8128 50376 8192
rect 50440 8128 50456 8192
rect 50520 8128 50536 8192
rect 50600 8128 50608 8192
rect 50288 8127 50608 8128
rect 81008 8192 81328 8193
rect 81008 8128 81016 8192
rect 81080 8128 81096 8192
rect 81160 8128 81176 8192
rect 81240 8128 81256 8192
rect 81320 8128 81328 8192
rect 81008 8127 81328 8128
rect 111728 8192 112048 8193
rect 111728 8128 111736 8192
rect 111800 8128 111816 8192
rect 111880 8128 111896 8192
rect 111960 8128 111976 8192
rect 112040 8128 112048 8192
rect 111728 8127 112048 8128
rect 142448 8192 142768 8193
rect 142448 8128 142456 8192
rect 142520 8128 142536 8192
rect 142600 8128 142616 8192
rect 142680 8128 142696 8192
rect 142760 8128 142768 8192
rect 142448 8127 142768 8128
rect 173168 8192 173488 8193
rect 173168 8128 173176 8192
rect 173240 8128 173256 8192
rect 173320 8128 173336 8192
rect 173400 8128 173416 8192
rect 173480 8128 173488 8192
rect 173168 8127 173488 8128
rect 32489 8122 32555 8125
rect 32949 8122 33015 8125
rect 32489 8120 33015 8122
rect 32489 8064 32494 8120
rect 32550 8064 32954 8120
rect 33010 8064 33015 8120
rect 32489 8062 33015 8064
rect 32489 8059 32555 8062
rect 32949 8059 33015 8062
rect 38653 8122 38719 8125
rect 39941 8122 40007 8125
rect 41229 8122 41295 8125
rect 38653 8120 41295 8122
rect 38653 8064 38658 8120
rect 38714 8064 39946 8120
rect 40002 8064 41234 8120
rect 41290 8064 41295 8120
rect 38653 8062 41295 8064
rect 38653 8059 38719 8062
rect 39941 8059 40007 8062
rect 41229 8059 41295 8062
rect 41597 8122 41663 8125
rect 47393 8122 47459 8125
rect 41597 8120 47459 8122
rect 41597 8064 41602 8120
rect 41658 8064 47398 8120
rect 47454 8064 47459 8120
rect 41597 8062 47459 8064
rect 41597 8059 41663 8062
rect 47393 8059 47459 8062
rect 20989 7986 21055 7989
rect 28165 7986 28231 7989
rect 20989 7984 28231 7986
rect 20989 7928 20994 7984
rect 21050 7928 28170 7984
rect 28226 7928 28231 7984
rect 20989 7926 28231 7928
rect 20989 7923 21055 7926
rect 28165 7923 28231 7926
rect 32765 7986 32831 7989
rect 39205 7986 39271 7989
rect 44173 7986 44239 7989
rect 32765 7984 44239 7986
rect 32765 7928 32770 7984
rect 32826 7928 39210 7984
rect 39266 7928 44178 7984
rect 44234 7928 44239 7984
rect 32765 7926 44239 7928
rect 32765 7923 32831 7926
rect 39205 7923 39271 7926
rect 44173 7923 44239 7926
rect 46013 7986 46079 7989
rect 47945 7986 48011 7989
rect 46013 7984 48011 7986
rect 46013 7928 46018 7984
rect 46074 7928 47950 7984
rect 48006 7928 48011 7984
rect 46013 7926 48011 7928
rect 46013 7923 46079 7926
rect 47945 7923 48011 7926
rect 48497 7986 48563 7989
rect 55857 7986 55923 7989
rect 48497 7984 55923 7986
rect 48497 7928 48502 7984
rect 48558 7928 55862 7984
rect 55918 7928 55923 7984
rect 48497 7926 55923 7928
rect 48497 7923 48563 7926
rect 55857 7923 55923 7926
rect 41045 7850 41111 7853
rect 42793 7850 42859 7853
rect 41045 7848 42859 7850
rect 41045 7792 41050 7848
rect 41106 7792 42798 7848
rect 42854 7792 42859 7848
rect 41045 7790 42859 7792
rect 41045 7787 41111 7790
rect 42793 7787 42859 7790
rect 46289 7850 46355 7853
rect 48681 7850 48747 7853
rect 46289 7848 48747 7850
rect 46289 7792 46294 7848
rect 46350 7792 48686 7848
rect 48742 7792 48747 7848
rect 46289 7790 48747 7792
rect 46289 7787 46355 7790
rect 48681 7787 48747 7790
rect 62573 7850 62639 7853
rect 64229 7850 64295 7853
rect 62573 7848 64295 7850
rect 62573 7792 62578 7848
rect 62634 7792 64234 7848
rect 64290 7792 64295 7848
rect 62573 7790 64295 7792
rect 62573 7787 62639 7790
rect 64229 7787 64295 7790
rect 28533 7714 28599 7717
rect 33961 7714 34027 7717
rect 28533 7712 34027 7714
rect 28533 7656 28538 7712
rect 28594 7656 33966 7712
rect 34022 7656 34027 7712
rect 28533 7654 34027 7656
rect 28533 7651 28599 7654
rect 33961 7651 34027 7654
rect 41873 7714 41939 7717
rect 46933 7714 46999 7717
rect 41873 7712 46999 7714
rect 41873 7656 41878 7712
rect 41934 7656 46938 7712
rect 46994 7656 46999 7712
rect 41873 7654 46999 7656
rect 41873 7651 41939 7654
rect 46933 7651 46999 7654
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 34928 7648 35248 7649
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 7583 35248 7584
rect 65648 7648 65968 7649
rect 65648 7584 65656 7648
rect 65720 7584 65736 7648
rect 65800 7584 65816 7648
rect 65880 7584 65896 7648
rect 65960 7584 65968 7648
rect 65648 7583 65968 7584
rect 96368 7648 96688 7649
rect 96368 7584 96376 7648
rect 96440 7584 96456 7648
rect 96520 7584 96536 7648
rect 96600 7584 96616 7648
rect 96680 7584 96688 7648
rect 96368 7583 96688 7584
rect 127088 7648 127408 7649
rect 127088 7584 127096 7648
rect 127160 7584 127176 7648
rect 127240 7584 127256 7648
rect 127320 7584 127336 7648
rect 127400 7584 127408 7648
rect 127088 7583 127408 7584
rect 157808 7648 158128 7649
rect 157808 7584 157816 7648
rect 157880 7584 157896 7648
rect 157960 7584 157976 7648
rect 158040 7584 158056 7648
rect 158120 7584 158128 7648
rect 157808 7583 158128 7584
rect 22185 7578 22251 7581
rect 28901 7578 28967 7581
rect 22185 7576 28967 7578
rect 22185 7520 22190 7576
rect 22246 7520 28906 7576
rect 28962 7520 28967 7576
rect 22185 7518 28967 7520
rect 22185 7515 22251 7518
rect 28901 7515 28967 7518
rect 39481 7578 39547 7581
rect 41505 7578 41571 7581
rect 39481 7576 41571 7578
rect 39481 7520 39486 7576
rect 39542 7520 41510 7576
rect 41566 7520 41571 7576
rect 39481 7518 41571 7520
rect 39481 7515 39547 7518
rect 41505 7515 41571 7518
rect 47209 7578 47275 7581
rect 49325 7578 49391 7581
rect 47209 7576 49391 7578
rect 47209 7520 47214 7576
rect 47270 7520 49330 7576
rect 49386 7520 49391 7576
rect 47209 7518 49391 7520
rect 47209 7515 47275 7518
rect 49325 7515 49391 7518
rect 26509 7442 26575 7445
rect 36169 7442 36235 7445
rect 26509 7440 36235 7442
rect 26509 7384 26514 7440
rect 26570 7384 36174 7440
rect 36230 7384 36235 7440
rect 26509 7382 36235 7384
rect 26509 7379 26575 7382
rect 36169 7379 36235 7382
rect 39389 7442 39455 7445
rect 42333 7442 42399 7445
rect 42609 7442 42675 7445
rect 39389 7440 42675 7442
rect 39389 7384 39394 7440
rect 39450 7384 42338 7440
rect 42394 7384 42614 7440
rect 42670 7384 42675 7440
rect 39389 7382 42675 7384
rect 39389 7379 39455 7382
rect 42333 7379 42399 7382
rect 42609 7379 42675 7382
rect 46933 7442 46999 7445
rect 49233 7442 49299 7445
rect 46933 7440 49299 7442
rect 46933 7384 46938 7440
rect 46994 7384 49238 7440
rect 49294 7384 49299 7440
rect 46933 7382 49299 7384
rect 46933 7379 46999 7382
rect 49233 7379 49299 7382
rect 50889 7442 50955 7445
rect 51073 7442 51139 7445
rect 50889 7440 51139 7442
rect 50889 7384 50894 7440
rect 50950 7384 51078 7440
rect 51134 7384 51139 7440
rect 50889 7382 51139 7384
rect 50889 7379 50955 7382
rect 51073 7379 51139 7382
rect 62297 7442 62363 7445
rect 63309 7442 63375 7445
rect 62297 7440 63375 7442
rect 62297 7384 62302 7440
rect 62358 7384 63314 7440
rect 63370 7384 63375 7440
rect 62297 7382 63375 7384
rect 62297 7379 62363 7382
rect 63309 7379 63375 7382
rect 28441 7306 28507 7309
rect 29637 7306 29703 7309
rect 28441 7304 29703 7306
rect 28441 7248 28446 7304
rect 28502 7248 29642 7304
rect 29698 7248 29703 7304
rect 28441 7246 29703 7248
rect 28441 7243 28507 7246
rect 29637 7243 29703 7246
rect 30465 7306 30531 7309
rect 31293 7306 31359 7309
rect 30465 7304 31359 7306
rect 30465 7248 30470 7304
rect 30526 7248 31298 7304
rect 31354 7248 31359 7304
rect 30465 7246 31359 7248
rect 30465 7243 30531 7246
rect 31293 7243 31359 7246
rect 34237 7306 34303 7309
rect 35249 7306 35315 7309
rect 34237 7304 35315 7306
rect 34237 7248 34242 7304
rect 34298 7248 35254 7304
rect 35310 7248 35315 7304
rect 34237 7246 35315 7248
rect 34237 7243 34303 7246
rect 35249 7243 35315 7246
rect 41689 7306 41755 7309
rect 43621 7306 43687 7309
rect 41689 7304 43687 7306
rect 41689 7248 41694 7304
rect 41750 7248 43626 7304
rect 43682 7248 43687 7304
rect 41689 7246 43687 7248
rect 41689 7243 41755 7246
rect 43621 7243 43687 7246
rect 61561 7306 61627 7309
rect 63861 7306 63927 7309
rect 61561 7304 63927 7306
rect 61561 7248 61566 7304
rect 61622 7248 63866 7304
rect 63922 7248 63927 7304
rect 61561 7246 63927 7248
rect 61561 7243 61627 7246
rect 63861 7243 63927 7246
rect 28625 7170 28691 7173
rect 28901 7170 28967 7173
rect 28625 7168 28967 7170
rect 28625 7112 28630 7168
rect 28686 7112 28906 7168
rect 28962 7112 28967 7168
rect 28625 7110 28967 7112
rect 28625 7107 28691 7110
rect 28901 7107 28967 7110
rect 34145 7170 34211 7173
rect 34789 7170 34855 7173
rect 34145 7168 34855 7170
rect 34145 7112 34150 7168
rect 34206 7112 34794 7168
rect 34850 7112 34855 7168
rect 34145 7110 34855 7112
rect 34145 7107 34211 7110
rect 34789 7107 34855 7110
rect 40033 7170 40099 7173
rect 49141 7170 49207 7173
rect 50153 7170 50219 7173
rect 40033 7168 50219 7170
rect 40033 7112 40038 7168
rect 40094 7112 49146 7168
rect 49202 7112 50158 7168
rect 50214 7112 50219 7168
rect 40033 7110 50219 7112
rect 40033 7107 40099 7110
rect 49141 7107 49207 7110
rect 50153 7107 50219 7110
rect 61193 7170 61259 7173
rect 65149 7170 65215 7173
rect 65333 7170 65399 7173
rect 61193 7168 65399 7170
rect 61193 7112 61198 7168
rect 61254 7112 65154 7168
rect 65210 7112 65338 7168
rect 65394 7112 65399 7168
rect 61193 7110 65399 7112
rect 61193 7107 61259 7110
rect 65149 7107 65215 7110
rect 65333 7107 65399 7110
rect 19568 7104 19888 7105
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 7039 19888 7040
rect 50288 7104 50608 7105
rect 50288 7040 50296 7104
rect 50360 7040 50376 7104
rect 50440 7040 50456 7104
rect 50520 7040 50536 7104
rect 50600 7040 50608 7104
rect 50288 7039 50608 7040
rect 81008 7104 81328 7105
rect 81008 7040 81016 7104
rect 81080 7040 81096 7104
rect 81160 7040 81176 7104
rect 81240 7040 81256 7104
rect 81320 7040 81328 7104
rect 81008 7039 81328 7040
rect 111728 7104 112048 7105
rect 111728 7040 111736 7104
rect 111800 7040 111816 7104
rect 111880 7040 111896 7104
rect 111960 7040 111976 7104
rect 112040 7040 112048 7104
rect 111728 7039 112048 7040
rect 142448 7104 142768 7105
rect 142448 7040 142456 7104
rect 142520 7040 142536 7104
rect 142600 7040 142616 7104
rect 142680 7040 142696 7104
rect 142760 7040 142768 7104
rect 142448 7039 142768 7040
rect 173168 7104 173488 7105
rect 173168 7040 173176 7104
rect 173240 7040 173256 7104
rect 173320 7040 173336 7104
rect 173400 7040 173416 7104
rect 173480 7040 173488 7104
rect 173168 7039 173488 7040
rect 31293 7034 31359 7037
rect 35893 7034 35959 7037
rect 31293 7032 35959 7034
rect 31293 6976 31298 7032
rect 31354 6976 35898 7032
rect 35954 6976 35959 7032
rect 31293 6974 35959 6976
rect 31293 6971 31359 6974
rect 35893 6971 35959 6974
rect 39941 7034 40007 7037
rect 41689 7034 41755 7037
rect 39941 7032 41755 7034
rect 39941 6976 39946 7032
rect 40002 6976 41694 7032
rect 41750 6976 41755 7032
rect 39941 6974 41755 6976
rect 39941 6971 40007 6974
rect 41689 6971 41755 6974
rect 44633 7034 44699 7037
rect 45001 7034 45067 7037
rect 47669 7034 47735 7037
rect 44633 7032 47735 7034
rect 44633 6976 44638 7032
rect 44694 6976 45006 7032
rect 45062 6976 47674 7032
rect 47730 6976 47735 7032
rect 44633 6974 47735 6976
rect 44633 6971 44699 6974
rect 45001 6971 45067 6974
rect 47669 6971 47735 6974
rect 62021 7034 62087 7037
rect 66253 7034 66319 7037
rect 62021 7032 66319 7034
rect 62021 6976 62026 7032
rect 62082 6976 66258 7032
rect 66314 6976 66319 7032
rect 62021 6974 66319 6976
rect 62021 6971 62087 6974
rect 66253 6971 66319 6974
rect 20529 6898 20595 6901
rect 23013 6898 23079 6901
rect 20529 6896 23079 6898
rect 20529 6840 20534 6896
rect 20590 6840 23018 6896
rect 23074 6840 23079 6896
rect 20529 6838 23079 6840
rect 20529 6835 20595 6838
rect 23013 6835 23079 6838
rect 33317 6898 33383 6901
rect 36077 6898 36143 6901
rect 33317 6896 36143 6898
rect 33317 6840 33322 6896
rect 33378 6840 36082 6896
rect 36138 6840 36143 6896
rect 33317 6838 36143 6840
rect 33317 6835 33383 6838
rect 36077 6835 36143 6838
rect 36629 6898 36695 6901
rect 37641 6898 37707 6901
rect 36629 6896 37707 6898
rect 36629 6840 36634 6896
rect 36690 6840 37646 6896
rect 37702 6840 37707 6896
rect 36629 6838 37707 6840
rect 36629 6835 36695 6838
rect 37641 6835 37707 6838
rect 41137 6898 41203 6901
rect 41873 6898 41939 6901
rect 41137 6896 41939 6898
rect 41137 6840 41142 6896
rect 41198 6840 41878 6896
rect 41934 6840 41939 6896
rect 41137 6838 41939 6840
rect 41137 6835 41203 6838
rect 41873 6835 41939 6838
rect 46657 6898 46723 6901
rect 47393 6898 47459 6901
rect 46657 6896 47459 6898
rect 46657 6840 46662 6896
rect 46718 6840 47398 6896
rect 47454 6840 47459 6896
rect 46657 6838 47459 6840
rect 46657 6835 46723 6838
rect 47393 6835 47459 6838
rect 64413 6898 64479 6901
rect 64781 6898 64847 6901
rect 64413 6896 64847 6898
rect 64413 6840 64418 6896
rect 64474 6840 64786 6896
rect 64842 6840 64847 6896
rect 64413 6838 64847 6840
rect 64413 6835 64479 6838
rect 64781 6835 64847 6838
rect 20989 6762 21055 6765
rect 21541 6762 21607 6765
rect 28533 6762 28599 6765
rect 20989 6760 28599 6762
rect 20989 6704 20994 6760
rect 21050 6704 21546 6760
rect 21602 6704 28538 6760
rect 28594 6704 28599 6760
rect 20989 6702 28599 6704
rect 20989 6699 21055 6702
rect 21541 6699 21607 6702
rect 28533 6699 28599 6702
rect 30281 6762 30347 6765
rect 31753 6762 31819 6765
rect 30281 6760 31819 6762
rect 30281 6704 30286 6760
rect 30342 6704 31758 6760
rect 31814 6704 31819 6760
rect 30281 6702 31819 6704
rect 30281 6699 30347 6702
rect 31753 6699 31819 6702
rect 40861 6762 40927 6765
rect 44081 6762 44147 6765
rect 47209 6762 47275 6765
rect 40861 6760 47275 6762
rect 40861 6704 40866 6760
rect 40922 6704 44086 6760
rect 44142 6704 47214 6760
rect 47270 6704 47275 6760
rect 40861 6702 47275 6704
rect 40861 6699 40927 6702
rect 44081 6699 44147 6702
rect 47209 6699 47275 6702
rect 58065 6762 58131 6765
rect 59169 6762 59235 6765
rect 62389 6762 62455 6765
rect 58065 6760 59235 6762
rect 58065 6704 58070 6760
rect 58126 6704 59174 6760
rect 59230 6704 59235 6760
rect 58065 6702 59235 6704
rect 58065 6699 58131 6702
rect 59169 6699 59235 6702
rect 59310 6760 62455 6762
rect 59310 6704 62394 6760
rect 62450 6704 62455 6760
rect 59310 6702 62455 6704
rect 46841 6626 46907 6629
rect 47853 6626 47919 6629
rect 46841 6624 47919 6626
rect 46841 6568 46846 6624
rect 46902 6568 47858 6624
rect 47914 6568 47919 6624
rect 46841 6566 47919 6568
rect 46841 6563 46907 6566
rect 47853 6563 47919 6566
rect 48957 6626 49023 6629
rect 57881 6626 57947 6629
rect 59310 6626 59370 6702
rect 62389 6699 62455 6702
rect 63309 6762 63375 6765
rect 65425 6762 65491 6765
rect 63309 6760 65491 6762
rect 63309 6704 63314 6760
rect 63370 6704 65430 6760
rect 65486 6704 65491 6760
rect 63309 6702 65491 6704
rect 63309 6699 63375 6702
rect 65425 6699 65491 6702
rect 48957 6624 57947 6626
rect 48957 6568 48962 6624
rect 49018 6568 57886 6624
rect 57942 6568 57947 6624
rect 48957 6566 57947 6568
rect 48957 6563 49023 6566
rect 57881 6563 57947 6566
rect 58206 6566 59370 6626
rect 61561 6626 61627 6629
rect 65517 6626 65583 6629
rect 61561 6624 65583 6626
rect 61561 6568 61566 6624
rect 61622 6568 65522 6624
rect 65578 6568 65583 6624
rect 61561 6566 65583 6568
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 34928 6560 35248 6561
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 6495 35248 6496
rect 46473 6490 46539 6493
rect 46933 6490 46999 6493
rect 46473 6488 46999 6490
rect 46473 6432 46478 6488
rect 46534 6432 46938 6488
rect 46994 6432 46999 6488
rect 46473 6430 46999 6432
rect 46473 6427 46539 6430
rect 46933 6427 46999 6430
rect 47485 6490 47551 6493
rect 49785 6490 49851 6493
rect 47485 6488 49851 6490
rect 47485 6432 47490 6488
rect 47546 6432 49790 6488
rect 49846 6432 49851 6488
rect 47485 6430 49851 6432
rect 47485 6427 47551 6430
rect 49785 6427 49851 6430
rect 50061 6490 50127 6493
rect 54201 6490 54267 6493
rect 50061 6488 54267 6490
rect 50061 6432 50066 6488
rect 50122 6432 54206 6488
rect 54262 6432 54267 6488
rect 50061 6430 54267 6432
rect 50061 6427 50127 6430
rect 54201 6427 54267 6430
rect 32121 6354 32187 6357
rect 58206 6354 58266 6566
rect 61561 6563 61627 6566
rect 65517 6563 65583 6566
rect 65648 6560 65968 6561
rect 65648 6496 65656 6560
rect 65720 6496 65736 6560
rect 65800 6496 65816 6560
rect 65880 6496 65896 6560
rect 65960 6496 65968 6560
rect 65648 6495 65968 6496
rect 96368 6560 96688 6561
rect 96368 6496 96376 6560
rect 96440 6496 96456 6560
rect 96520 6496 96536 6560
rect 96600 6496 96616 6560
rect 96680 6496 96688 6560
rect 96368 6495 96688 6496
rect 127088 6560 127408 6561
rect 127088 6496 127096 6560
rect 127160 6496 127176 6560
rect 127240 6496 127256 6560
rect 127320 6496 127336 6560
rect 127400 6496 127408 6560
rect 127088 6495 127408 6496
rect 157808 6560 158128 6561
rect 157808 6496 157816 6560
rect 157880 6496 157896 6560
rect 157960 6496 157976 6560
rect 158040 6496 158056 6560
rect 158120 6496 158128 6560
rect 157808 6495 158128 6496
rect 58341 6490 58407 6493
rect 63125 6490 63191 6493
rect 58341 6488 63191 6490
rect 58341 6432 58346 6488
rect 58402 6432 63130 6488
rect 63186 6432 63191 6488
rect 58341 6430 63191 6432
rect 58341 6427 58407 6430
rect 63125 6427 63191 6430
rect 32121 6352 58266 6354
rect 32121 6296 32126 6352
rect 32182 6296 58266 6352
rect 32121 6294 58266 6296
rect 58709 6354 58775 6357
rect 60641 6354 60707 6357
rect 58709 6352 60707 6354
rect 58709 6296 58714 6352
rect 58770 6296 60646 6352
rect 60702 6296 60707 6352
rect 58709 6294 60707 6296
rect 32121 6291 32187 6294
rect 58709 6291 58775 6294
rect 60641 6291 60707 6294
rect 64597 6354 64663 6357
rect 66897 6354 66963 6357
rect 64597 6352 66963 6354
rect 64597 6296 64602 6352
rect 64658 6296 66902 6352
rect 66958 6296 66963 6352
rect 64597 6294 66963 6296
rect 64597 6291 64663 6294
rect 66897 6291 66963 6294
rect 33133 6218 33199 6221
rect 36169 6218 36235 6221
rect 37181 6218 37247 6221
rect 38285 6218 38351 6221
rect 33133 6216 38351 6218
rect 33133 6160 33138 6216
rect 33194 6160 36174 6216
rect 36230 6160 37186 6216
rect 37242 6160 38290 6216
rect 38346 6160 38351 6216
rect 33133 6158 38351 6160
rect 33133 6155 33199 6158
rect 36169 6155 36235 6158
rect 37181 6155 37247 6158
rect 38285 6155 38351 6158
rect 41137 6218 41203 6221
rect 44265 6218 44331 6221
rect 41137 6216 44331 6218
rect 41137 6160 41142 6216
rect 41198 6160 44270 6216
rect 44326 6160 44331 6216
rect 41137 6158 44331 6160
rect 41137 6155 41203 6158
rect 44265 6155 44331 6158
rect 45553 6218 45619 6221
rect 47853 6218 47919 6221
rect 45553 6216 47919 6218
rect 45553 6160 45558 6216
rect 45614 6160 47858 6216
rect 47914 6160 47919 6216
rect 45553 6158 47919 6160
rect 45553 6155 45619 6158
rect 47853 6155 47919 6158
rect 48957 6218 49023 6221
rect 70393 6218 70459 6221
rect 73245 6218 73311 6221
rect 48957 6216 73311 6218
rect 48957 6160 48962 6216
rect 49018 6160 70398 6216
rect 70454 6160 73250 6216
rect 73306 6160 73311 6216
rect 48957 6158 73311 6160
rect 48957 6155 49023 6158
rect 70393 6155 70459 6158
rect 73245 6155 73311 6158
rect 31661 6082 31727 6085
rect 32857 6082 32923 6085
rect 33777 6082 33843 6085
rect 31661 6080 33843 6082
rect 31661 6024 31666 6080
rect 31722 6024 32862 6080
rect 32918 6024 33782 6080
rect 33838 6024 33843 6080
rect 31661 6022 33843 6024
rect 31661 6019 31727 6022
rect 32857 6019 32923 6022
rect 33777 6019 33843 6022
rect 46841 6082 46907 6085
rect 47577 6082 47643 6085
rect 46841 6080 47643 6082
rect 46841 6024 46846 6080
rect 46902 6024 47582 6080
rect 47638 6024 47643 6080
rect 46841 6022 47643 6024
rect 46841 6019 46907 6022
rect 47577 6019 47643 6022
rect 48681 6082 48747 6085
rect 50061 6082 50127 6085
rect 48681 6080 50127 6082
rect 48681 6024 48686 6080
rect 48742 6024 50066 6080
rect 50122 6024 50127 6080
rect 48681 6022 50127 6024
rect 48681 6019 48747 6022
rect 50061 6019 50127 6022
rect 64413 6082 64479 6085
rect 65977 6082 66043 6085
rect 64413 6080 66043 6082
rect 64413 6024 64418 6080
rect 64474 6024 65982 6080
rect 66038 6024 66043 6080
rect 64413 6022 66043 6024
rect 64413 6019 64479 6022
rect 65977 6019 66043 6022
rect 19568 6016 19888 6017
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 5951 19888 5952
rect 50288 6016 50608 6017
rect 50288 5952 50296 6016
rect 50360 5952 50376 6016
rect 50440 5952 50456 6016
rect 50520 5952 50536 6016
rect 50600 5952 50608 6016
rect 50288 5951 50608 5952
rect 81008 6016 81328 6017
rect 81008 5952 81016 6016
rect 81080 5952 81096 6016
rect 81160 5952 81176 6016
rect 81240 5952 81256 6016
rect 81320 5952 81328 6016
rect 81008 5951 81328 5952
rect 111728 6016 112048 6017
rect 111728 5952 111736 6016
rect 111800 5952 111816 6016
rect 111880 5952 111896 6016
rect 111960 5952 111976 6016
rect 112040 5952 112048 6016
rect 111728 5951 112048 5952
rect 142448 6016 142768 6017
rect 142448 5952 142456 6016
rect 142520 5952 142536 6016
rect 142600 5952 142616 6016
rect 142680 5952 142696 6016
rect 142760 5952 142768 6016
rect 142448 5951 142768 5952
rect 173168 6016 173488 6017
rect 173168 5952 173176 6016
rect 173240 5952 173256 6016
rect 173320 5952 173336 6016
rect 173400 5952 173416 6016
rect 173480 5952 173488 6016
rect 173168 5951 173488 5952
rect 46013 5946 46079 5949
rect 47485 5946 47551 5949
rect 46013 5944 47551 5946
rect 46013 5888 46018 5944
rect 46074 5888 47490 5944
rect 47546 5888 47551 5944
rect 46013 5886 47551 5888
rect 46013 5883 46079 5886
rect 47485 5883 47551 5886
rect 63125 5946 63191 5949
rect 65241 5946 65307 5949
rect 63125 5944 65307 5946
rect 63125 5888 63130 5944
rect 63186 5888 65246 5944
rect 65302 5888 65307 5944
rect 63125 5886 65307 5888
rect 63125 5883 63191 5886
rect 65241 5883 65307 5886
rect 37733 5810 37799 5813
rect 39481 5810 39547 5813
rect 37733 5808 39547 5810
rect 37733 5752 37738 5808
rect 37794 5752 39486 5808
rect 39542 5752 39547 5808
rect 37733 5750 39547 5752
rect 37733 5747 37799 5750
rect 39481 5747 39547 5750
rect 43805 5810 43871 5813
rect 48773 5810 48839 5813
rect 43805 5808 48839 5810
rect 43805 5752 43810 5808
rect 43866 5752 48778 5808
rect 48834 5752 48839 5808
rect 43805 5750 48839 5752
rect 43805 5747 43871 5750
rect 48773 5747 48839 5750
rect 53189 5810 53255 5813
rect 54293 5810 54359 5813
rect 53189 5808 54359 5810
rect 53189 5752 53194 5808
rect 53250 5752 54298 5808
rect 54354 5752 54359 5808
rect 53189 5750 54359 5752
rect 53189 5747 53255 5750
rect 54293 5747 54359 5750
rect 64229 5810 64295 5813
rect 65241 5810 65307 5813
rect 64229 5808 65307 5810
rect 64229 5752 64234 5808
rect 64290 5752 65246 5808
rect 65302 5752 65307 5808
rect 64229 5750 65307 5752
rect 64229 5747 64295 5750
rect 65241 5747 65307 5750
rect 82537 5810 82603 5813
rect 84561 5810 84627 5813
rect 82537 5808 84627 5810
rect 82537 5752 82542 5808
rect 82598 5752 84566 5808
rect 84622 5752 84627 5808
rect 82537 5750 84627 5752
rect 82537 5747 82603 5750
rect 84561 5747 84627 5750
rect 20621 5674 20687 5677
rect 21633 5674 21699 5677
rect 20621 5672 21699 5674
rect 20621 5616 20626 5672
rect 20682 5616 21638 5672
rect 21694 5616 21699 5672
rect 20621 5614 21699 5616
rect 20621 5611 20687 5614
rect 21633 5611 21699 5614
rect 31845 5674 31911 5677
rect 35249 5674 35315 5677
rect 38101 5674 38167 5677
rect 31845 5672 38167 5674
rect 31845 5616 31850 5672
rect 31906 5616 35254 5672
rect 35310 5616 38106 5672
rect 38162 5616 38167 5672
rect 31845 5614 38167 5616
rect 31845 5611 31911 5614
rect 35249 5611 35315 5614
rect 38101 5611 38167 5614
rect 46657 5674 46723 5677
rect 47485 5674 47551 5677
rect 46657 5672 47551 5674
rect 46657 5616 46662 5672
rect 46718 5616 47490 5672
rect 47546 5616 47551 5672
rect 46657 5614 47551 5616
rect 46657 5611 46723 5614
rect 47485 5611 47551 5614
rect 63401 5674 63467 5677
rect 64597 5674 64663 5677
rect 65793 5674 65859 5677
rect 63401 5672 65859 5674
rect 63401 5616 63406 5672
rect 63462 5616 64602 5672
rect 64658 5616 65798 5672
rect 65854 5616 65859 5672
rect 63401 5614 65859 5616
rect 63401 5611 63467 5614
rect 64597 5611 64663 5614
rect 65793 5611 65859 5614
rect 79041 5674 79107 5677
rect 84009 5674 84075 5677
rect 79041 5672 84075 5674
rect 79041 5616 79046 5672
rect 79102 5616 84014 5672
rect 84070 5616 84075 5672
rect 79041 5614 84075 5616
rect 79041 5611 79107 5614
rect 84009 5611 84075 5614
rect 46013 5538 46079 5541
rect 47853 5538 47919 5541
rect 46013 5536 47919 5538
rect 46013 5480 46018 5536
rect 46074 5480 47858 5536
rect 47914 5480 47919 5536
rect 46013 5478 47919 5480
rect 46013 5475 46079 5478
rect 47853 5475 47919 5478
rect 61009 5538 61075 5541
rect 65517 5538 65583 5541
rect 61009 5536 65583 5538
rect 61009 5480 61014 5536
rect 61070 5480 65522 5536
rect 65578 5480 65583 5536
rect 61009 5478 65583 5480
rect 61009 5475 61075 5478
rect 65517 5475 65583 5478
rect 83365 5538 83431 5541
rect 85757 5538 85823 5541
rect 83365 5536 85823 5538
rect 83365 5480 83370 5536
rect 83426 5480 85762 5536
rect 85818 5480 85823 5536
rect 83365 5478 85823 5480
rect 83365 5475 83431 5478
rect 85757 5475 85823 5478
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 34928 5472 35248 5473
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 5407 35248 5408
rect 65648 5472 65968 5473
rect 65648 5408 65656 5472
rect 65720 5408 65736 5472
rect 65800 5408 65816 5472
rect 65880 5408 65896 5472
rect 65960 5408 65968 5472
rect 65648 5407 65968 5408
rect 96368 5472 96688 5473
rect 96368 5408 96376 5472
rect 96440 5408 96456 5472
rect 96520 5408 96536 5472
rect 96600 5408 96616 5472
rect 96680 5408 96688 5472
rect 96368 5407 96688 5408
rect 127088 5472 127408 5473
rect 127088 5408 127096 5472
rect 127160 5408 127176 5472
rect 127240 5408 127256 5472
rect 127320 5408 127336 5472
rect 127400 5408 127408 5472
rect 127088 5407 127408 5408
rect 157808 5472 158128 5473
rect 157808 5408 157816 5472
rect 157880 5408 157896 5472
rect 157960 5408 157976 5472
rect 158040 5408 158056 5472
rect 158120 5408 158128 5472
rect 157808 5407 158128 5408
rect 78857 5402 78923 5405
rect 83733 5402 83799 5405
rect 84745 5402 84811 5405
rect 78857 5400 84811 5402
rect 78857 5344 78862 5400
rect 78918 5344 83738 5400
rect 83794 5344 84750 5400
rect 84806 5344 84811 5400
rect 78857 5342 84811 5344
rect 78857 5339 78923 5342
rect 83733 5339 83799 5342
rect 84745 5339 84811 5342
rect 43713 5266 43779 5269
rect 47393 5266 47459 5269
rect 43713 5264 47459 5266
rect 43713 5208 43718 5264
rect 43774 5208 47398 5264
rect 47454 5208 47459 5264
rect 43713 5206 47459 5208
rect 43713 5203 43779 5206
rect 47393 5203 47459 5206
rect 81801 5266 81867 5269
rect 85021 5266 85087 5269
rect 81801 5264 85087 5266
rect 81801 5208 81806 5264
rect 81862 5208 85026 5264
rect 85082 5208 85087 5264
rect 81801 5206 85087 5208
rect 81801 5203 81867 5206
rect 85021 5203 85087 5206
rect 33041 5130 33107 5133
rect 34513 5130 34579 5133
rect 80329 5130 80395 5133
rect 82261 5130 82327 5133
rect 92197 5130 92263 5133
rect 33041 5128 34579 5130
rect 33041 5072 33046 5128
rect 33102 5072 34518 5128
rect 34574 5072 34579 5128
rect 33041 5070 34579 5072
rect 33041 5067 33107 5070
rect 34513 5067 34579 5070
rect 80010 5128 81450 5130
rect 80010 5072 80334 5128
rect 80390 5072 81450 5128
rect 80010 5070 81450 5072
rect 19568 4928 19888 4929
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 4863 19888 4864
rect 50288 4928 50608 4929
rect 50288 4864 50296 4928
rect 50360 4864 50376 4928
rect 50440 4864 50456 4928
rect 50520 4864 50536 4928
rect 50600 4864 50608 4928
rect 50288 4863 50608 4864
rect 31753 4858 31819 4861
rect 37273 4858 37339 4861
rect 31753 4856 37339 4858
rect 31753 4800 31758 4856
rect 31814 4800 37278 4856
rect 37334 4800 37339 4856
rect 31753 4798 37339 4800
rect 31753 4795 31819 4798
rect 37273 4795 37339 4798
rect 69381 4722 69447 4725
rect 80010 4722 80070 5070
rect 80329 5067 80395 5070
rect 81390 4994 81450 5070
rect 82261 5128 92263 5130
rect 82261 5072 82266 5128
rect 82322 5072 92202 5128
rect 92258 5072 92263 5128
rect 82261 5070 92263 5072
rect 82261 5067 82327 5070
rect 92197 5067 92263 5070
rect 84837 4994 84903 4997
rect 81390 4992 84903 4994
rect 81390 4936 84842 4992
rect 84898 4936 84903 4992
rect 81390 4934 84903 4936
rect 84837 4931 84903 4934
rect 81008 4928 81328 4929
rect 81008 4864 81016 4928
rect 81080 4864 81096 4928
rect 81160 4864 81176 4928
rect 81240 4864 81256 4928
rect 81320 4864 81328 4928
rect 81008 4863 81328 4864
rect 111728 4928 112048 4929
rect 111728 4864 111736 4928
rect 111800 4864 111816 4928
rect 111880 4864 111896 4928
rect 111960 4864 111976 4928
rect 112040 4864 112048 4928
rect 111728 4863 112048 4864
rect 142448 4928 142768 4929
rect 142448 4864 142456 4928
rect 142520 4864 142536 4928
rect 142600 4864 142616 4928
rect 142680 4864 142696 4928
rect 142760 4864 142768 4928
rect 142448 4863 142768 4864
rect 173168 4928 173488 4929
rect 173168 4864 173176 4928
rect 173240 4864 173256 4928
rect 173320 4864 173336 4928
rect 173400 4864 173416 4928
rect 173480 4864 173488 4928
rect 173168 4863 173488 4864
rect 81709 4858 81775 4861
rect 87873 4858 87939 4861
rect 88517 4858 88583 4861
rect 89621 4858 89687 4861
rect 81709 4856 89687 4858
rect 81709 4800 81714 4856
rect 81770 4800 87878 4856
rect 87934 4800 88522 4856
rect 88578 4800 89626 4856
rect 89682 4800 89687 4856
rect 81709 4798 89687 4800
rect 81709 4795 81775 4798
rect 87873 4795 87939 4798
rect 88517 4795 88583 4798
rect 89621 4795 89687 4798
rect 69381 4720 80070 4722
rect 69381 4664 69386 4720
rect 69442 4664 80070 4720
rect 69381 4662 80070 4664
rect 69381 4659 69447 4662
rect 80646 4660 80652 4724
rect 80716 4722 80722 4724
rect 86493 4722 86559 4725
rect 80716 4720 86559 4722
rect 80716 4664 86498 4720
rect 86554 4664 86559 4720
rect 80716 4662 86559 4664
rect 80716 4660 80722 4662
rect 86493 4659 86559 4662
rect 75269 4586 75335 4589
rect 88425 4586 88491 4589
rect 75269 4584 88491 4586
rect 75269 4528 75274 4584
rect 75330 4528 88430 4584
rect 88486 4528 88491 4584
rect 75269 4526 88491 4528
rect 75269 4523 75335 4526
rect 88425 4523 88491 4526
rect 31661 4450 31727 4453
rect 31845 4450 31911 4453
rect 31661 4448 31911 4450
rect 31661 4392 31666 4448
rect 31722 4392 31850 4448
rect 31906 4392 31911 4448
rect 31661 4390 31911 4392
rect 31661 4387 31727 4390
rect 31845 4387 31911 4390
rect 78397 4450 78463 4453
rect 82997 4450 83063 4453
rect 78397 4448 83063 4450
rect 78397 4392 78402 4448
rect 78458 4392 83002 4448
rect 83058 4392 83063 4448
rect 78397 4390 83063 4392
rect 78397 4387 78463 4390
rect 82997 4387 83063 4390
rect 83917 4450 83983 4453
rect 85849 4450 85915 4453
rect 83917 4448 85915 4450
rect 83917 4392 83922 4448
rect 83978 4392 85854 4448
rect 85910 4392 85915 4448
rect 83917 4390 85915 4392
rect 83917 4387 83983 4390
rect 85849 4387 85915 4390
rect 87597 4450 87663 4453
rect 89713 4450 89779 4453
rect 87597 4448 89779 4450
rect 87597 4392 87602 4448
rect 87658 4392 89718 4448
rect 89774 4392 89779 4448
rect 87597 4390 89779 4392
rect 87597 4387 87663 4390
rect 89713 4387 89779 4390
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 34928 4384 35248 4385
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 4319 35248 4320
rect 65648 4384 65968 4385
rect 65648 4320 65656 4384
rect 65720 4320 65736 4384
rect 65800 4320 65816 4384
rect 65880 4320 65896 4384
rect 65960 4320 65968 4384
rect 65648 4319 65968 4320
rect 96368 4384 96688 4385
rect 96368 4320 96376 4384
rect 96440 4320 96456 4384
rect 96520 4320 96536 4384
rect 96600 4320 96616 4384
rect 96680 4320 96688 4384
rect 96368 4319 96688 4320
rect 127088 4384 127408 4385
rect 127088 4320 127096 4384
rect 127160 4320 127176 4384
rect 127240 4320 127256 4384
rect 127320 4320 127336 4384
rect 127400 4320 127408 4384
rect 127088 4319 127408 4320
rect 157808 4384 158128 4385
rect 157808 4320 157816 4384
rect 157880 4320 157896 4384
rect 157960 4320 157976 4384
rect 158040 4320 158056 4384
rect 158120 4320 158128 4384
rect 157808 4319 158128 4320
rect 79685 4314 79751 4317
rect 80421 4314 80487 4317
rect 79685 4312 80487 4314
rect 79685 4256 79690 4312
rect 79746 4256 80426 4312
rect 80482 4256 80487 4312
rect 79685 4254 80487 4256
rect 79685 4251 79751 4254
rect 80421 4251 80487 4254
rect 84193 4314 84259 4317
rect 84837 4314 84903 4317
rect 84193 4312 84903 4314
rect 84193 4256 84198 4312
rect 84254 4256 84842 4312
rect 84898 4256 84903 4312
rect 84193 4254 84903 4256
rect 84193 4251 84259 4254
rect 84837 4251 84903 4254
rect 86534 4252 86540 4316
rect 86604 4314 86610 4316
rect 86769 4314 86835 4317
rect 86604 4312 86835 4314
rect 86604 4256 86774 4312
rect 86830 4256 86835 4312
rect 86604 4254 86835 4256
rect 86604 4252 86610 4254
rect 86769 4251 86835 4254
rect 87965 4314 88031 4317
rect 95049 4314 95115 4317
rect 87965 4312 95115 4314
rect 87965 4256 87970 4312
rect 88026 4256 95054 4312
rect 95110 4256 95115 4312
rect 87965 4254 95115 4256
rect 87965 4251 88031 4254
rect 95049 4251 95115 4254
rect 36077 4178 36143 4181
rect 39849 4178 39915 4181
rect 36077 4176 39915 4178
rect 36077 4120 36082 4176
rect 36138 4120 39854 4176
rect 39910 4120 39915 4176
rect 36077 4118 39915 4120
rect 36077 4115 36143 4118
rect 39849 4115 39915 4118
rect 79409 4178 79475 4181
rect 91001 4178 91067 4181
rect 79409 4176 91067 4178
rect 79409 4120 79414 4176
rect 79470 4120 91006 4176
rect 91062 4120 91067 4176
rect 79409 4118 91067 4120
rect 79409 4115 79475 4118
rect 91001 4115 91067 4118
rect 12433 4042 12499 4045
rect 21633 4042 21699 4045
rect 12433 4040 21699 4042
rect 12433 3984 12438 4040
rect 12494 3984 21638 4040
rect 21694 3984 21699 4040
rect 12433 3982 21699 3984
rect 12433 3979 12499 3982
rect 21633 3979 21699 3982
rect 22093 4042 22159 4045
rect 30557 4042 30623 4045
rect 22093 4040 30623 4042
rect 22093 3984 22098 4040
rect 22154 3984 30562 4040
rect 30618 3984 30623 4040
rect 22093 3982 30623 3984
rect 22093 3979 22159 3982
rect 30557 3979 30623 3982
rect 73245 4042 73311 4045
rect 86217 4042 86283 4045
rect 86769 4044 86835 4045
rect 86718 4042 86724 4044
rect 73245 4040 86283 4042
rect 73245 3984 73250 4040
rect 73306 3984 86222 4040
rect 86278 3984 86283 4040
rect 73245 3982 86283 3984
rect 86678 3982 86724 4042
rect 86788 4040 86835 4044
rect 86830 3984 86835 4040
rect 73245 3979 73311 3982
rect 86217 3979 86283 3982
rect 86718 3980 86724 3982
rect 86788 3980 86835 3984
rect 86769 3979 86835 3980
rect 88609 4042 88675 4045
rect 101581 4042 101647 4045
rect 88609 4040 101647 4042
rect 88609 3984 88614 4040
rect 88670 3984 101586 4040
rect 101642 3984 101647 4040
rect 88609 3982 101647 3984
rect 88609 3979 88675 3982
rect 101581 3979 101647 3982
rect 71497 3906 71563 3909
rect 77845 3906 77911 3909
rect 71497 3904 77911 3906
rect 71497 3848 71502 3904
rect 71558 3848 77850 3904
rect 77906 3848 77911 3904
rect 71497 3846 77911 3848
rect 71497 3843 71563 3846
rect 77845 3843 77911 3846
rect 82813 3906 82879 3909
rect 85389 3906 85455 3909
rect 82813 3904 85455 3906
rect 82813 3848 82818 3904
rect 82874 3848 85394 3904
rect 85450 3848 85455 3904
rect 82813 3846 85455 3848
rect 82813 3843 82879 3846
rect 85389 3843 85455 3846
rect 86217 3906 86283 3909
rect 97993 3906 98059 3909
rect 86217 3904 98059 3906
rect 86217 3848 86222 3904
rect 86278 3848 97998 3904
rect 98054 3848 98059 3904
rect 86217 3846 98059 3848
rect 86217 3843 86283 3846
rect 97993 3843 98059 3846
rect 19568 3840 19888 3841
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 3775 19888 3776
rect 50288 3840 50608 3841
rect 50288 3776 50296 3840
rect 50360 3776 50376 3840
rect 50440 3776 50456 3840
rect 50520 3776 50536 3840
rect 50600 3776 50608 3840
rect 50288 3775 50608 3776
rect 81008 3840 81328 3841
rect 81008 3776 81016 3840
rect 81080 3776 81096 3840
rect 81160 3776 81176 3840
rect 81240 3776 81256 3840
rect 81320 3776 81328 3840
rect 81008 3775 81328 3776
rect 111728 3840 112048 3841
rect 111728 3776 111736 3840
rect 111800 3776 111816 3840
rect 111880 3776 111896 3840
rect 111960 3776 111976 3840
rect 112040 3776 112048 3840
rect 111728 3775 112048 3776
rect 142448 3840 142768 3841
rect 142448 3776 142456 3840
rect 142520 3776 142536 3840
rect 142600 3776 142616 3840
rect 142680 3776 142696 3840
rect 142760 3776 142768 3840
rect 142448 3775 142768 3776
rect 173168 3840 173488 3841
rect 173168 3776 173176 3840
rect 173240 3776 173256 3840
rect 173320 3776 173336 3840
rect 173400 3776 173416 3840
rect 173480 3776 173488 3840
rect 173168 3775 173488 3776
rect 11881 3770 11947 3773
rect 12617 3770 12683 3773
rect 11881 3768 12683 3770
rect 11881 3712 11886 3768
rect 11942 3712 12622 3768
rect 12678 3712 12683 3768
rect 11881 3710 12683 3712
rect 11881 3707 11947 3710
rect 12617 3707 12683 3710
rect 68277 3770 68343 3773
rect 79685 3770 79751 3773
rect 68277 3768 79751 3770
rect 68277 3712 68282 3768
rect 68338 3712 79690 3768
rect 79746 3712 79751 3768
rect 68277 3710 79751 3712
rect 68277 3707 68343 3710
rect 79685 3707 79751 3710
rect 84101 3770 84167 3773
rect 85481 3770 85547 3773
rect 88374 3770 88380 3772
rect 84101 3768 88380 3770
rect 84101 3712 84106 3768
rect 84162 3712 85486 3768
rect 85542 3712 88380 3768
rect 84101 3710 88380 3712
rect 84101 3707 84167 3710
rect 85481 3707 85547 3710
rect 88374 3708 88380 3710
rect 88444 3708 88450 3772
rect 88701 3770 88767 3773
rect 101857 3770 101923 3773
rect 88701 3768 101923 3770
rect 88701 3712 88706 3768
rect 88762 3712 101862 3768
rect 101918 3712 101923 3768
rect 88701 3710 101923 3712
rect 88701 3707 88767 3710
rect 101857 3707 101923 3710
rect 20897 3634 20963 3637
rect 28901 3634 28967 3637
rect 20897 3632 28967 3634
rect 20897 3576 20902 3632
rect 20958 3576 28906 3632
rect 28962 3576 28967 3632
rect 20897 3574 28967 3576
rect 20897 3571 20963 3574
rect 28901 3571 28967 3574
rect 72141 3634 72207 3637
rect 75821 3634 75887 3637
rect 72141 3632 75887 3634
rect 72141 3576 72146 3632
rect 72202 3576 75826 3632
rect 75882 3576 75887 3632
rect 72141 3574 75887 3576
rect 72141 3571 72207 3574
rect 75821 3571 75887 3574
rect 76281 3634 76347 3637
rect 88609 3634 88675 3637
rect 76281 3632 88675 3634
rect 76281 3576 76286 3632
rect 76342 3576 88614 3632
rect 88670 3576 88675 3632
rect 76281 3574 88675 3576
rect 76281 3571 76347 3574
rect 88609 3571 88675 3574
rect 88742 3572 88748 3636
rect 88812 3634 88818 3636
rect 89662 3634 89668 3636
rect 88812 3574 89668 3634
rect 88812 3572 88818 3574
rect 89662 3572 89668 3574
rect 89732 3572 89738 3636
rect 89846 3572 89852 3636
rect 89916 3634 89922 3636
rect 95601 3634 95667 3637
rect 101765 3634 101831 3637
rect 89916 3632 95667 3634
rect 89916 3576 95606 3632
rect 95662 3576 95667 3632
rect 89916 3574 95667 3576
rect 89916 3572 89922 3574
rect 95601 3571 95667 3574
rect 96570 3632 101831 3634
rect 96570 3576 101770 3632
rect 101826 3576 101831 3632
rect 96570 3574 101831 3576
rect 10133 3498 10199 3501
rect 15653 3498 15719 3501
rect 10133 3496 15719 3498
rect 10133 3440 10138 3496
rect 10194 3440 15658 3496
rect 15714 3440 15719 3496
rect 10133 3438 15719 3440
rect 10133 3435 10199 3438
rect 15653 3435 15719 3438
rect 21265 3498 21331 3501
rect 22277 3498 22343 3501
rect 21265 3496 22343 3498
rect 21265 3440 21270 3496
rect 21326 3440 22282 3496
rect 22338 3440 22343 3496
rect 21265 3438 22343 3440
rect 21265 3435 21331 3438
rect 22277 3435 22343 3438
rect 69749 3498 69815 3501
rect 75085 3498 75151 3501
rect 69749 3496 75151 3498
rect 69749 3440 69754 3496
rect 69810 3440 75090 3496
rect 75146 3440 75151 3496
rect 69749 3438 75151 3440
rect 69749 3435 69815 3438
rect 75085 3435 75151 3438
rect 75821 3498 75887 3501
rect 79869 3498 79935 3501
rect 80605 3498 80671 3501
rect 75821 3496 80671 3498
rect 75821 3440 75826 3496
rect 75882 3440 79874 3496
rect 79930 3440 80610 3496
rect 80666 3440 80671 3496
rect 75821 3438 80671 3440
rect 75821 3435 75887 3438
rect 79869 3435 79935 3438
rect 80605 3435 80671 3438
rect 81065 3498 81131 3501
rect 85665 3498 85731 3501
rect 81065 3496 85731 3498
rect 81065 3440 81070 3496
rect 81126 3440 85670 3496
rect 85726 3440 85731 3496
rect 81065 3438 85731 3440
rect 81065 3435 81131 3438
rect 85665 3435 85731 3438
rect 86166 3436 86172 3500
rect 86236 3498 86242 3500
rect 88425 3498 88491 3501
rect 96570 3498 96630 3574
rect 101765 3571 101831 3574
rect 86236 3438 88258 3498
rect 86236 3436 86242 3438
rect 68553 3362 68619 3365
rect 77385 3362 77451 3365
rect 77753 3362 77819 3365
rect 68553 3360 77819 3362
rect 68553 3304 68558 3360
rect 68614 3304 77390 3360
rect 77446 3304 77758 3360
rect 77814 3304 77819 3360
rect 68553 3302 77819 3304
rect 68553 3299 68619 3302
rect 77385 3299 77451 3302
rect 77753 3299 77819 3302
rect 79041 3362 79107 3365
rect 87965 3362 88031 3365
rect 79041 3360 88031 3362
rect 79041 3304 79046 3360
rect 79102 3304 87970 3360
rect 88026 3304 88031 3360
rect 79041 3302 88031 3304
rect 88198 3362 88258 3438
rect 88425 3496 96630 3498
rect 88425 3440 88430 3496
rect 88486 3440 96630 3496
rect 88425 3438 96630 3440
rect 88425 3435 88491 3438
rect 93209 3362 93275 3365
rect 88198 3360 93275 3362
rect 88198 3304 93214 3360
rect 93270 3304 93275 3360
rect 88198 3302 93275 3304
rect 79041 3299 79107 3302
rect 87965 3299 88031 3302
rect 93209 3299 93275 3302
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 34928 3296 35248 3297
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 3231 35248 3232
rect 65648 3296 65968 3297
rect 65648 3232 65656 3296
rect 65720 3232 65736 3296
rect 65800 3232 65816 3296
rect 65880 3232 65896 3296
rect 65960 3232 65968 3296
rect 65648 3231 65968 3232
rect 96368 3296 96688 3297
rect 96368 3232 96376 3296
rect 96440 3232 96456 3296
rect 96520 3232 96536 3296
rect 96600 3232 96616 3296
rect 96680 3232 96688 3296
rect 96368 3231 96688 3232
rect 127088 3296 127408 3297
rect 127088 3232 127096 3296
rect 127160 3232 127176 3296
rect 127240 3232 127256 3296
rect 127320 3232 127336 3296
rect 127400 3232 127408 3296
rect 127088 3231 127408 3232
rect 157808 3296 158128 3297
rect 157808 3232 157816 3296
rect 157880 3232 157896 3296
rect 157960 3232 157976 3296
rect 158040 3232 158056 3296
rect 158120 3232 158128 3296
rect 157808 3231 158128 3232
rect 17677 3226 17743 3229
rect 19057 3226 19123 3229
rect 17677 3224 19123 3226
rect 17677 3168 17682 3224
rect 17738 3168 19062 3224
rect 19118 3168 19123 3224
rect 17677 3166 19123 3168
rect 17677 3163 17743 3166
rect 19057 3163 19123 3166
rect 21081 3226 21147 3229
rect 28165 3226 28231 3229
rect 21081 3224 28231 3226
rect 21081 3168 21086 3224
rect 21142 3168 28170 3224
rect 28226 3168 28231 3224
rect 21081 3166 28231 3168
rect 21081 3163 21147 3166
rect 28165 3163 28231 3166
rect 70669 3226 70735 3229
rect 78581 3226 78647 3229
rect 70669 3224 78647 3226
rect 70669 3168 70674 3224
rect 70730 3168 78586 3224
rect 78642 3168 78647 3224
rect 70669 3166 78647 3168
rect 70669 3163 70735 3166
rect 78581 3163 78647 3166
rect 78765 3226 78831 3229
rect 90817 3226 90883 3229
rect 103513 3226 103579 3229
rect 78765 3224 90883 3226
rect 78765 3168 78770 3224
rect 78826 3168 90822 3224
rect 90878 3168 90883 3224
rect 78765 3166 90883 3168
rect 78765 3163 78831 3166
rect 90817 3163 90883 3166
rect 99330 3224 103579 3226
rect 99330 3168 103518 3224
rect 103574 3168 103579 3224
rect 99330 3166 103579 3168
rect 1669 3090 1735 3093
rect 2630 3090 2636 3092
rect 1669 3088 2636 3090
rect 1669 3032 1674 3088
rect 1730 3032 2636 3088
rect 1669 3030 2636 3032
rect 1669 3027 1735 3030
rect 2630 3028 2636 3030
rect 2700 3028 2706 3092
rect 11973 3090 12039 3093
rect 12525 3090 12591 3093
rect 11973 3088 12591 3090
rect 11973 3032 11978 3088
rect 12034 3032 12530 3088
rect 12586 3032 12591 3088
rect 11973 3030 12591 3032
rect 11973 3027 12039 3030
rect 12525 3027 12591 3030
rect 22369 3090 22435 3093
rect 28165 3090 28231 3093
rect 22369 3088 28231 3090
rect 22369 3032 22374 3088
rect 22430 3032 28170 3088
rect 28226 3032 28231 3088
rect 22369 3030 28231 3032
rect 22369 3027 22435 3030
rect 28165 3027 28231 3030
rect 70025 3090 70091 3093
rect 71957 3090 72023 3093
rect 70025 3088 72023 3090
rect 70025 3032 70030 3088
rect 70086 3032 71962 3088
rect 72018 3032 72023 3088
rect 70025 3030 72023 3032
rect 70025 3027 70091 3030
rect 71957 3027 72023 3030
rect 73429 3090 73495 3093
rect 75545 3090 75611 3093
rect 73429 3088 75611 3090
rect 73429 3032 73434 3088
rect 73490 3032 75550 3088
rect 75606 3032 75611 3088
rect 73429 3030 75611 3032
rect 73429 3027 73495 3030
rect 75545 3027 75611 3030
rect 76649 3090 76715 3093
rect 85757 3090 85823 3093
rect 86493 3090 86559 3093
rect 76649 3088 84946 3090
rect 76649 3032 76654 3088
rect 76710 3032 84946 3088
rect 76649 3030 84946 3032
rect 76649 3027 76715 3030
rect 15193 2954 15259 2957
rect 17493 2954 17559 2957
rect 15193 2952 17559 2954
rect 15193 2896 15198 2952
rect 15254 2896 17498 2952
rect 17554 2896 17559 2952
rect 15193 2894 17559 2896
rect 15193 2891 15259 2894
rect 17493 2891 17559 2894
rect 68645 2954 68711 2957
rect 70485 2954 70551 2957
rect 68645 2952 70551 2954
rect 68645 2896 68650 2952
rect 68706 2896 70490 2952
rect 70546 2896 70551 2952
rect 68645 2894 70551 2896
rect 68645 2891 68711 2894
rect 70485 2891 70551 2894
rect 71313 2954 71379 2957
rect 74625 2954 74691 2957
rect 71313 2952 74691 2954
rect 71313 2896 71318 2952
rect 71374 2896 74630 2952
rect 74686 2896 74691 2952
rect 71313 2894 74691 2896
rect 71313 2891 71379 2894
rect 74625 2891 74691 2894
rect 79041 2954 79107 2957
rect 84886 2954 84946 3030
rect 85757 3088 86559 3090
rect 85757 3032 85762 3088
rect 85818 3032 86498 3088
rect 86554 3032 86559 3088
rect 85757 3030 86559 3032
rect 85757 3027 85823 3030
rect 86493 3027 86559 3030
rect 86953 3090 87019 3093
rect 87229 3090 87295 3093
rect 86953 3088 87295 3090
rect 86953 3032 86958 3088
rect 87014 3032 87234 3088
rect 87290 3032 87295 3088
rect 86953 3030 87295 3032
rect 86953 3027 87019 3030
rect 87229 3027 87295 3030
rect 88057 3090 88123 3093
rect 99330 3090 99390 3166
rect 103513 3163 103579 3166
rect 88057 3088 99390 3090
rect 88057 3032 88062 3088
rect 88118 3032 99390 3088
rect 88057 3030 99390 3032
rect 102133 3092 102199 3093
rect 102133 3088 102180 3092
rect 102244 3090 102250 3092
rect 102133 3032 102138 3088
rect 88057 3027 88123 3030
rect 102133 3028 102180 3032
rect 102244 3030 102290 3090
rect 102244 3028 102250 3030
rect 102133 3027 102199 3028
rect 89161 2954 89227 2957
rect 79041 2952 84762 2954
rect 79041 2896 79046 2952
rect 79102 2896 84762 2952
rect 79041 2894 84762 2896
rect 84886 2952 89227 2954
rect 84886 2896 89166 2952
rect 89222 2896 89227 2952
rect 84886 2894 89227 2896
rect 79041 2891 79107 2894
rect 17677 2818 17743 2821
rect 18505 2818 18571 2821
rect 17677 2816 18571 2818
rect 17677 2760 17682 2816
rect 17738 2760 18510 2816
rect 18566 2760 18571 2816
rect 17677 2758 18571 2760
rect 17677 2755 17743 2758
rect 18505 2755 18571 2758
rect 75637 2818 75703 2821
rect 79685 2818 79751 2821
rect 75637 2816 79751 2818
rect 75637 2760 75642 2816
rect 75698 2760 79690 2816
rect 79746 2760 79751 2816
rect 75637 2758 79751 2760
rect 75637 2755 75703 2758
rect 79685 2755 79751 2758
rect 80646 2756 80652 2820
rect 80716 2818 80722 2820
rect 80881 2818 80947 2821
rect 80716 2816 80947 2818
rect 80716 2760 80886 2816
rect 80942 2760 80947 2816
rect 80716 2758 80947 2760
rect 80716 2756 80722 2758
rect 19568 2752 19888 2753
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2687 19888 2688
rect 50288 2752 50608 2753
rect 50288 2688 50296 2752
rect 50360 2688 50376 2752
rect 50440 2688 50456 2752
rect 50520 2688 50536 2752
rect 50600 2688 50608 2752
rect 50288 2687 50608 2688
rect 78857 2682 78923 2685
rect 80654 2682 80714 2756
rect 80881 2755 80947 2758
rect 83733 2818 83799 2821
rect 84193 2818 84259 2821
rect 83733 2816 84259 2818
rect 83733 2760 83738 2816
rect 83794 2760 84198 2816
rect 84254 2760 84259 2816
rect 83733 2758 84259 2760
rect 84702 2818 84762 2894
rect 89161 2891 89227 2894
rect 101397 2954 101463 2957
rect 102869 2954 102935 2957
rect 101397 2952 102935 2954
rect 101397 2896 101402 2952
rect 101458 2896 102874 2952
rect 102930 2896 102935 2952
rect 101397 2894 102935 2896
rect 101397 2891 101463 2894
rect 102869 2891 102935 2894
rect 86166 2818 86172 2820
rect 84702 2758 86172 2818
rect 83733 2755 83799 2758
rect 84193 2755 84259 2758
rect 86166 2756 86172 2758
rect 86236 2756 86242 2820
rect 86401 2818 86467 2821
rect 86534 2818 86540 2820
rect 86401 2816 86540 2818
rect 86401 2760 86406 2816
rect 86462 2760 86540 2816
rect 86401 2758 86540 2760
rect 86401 2755 86467 2758
rect 86534 2756 86540 2758
rect 86604 2756 86610 2820
rect 86769 2818 86835 2821
rect 87321 2818 87387 2821
rect 86769 2816 87387 2818
rect 86769 2760 86774 2816
rect 86830 2760 87326 2816
rect 87382 2760 87387 2816
rect 86769 2758 87387 2760
rect 86769 2755 86835 2758
rect 87321 2755 87387 2758
rect 89621 2818 89687 2821
rect 101029 2818 101095 2821
rect 89621 2816 101095 2818
rect 89621 2760 89626 2816
rect 89682 2760 101034 2816
rect 101090 2760 101095 2816
rect 89621 2758 101095 2760
rect 89621 2755 89687 2758
rect 101029 2755 101095 2758
rect 81008 2752 81328 2753
rect 81008 2688 81016 2752
rect 81080 2688 81096 2752
rect 81160 2688 81176 2752
rect 81240 2688 81256 2752
rect 81320 2688 81328 2752
rect 81008 2687 81328 2688
rect 111728 2752 112048 2753
rect 111728 2688 111736 2752
rect 111800 2688 111816 2752
rect 111880 2688 111896 2752
rect 111960 2688 111976 2752
rect 112040 2688 112048 2752
rect 111728 2687 112048 2688
rect 142448 2752 142768 2753
rect 142448 2688 142456 2752
rect 142520 2688 142536 2752
rect 142600 2688 142616 2752
rect 142680 2688 142696 2752
rect 142760 2688 142768 2752
rect 142448 2687 142768 2688
rect 173168 2752 173488 2753
rect 173168 2688 173176 2752
rect 173240 2688 173256 2752
rect 173320 2688 173336 2752
rect 173400 2688 173416 2752
rect 173480 2688 173488 2752
rect 173168 2687 173488 2688
rect 78857 2680 80714 2682
rect 78857 2624 78862 2680
rect 78918 2624 80714 2680
rect 78857 2622 80714 2624
rect 81709 2682 81775 2685
rect 95141 2682 95207 2685
rect 81709 2680 95207 2682
rect 81709 2624 81714 2680
rect 81770 2624 95146 2680
rect 95202 2624 95207 2680
rect 81709 2622 95207 2624
rect 78857 2619 78923 2622
rect 81709 2619 81775 2622
rect 95141 2619 95207 2622
rect 1669 2546 1735 2549
rect 94681 2546 94747 2549
rect 1669 2544 94747 2546
rect 1669 2488 1674 2544
rect 1730 2488 94686 2544
rect 94742 2488 94747 2544
rect 1669 2486 94747 2488
rect 1669 2483 1735 2486
rect 94681 2483 94747 2486
rect 74901 2410 74967 2413
rect 83181 2410 83247 2413
rect 74901 2408 83247 2410
rect 74901 2352 74906 2408
rect 74962 2352 83186 2408
rect 83242 2352 83247 2408
rect 74901 2350 83247 2352
rect 74901 2347 74967 2350
rect 83181 2347 83247 2350
rect 84561 2410 84627 2413
rect 86677 2410 86743 2413
rect 84561 2408 86743 2410
rect 84561 2352 84566 2408
rect 84622 2352 86682 2408
rect 86738 2352 86743 2408
rect 84561 2350 86743 2352
rect 84561 2347 84627 2350
rect 86677 2347 86743 2350
rect 78949 2274 79015 2277
rect 87689 2274 87755 2277
rect 93577 2274 93643 2277
rect 78949 2272 85590 2274
rect 78949 2216 78954 2272
rect 79010 2216 85590 2272
rect 78949 2214 85590 2216
rect 78949 2211 79015 2214
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 34928 2208 35248 2209
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2143 35248 2144
rect 65648 2208 65968 2209
rect 65648 2144 65656 2208
rect 65720 2144 65736 2208
rect 65800 2144 65816 2208
rect 65880 2144 65896 2208
rect 65960 2144 65968 2208
rect 65648 2143 65968 2144
rect 80421 2138 80487 2141
rect 85205 2138 85271 2141
rect 80421 2136 85271 2138
rect 80421 2080 80426 2136
rect 80482 2080 85210 2136
rect 85266 2080 85271 2136
rect 80421 2078 85271 2080
rect 85530 2138 85590 2214
rect 87689 2272 93643 2274
rect 87689 2216 87694 2272
rect 87750 2216 93582 2272
rect 93638 2216 93643 2272
rect 87689 2214 93643 2216
rect 87689 2211 87755 2214
rect 93577 2211 93643 2214
rect 96368 2208 96688 2209
rect 96368 2144 96376 2208
rect 96440 2144 96456 2208
rect 96520 2144 96536 2208
rect 96600 2144 96616 2208
rect 96680 2144 96688 2208
rect 96368 2143 96688 2144
rect 127088 2208 127408 2209
rect 127088 2144 127096 2208
rect 127160 2144 127176 2208
rect 127240 2144 127256 2208
rect 127320 2144 127336 2208
rect 127400 2144 127408 2208
rect 127088 2143 127408 2144
rect 157808 2208 158128 2209
rect 157808 2144 157816 2208
rect 157880 2144 157896 2208
rect 157960 2144 157976 2208
rect 158040 2144 158056 2208
rect 158120 2144 158128 2208
rect 157808 2143 158128 2144
rect 86493 2138 86559 2141
rect 91829 2138 91895 2141
rect 85530 2136 91895 2138
rect 85530 2080 86498 2136
rect 86554 2080 91834 2136
rect 91890 2080 91895 2136
rect 85530 2078 91895 2080
rect 80421 2075 80487 2078
rect 85205 2075 85271 2078
rect 86493 2075 86559 2078
rect 91829 2075 91895 2078
rect 86769 2004 86835 2005
rect 86718 1940 86724 2004
rect 86788 2002 86835 2004
rect 86788 2000 86880 2002
rect 86830 1944 86880 2000
rect 86788 1942 86880 1944
rect 86788 1940 86835 1942
rect 86769 1939 86835 1940
<< via3 >>
rect 4216 117532 4280 117536
rect 4216 117476 4220 117532
rect 4220 117476 4276 117532
rect 4276 117476 4280 117532
rect 4216 117472 4280 117476
rect 4296 117532 4360 117536
rect 4296 117476 4300 117532
rect 4300 117476 4356 117532
rect 4356 117476 4360 117532
rect 4296 117472 4360 117476
rect 4376 117532 4440 117536
rect 4376 117476 4380 117532
rect 4380 117476 4436 117532
rect 4436 117476 4440 117532
rect 4376 117472 4440 117476
rect 4456 117532 4520 117536
rect 4456 117476 4460 117532
rect 4460 117476 4516 117532
rect 4516 117476 4520 117532
rect 4456 117472 4520 117476
rect 34936 117532 35000 117536
rect 34936 117476 34940 117532
rect 34940 117476 34996 117532
rect 34996 117476 35000 117532
rect 34936 117472 35000 117476
rect 35016 117532 35080 117536
rect 35016 117476 35020 117532
rect 35020 117476 35076 117532
rect 35076 117476 35080 117532
rect 35016 117472 35080 117476
rect 35096 117532 35160 117536
rect 35096 117476 35100 117532
rect 35100 117476 35156 117532
rect 35156 117476 35160 117532
rect 35096 117472 35160 117476
rect 35176 117532 35240 117536
rect 35176 117476 35180 117532
rect 35180 117476 35236 117532
rect 35236 117476 35240 117532
rect 35176 117472 35240 117476
rect 65656 117532 65720 117536
rect 65656 117476 65660 117532
rect 65660 117476 65716 117532
rect 65716 117476 65720 117532
rect 65656 117472 65720 117476
rect 65736 117532 65800 117536
rect 65736 117476 65740 117532
rect 65740 117476 65796 117532
rect 65796 117476 65800 117532
rect 65736 117472 65800 117476
rect 65816 117532 65880 117536
rect 65816 117476 65820 117532
rect 65820 117476 65876 117532
rect 65876 117476 65880 117532
rect 65816 117472 65880 117476
rect 65896 117532 65960 117536
rect 65896 117476 65900 117532
rect 65900 117476 65956 117532
rect 65956 117476 65960 117532
rect 65896 117472 65960 117476
rect 96376 117532 96440 117536
rect 96376 117476 96380 117532
rect 96380 117476 96436 117532
rect 96436 117476 96440 117532
rect 96376 117472 96440 117476
rect 96456 117532 96520 117536
rect 96456 117476 96460 117532
rect 96460 117476 96516 117532
rect 96516 117476 96520 117532
rect 96456 117472 96520 117476
rect 96536 117532 96600 117536
rect 96536 117476 96540 117532
rect 96540 117476 96596 117532
rect 96596 117476 96600 117532
rect 96536 117472 96600 117476
rect 96616 117532 96680 117536
rect 96616 117476 96620 117532
rect 96620 117476 96676 117532
rect 96676 117476 96680 117532
rect 96616 117472 96680 117476
rect 127096 117532 127160 117536
rect 127096 117476 127100 117532
rect 127100 117476 127156 117532
rect 127156 117476 127160 117532
rect 127096 117472 127160 117476
rect 127176 117532 127240 117536
rect 127176 117476 127180 117532
rect 127180 117476 127236 117532
rect 127236 117476 127240 117532
rect 127176 117472 127240 117476
rect 127256 117532 127320 117536
rect 127256 117476 127260 117532
rect 127260 117476 127316 117532
rect 127316 117476 127320 117532
rect 127256 117472 127320 117476
rect 127336 117532 127400 117536
rect 127336 117476 127340 117532
rect 127340 117476 127396 117532
rect 127396 117476 127400 117532
rect 127336 117472 127400 117476
rect 157816 117532 157880 117536
rect 157816 117476 157820 117532
rect 157820 117476 157876 117532
rect 157876 117476 157880 117532
rect 157816 117472 157880 117476
rect 157896 117532 157960 117536
rect 157896 117476 157900 117532
rect 157900 117476 157956 117532
rect 157956 117476 157960 117532
rect 157896 117472 157960 117476
rect 157976 117532 158040 117536
rect 157976 117476 157980 117532
rect 157980 117476 158036 117532
rect 158036 117476 158040 117532
rect 157976 117472 158040 117476
rect 158056 117532 158120 117536
rect 158056 117476 158060 117532
rect 158060 117476 158116 117532
rect 158116 117476 158120 117532
rect 158056 117472 158120 117476
rect 19576 116988 19640 116992
rect 19576 116932 19580 116988
rect 19580 116932 19636 116988
rect 19636 116932 19640 116988
rect 19576 116928 19640 116932
rect 19656 116988 19720 116992
rect 19656 116932 19660 116988
rect 19660 116932 19716 116988
rect 19716 116932 19720 116988
rect 19656 116928 19720 116932
rect 19736 116988 19800 116992
rect 19736 116932 19740 116988
rect 19740 116932 19796 116988
rect 19796 116932 19800 116988
rect 19736 116928 19800 116932
rect 19816 116988 19880 116992
rect 19816 116932 19820 116988
rect 19820 116932 19876 116988
rect 19876 116932 19880 116988
rect 19816 116928 19880 116932
rect 50296 116988 50360 116992
rect 50296 116932 50300 116988
rect 50300 116932 50356 116988
rect 50356 116932 50360 116988
rect 50296 116928 50360 116932
rect 50376 116988 50440 116992
rect 50376 116932 50380 116988
rect 50380 116932 50436 116988
rect 50436 116932 50440 116988
rect 50376 116928 50440 116932
rect 50456 116988 50520 116992
rect 50456 116932 50460 116988
rect 50460 116932 50516 116988
rect 50516 116932 50520 116988
rect 50456 116928 50520 116932
rect 50536 116988 50600 116992
rect 50536 116932 50540 116988
rect 50540 116932 50596 116988
rect 50596 116932 50600 116988
rect 50536 116928 50600 116932
rect 81016 116988 81080 116992
rect 81016 116932 81020 116988
rect 81020 116932 81076 116988
rect 81076 116932 81080 116988
rect 81016 116928 81080 116932
rect 81096 116988 81160 116992
rect 81096 116932 81100 116988
rect 81100 116932 81156 116988
rect 81156 116932 81160 116988
rect 81096 116928 81160 116932
rect 81176 116988 81240 116992
rect 81176 116932 81180 116988
rect 81180 116932 81236 116988
rect 81236 116932 81240 116988
rect 81176 116928 81240 116932
rect 81256 116988 81320 116992
rect 81256 116932 81260 116988
rect 81260 116932 81316 116988
rect 81316 116932 81320 116988
rect 81256 116928 81320 116932
rect 111736 116988 111800 116992
rect 111736 116932 111740 116988
rect 111740 116932 111796 116988
rect 111796 116932 111800 116988
rect 111736 116928 111800 116932
rect 111816 116988 111880 116992
rect 111816 116932 111820 116988
rect 111820 116932 111876 116988
rect 111876 116932 111880 116988
rect 111816 116928 111880 116932
rect 111896 116988 111960 116992
rect 111896 116932 111900 116988
rect 111900 116932 111956 116988
rect 111956 116932 111960 116988
rect 111896 116928 111960 116932
rect 111976 116988 112040 116992
rect 111976 116932 111980 116988
rect 111980 116932 112036 116988
rect 112036 116932 112040 116988
rect 111976 116928 112040 116932
rect 142456 116988 142520 116992
rect 142456 116932 142460 116988
rect 142460 116932 142516 116988
rect 142516 116932 142520 116988
rect 142456 116928 142520 116932
rect 142536 116988 142600 116992
rect 142536 116932 142540 116988
rect 142540 116932 142596 116988
rect 142596 116932 142600 116988
rect 142536 116928 142600 116932
rect 142616 116988 142680 116992
rect 142616 116932 142620 116988
rect 142620 116932 142676 116988
rect 142676 116932 142680 116988
rect 142616 116928 142680 116932
rect 142696 116988 142760 116992
rect 142696 116932 142700 116988
rect 142700 116932 142756 116988
rect 142756 116932 142760 116988
rect 142696 116928 142760 116932
rect 173176 116988 173240 116992
rect 173176 116932 173180 116988
rect 173180 116932 173236 116988
rect 173236 116932 173240 116988
rect 173176 116928 173240 116932
rect 173256 116988 173320 116992
rect 173256 116932 173260 116988
rect 173260 116932 173316 116988
rect 173316 116932 173320 116988
rect 173256 116928 173320 116932
rect 173336 116988 173400 116992
rect 173336 116932 173340 116988
rect 173340 116932 173396 116988
rect 173396 116932 173400 116988
rect 173336 116928 173400 116932
rect 173416 116988 173480 116992
rect 173416 116932 173420 116988
rect 173420 116932 173476 116988
rect 173476 116932 173480 116988
rect 173416 116928 173480 116932
rect 4216 116444 4280 116448
rect 4216 116388 4220 116444
rect 4220 116388 4276 116444
rect 4276 116388 4280 116444
rect 4216 116384 4280 116388
rect 4296 116444 4360 116448
rect 4296 116388 4300 116444
rect 4300 116388 4356 116444
rect 4356 116388 4360 116444
rect 4296 116384 4360 116388
rect 4376 116444 4440 116448
rect 4376 116388 4380 116444
rect 4380 116388 4436 116444
rect 4436 116388 4440 116444
rect 4376 116384 4440 116388
rect 4456 116444 4520 116448
rect 4456 116388 4460 116444
rect 4460 116388 4516 116444
rect 4516 116388 4520 116444
rect 4456 116384 4520 116388
rect 34936 116444 35000 116448
rect 34936 116388 34940 116444
rect 34940 116388 34996 116444
rect 34996 116388 35000 116444
rect 34936 116384 35000 116388
rect 35016 116444 35080 116448
rect 35016 116388 35020 116444
rect 35020 116388 35076 116444
rect 35076 116388 35080 116444
rect 35016 116384 35080 116388
rect 35096 116444 35160 116448
rect 35096 116388 35100 116444
rect 35100 116388 35156 116444
rect 35156 116388 35160 116444
rect 35096 116384 35160 116388
rect 35176 116444 35240 116448
rect 35176 116388 35180 116444
rect 35180 116388 35236 116444
rect 35236 116388 35240 116444
rect 35176 116384 35240 116388
rect 65656 116444 65720 116448
rect 65656 116388 65660 116444
rect 65660 116388 65716 116444
rect 65716 116388 65720 116444
rect 65656 116384 65720 116388
rect 65736 116444 65800 116448
rect 65736 116388 65740 116444
rect 65740 116388 65796 116444
rect 65796 116388 65800 116444
rect 65736 116384 65800 116388
rect 65816 116444 65880 116448
rect 65816 116388 65820 116444
rect 65820 116388 65876 116444
rect 65876 116388 65880 116444
rect 65816 116384 65880 116388
rect 65896 116444 65960 116448
rect 65896 116388 65900 116444
rect 65900 116388 65956 116444
rect 65956 116388 65960 116444
rect 65896 116384 65960 116388
rect 96376 116444 96440 116448
rect 96376 116388 96380 116444
rect 96380 116388 96436 116444
rect 96436 116388 96440 116444
rect 96376 116384 96440 116388
rect 96456 116444 96520 116448
rect 96456 116388 96460 116444
rect 96460 116388 96516 116444
rect 96516 116388 96520 116444
rect 96456 116384 96520 116388
rect 96536 116444 96600 116448
rect 96536 116388 96540 116444
rect 96540 116388 96596 116444
rect 96596 116388 96600 116444
rect 96536 116384 96600 116388
rect 96616 116444 96680 116448
rect 96616 116388 96620 116444
rect 96620 116388 96676 116444
rect 96676 116388 96680 116444
rect 96616 116384 96680 116388
rect 127096 116444 127160 116448
rect 127096 116388 127100 116444
rect 127100 116388 127156 116444
rect 127156 116388 127160 116444
rect 127096 116384 127160 116388
rect 127176 116444 127240 116448
rect 127176 116388 127180 116444
rect 127180 116388 127236 116444
rect 127236 116388 127240 116444
rect 127176 116384 127240 116388
rect 127256 116444 127320 116448
rect 127256 116388 127260 116444
rect 127260 116388 127316 116444
rect 127316 116388 127320 116444
rect 127256 116384 127320 116388
rect 127336 116444 127400 116448
rect 127336 116388 127340 116444
rect 127340 116388 127396 116444
rect 127396 116388 127400 116444
rect 127336 116384 127400 116388
rect 157816 116444 157880 116448
rect 157816 116388 157820 116444
rect 157820 116388 157876 116444
rect 157876 116388 157880 116444
rect 157816 116384 157880 116388
rect 157896 116444 157960 116448
rect 157896 116388 157900 116444
rect 157900 116388 157956 116444
rect 157956 116388 157960 116444
rect 157896 116384 157960 116388
rect 157976 116444 158040 116448
rect 157976 116388 157980 116444
rect 157980 116388 158036 116444
rect 158036 116388 158040 116444
rect 157976 116384 158040 116388
rect 158056 116444 158120 116448
rect 158056 116388 158060 116444
rect 158060 116388 158116 116444
rect 158116 116388 158120 116444
rect 158056 116384 158120 116388
rect 19576 115900 19640 115904
rect 19576 115844 19580 115900
rect 19580 115844 19636 115900
rect 19636 115844 19640 115900
rect 19576 115840 19640 115844
rect 19656 115900 19720 115904
rect 19656 115844 19660 115900
rect 19660 115844 19716 115900
rect 19716 115844 19720 115900
rect 19656 115840 19720 115844
rect 19736 115900 19800 115904
rect 19736 115844 19740 115900
rect 19740 115844 19796 115900
rect 19796 115844 19800 115900
rect 19736 115840 19800 115844
rect 19816 115900 19880 115904
rect 19816 115844 19820 115900
rect 19820 115844 19876 115900
rect 19876 115844 19880 115900
rect 19816 115840 19880 115844
rect 50296 115900 50360 115904
rect 50296 115844 50300 115900
rect 50300 115844 50356 115900
rect 50356 115844 50360 115900
rect 50296 115840 50360 115844
rect 50376 115900 50440 115904
rect 50376 115844 50380 115900
rect 50380 115844 50436 115900
rect 50436 115844 50440 115900
rect 50376 115840 50440 115844
rect 50456 115900 50520 115904
rect 50456 115844 50460 115900
rect 50460 115844 50516 115900
rect 50516 115844 50520 115900
rect 50456 115840 50520 115844
rect 50536 115900 50600 115904
rect 50536 115844 50540 115900
rect 50540 115844 50596 115900
rect 50596 115844 50600 115900
rect 50536 115840 50600 115844
rect 81016 115900 81080 115904
rect 81016 115844 81020 115900
rect 81020 115844 81076 115900
rect 81076 115844 81080 115900
rect 81016 115840 81080 115844
rect 81096 115900 81160 115904
rect 81096 115844 81100 115900
rect 81100 115844 81156 115900
rect 81156 115844 81160 115900
rect 81096 115840 81160 115844
rect 81176 115900 81240 115904
rect 81176 115844 81180 115900
rect 81180 115844 81236 115900
rect 81236 115844 81240 115900
rect 81176 115840 81240 115844
rect 81256 115900 81320 115904
rect 81256 115844 81260 115900
rect 81260 115844 81316 115900
rect 81316 115844 81320 115900
rect 81256 115840 81320 115844
rect 111736 115900 111800 115904
rect 111736 115844 111740 115900
rect 111740 115844 111796 115900
rect 111796 115844 111800 115900
rect 111736 115840 111800 115844
rect 111816 115900 111880 115904
rect 111816 115844 111820 115900
rect 111820 115844 111876 115900
rect 111876 115844 111880 115900
rect 111816 115840 111880 115844
rect 111896 115900 111960 115904
rect 111896 115844 111900 115900
rect 111900 115844 111956 115900
rect 111956 115844 111960 115900
rect 111896 115840 111960 115844
rect 111976 115900 112040 115904
rect 111976 115844 111980 115900
rect 111980 115844 112036 115900
rect 112036 115844 112040 115900
rect 111976 115840 112040 115844
rect 142456 115900 142520 115904
rect 142456 115844 142460 115900
rect 142460 115844 142516 115900
rect 142516 115844 142520 115900
rect 142456 115840 142520 115844
rect 142536 115900 142600 115904
rect 142536 115844 142540 115900
rect 142540 115844 142596 115900
rect 142596 115844 142600 115900
rect 142536 115840 142600 115844
rect 142616 115900 142680 115904
rect 142616 115844 142620 115900
rect 142620 115844 142676 115900
rect 142676 115844 142680 115900
rect 142616 115840 142680 115844
rect 142696 115900 142760 115904
rect 142696 115844 142700 115900
rect 142700 115844 142756 115900
rect 142756 115844 142760 115900
rect 142696 115840 142760 115844
rect 173176 115900 173240 115904
rect 173176 115844 173180 115900
rect 173180 115844 173236 115900
rect 173236 115844 173240 115900
rect 173176 115840 173240 115844
rect 173256 115900 173320 115904
rect 173256 115844 173260 115900
rect 173260 115844 173316 115900
rect 173316 115844 173320 115900
rect 173256 115840 173320 115844
rect 173336 115900 173400 115904
rect 173336 115844 173340 115900
rect 173340 115844 173396 115900
rect 173396 115844 173400 115900
rect 173336 115840 173400 115844
rect 173416 115900 173480 115904
rect 173416 115844 173420 115900
rect 173420 115844 173476 115900
rect 173476 115844 173480 115900
rect 173416 115840 173480 115844
rect 4216 115356 4280 115360
rect 4216 115300 4220 115356
rect 4220 115300 4276 115356
rect 4276 115300 4280 115356
rect 4216 115296 4280 115300
rect 4296 115356 4360 115360
rect 4296 115300 4300 115356
rect 4300 115300 4356 115356
rect 4356 115300 4360 115356
rect 4296 115296 4360 115300
rect 4376 115356 4440 115360
rect 4376 115300 4380 115356
rect 4380 115300 4436 115356
rect 4436 115300 4440 115356
rect 4376 115296 4440 115300
rect 4456 115356 4520 115360
rect 4456 115300 4460 115356
rect 4460 115300 4516 115356
rect 4516 115300 4520 115356
rect 4456 115296 4520 115300
rect 34936 115356 35000 115360
rect 34936 115300 34940 115356
rect 34940 115300 34996 115356
rect 34996 115300 35000 115356
rect 34936 115296 35000 115300
rect 35016 115356 35080 115360
rect 35016 115300 35020 115356
rect 35020 115300 35076 115356
rect 35076 115300 35080 115356
rect 35016 115296 35080 115300
rect 35096 115356 35160 115360
rect 35096 115300 35100 115356
rect 35100 115300 35156 115356
rect 35156 115300 35160 115356
rect 35096 115296 35160 115300
rect 35176 115356 35240 115360
rect 35176 115300 35180 115356
rect 35180 115300 35236 115356
rect 35236 115300 35240 115356
rect 35176 115296 35240 115300
rect 65656 115356 65720 115360
rect 65656 115300 65660 115356
rect 65660 115300 65716 115356
rect 65716 115300 65720 115356
rect 65656 115296 65720 115300
rect 65736 115356 65800 115360
rect 65736 115300 65740 115356
rect 65740 115300 65796 115356
rect 65796 115300 65800 115356
rect 65736 115296 65800 115300
rect 65816 115356 65880 115360
rect 65816 115300 65820 115356
rect 65820 115300 65876 115356
rect 65876 115300 65880 115356
rect 65816 115296 65880 115300
rect 65896 115356 65960 115360
rect 65896 115300 65900 115356
rect 65900 115300 65956 115356
rect 65956 115300 65960 115356
rect 65896 115296 65960 115300
rect 96376 115356 96440 115360
rect 96376 115300 96380 115356
rect 96380 115300 96436 115356
rect 96436 115300 96440 115356
rect 96376 115296 96440 115300
rect 96456 115356 96520 115360
rect 96456 115300 96460 115356
rect 96460 115300 96516 115356
rect 96516 115300 96520 115356
rect 96456 115296 96520 115300
rect 96536 115356 96600 115360
rect 96536 115300 96540 115356
rect 96540 115300 96596 115356
rect 96596 115300 96600 115356
rect 96536 115296 96600 115300
rect 96616 115356 96680 115360
rect 96616 115300 96620 115356
rect 96620 115300 96676 115356
rect 96676 115300 96680 115356
rect 96616 115296 96680 115300
rect 127096 115356 127160 115360
rect 127096 115300 127100 115356
rect 127100 115300 127156 115356
rect 127156 115300 127160 115356
rect 127096 115296 127160 115300
rect 127176 115356 127240 115360
rect 127176 115300 127180 115356
rect 127180 115300 127236 115356
rect 127236 115300 127240 115356
rect 127176 115296 127240 115300
rect 127256 115356 127320 115360
rect 127256 115300 127260 115356
rect 127260 115300 127316 115356
rect 127316 115300 127320 115356
rect 127256 115296 127320 115300
rect 127336 115356 127400 115360
rect 127336 115300 127340 115356
rect 127340 115300 127396 115356
rect 127396 115300 127400 115356
rect 127336 115296 127400 115300
rect 157816 115356 157880 115360
rect 157816 115300 157820 115356
rect 157820 115300 157876 115356
rect 157876 115300 157880 115356
rect 157816 115296 157880 115300
rect 157896 115356 157960 115360
rect 157896 115300 157900 115356
rect 157900 115300 157956 115356
rect 157956 115300 157960 115356
rect 157896 115296 157960 115300
rect 157976 115356 158040 115360
rect 157976 115300 157980 115356
rect 157980 115300 158036 115356
rect 158036 115300 158040 115356
rect 157976 115296 158040 115300
rect 158056 115356 158120 115360
rect 158056 115300 158060 115356
rect 158060 115300 158116 115356
rect 158116 115300 158120 115356
rect 158056 115296 158120 115300
rect 19576 114812 19640 114816
rect 19576 114756 19580 114812
rect 19580 114756 19636 114812
rect 19636 114756 19640 114812
rect 19576 114752 19640 114756
rect 19656 114812 19720 114816
rect 19656 114756 19660 114812
rect 19660 114756 19716 114812
rect 19716 114756 19720 114812
rect 19656 114752 19720 114756
rect 19736 114812 19800 114816
rect 19736 114756 19740 114812
rect 19740 114756 19796 114812
rect 19796 114756 19800 114812
rect 19736 114752 19800 114756
rect 19816 114812 19880 114816
rect 19816 114756 19820 114812
rect 19820 114756 19876 114812
rect 19876 114756 19880 114812
rect 19816 114752 19880 114756
rect 50296 114812 50360 114816
rect 50296 114756 50300 114812
rect 50300 114756 50356 114812
rect 50356 114756 50360 114812
rect 50296 114752 50360 114756
rect 50376 114812 50440 114816
rect 50376 114756 50380 114812
rect 50380 114756 50436 114812
rect 50436 114756 50440 114812
rect 50376 114752 50440 114756
rect 50456 114812 50520 114816
rect 50456 114756 50460 114812
rect 50460 114756 50516 114812
rect 50516 114756 50520 114812
rect 50456 114752 50520 114756
rect 50536 114812 50600 114816
rect 50536 114756 50540 114812
rect 50540 114756 50596 114812
rect 50596 114756 50600 114812
rect 50536 114752 50600 114756
rect 81016 114812 81080 114816
rect 81016 114756 81020 114812
rect 81020 114756 81076 114812
rect 81076 114756 81080 114812
rect 81016 114752 81080 114756
rect 81096 114812 81160 114816
rect 81096 114756 81100 114812
rect 81100 114756 81156 114812
rect 81156 114756 81160 114812
rect 81096 114752 81160 114756
rect 81176 114812 81240 114816
rect 81176 114756 81180 114812
rect 81180 114756 81236 114812
rect 81236 114756 81240 114812
rect 81176 114752 81240 114756
rect 81256 114812 81320 114816
rect 81256 114756 81260 114812
rect 81260 114756 81316 114812
rect 81316 114756 81320 114812
rect 81256 114752 81320 114756
rect 111736 114812 111800 114816
rect 111736 114756 111740 114812
rect 111740 114756 111796 114812
rect 111796 114756 111800 114812
rect 111736 114752 111800 114756
rect 111816 114812 111880 114816
rect 111816 114756 111820 114812
rect 111820 114756 111876 114812
rect 111876 114756 111880 114812
rect 111816 114752 111880 114756
rect 111896 114812 111960 114816
rect 111896 114756 111900 114812
rect 111900 114756 111956 114812
rect 111956 114756 111960 114812
rect 111896 114752 111960 114756
rect 111976 114812 112040 114816
rect 111976 114756 111980 114812
rect 111980 114756 112036 114812
rect 112036 114756 112040 114812
rect 111976 114752 112040 114756
rect 142456 114812 142520 114816
rect 142456 114756 142460 114812
rect 142460 114756 142516 114812
rect 142516 114756 142520 114812
rect 142456 114752 142520 114756
rect 142536 114812 142600 114816
rect 142536 114756 142540 114812
rect 142540 114756 142596 114812
rect 142596 114756 142600 114812
rect 142536 114752 142600 114756
rect 142616 114812 142680 114816
rect 142616 114756 142620 114812
rect 142620 114756 142676 114812
rect 142676 114756 142680 114812
rect 142616 114752 142680 114756
rect 142696 114812 142760 114816
rect 142696 114756 142700 114812
rect 142700 114756 142756 114812
rect 142756 114756 142760 114812
rect 142696 114752 142760 114756
rect 173176 114812 173240 114816
rect 173176 114756 173180 114812
rect 173180 114756 173236 114812
rect 173236 114756 173240 114812
rect 173176 114752 173240 114756
rect 173256 114812 173320 114816
rect 173256 114756 173260 114812
rect 173260 114756 173316 114812
rect 173316 114756 173320 114812
rect 173256 114752 173320 114756
rect 173336 114812 173400 114816
rect 173336 114756 173340 114812
rect 173340 114756 173396 114812
rect 173396 114756 173400 114812
rect 173336 114752 173400 114756
rect 173416 114812 173480 114816
rect 173416 114756 173420 114812
rect 173420 114756 173476 114812
rect 173476 114756 173480 114812
rect 173416 114752 173480 114756
rect 4216 114268 4280 114272
rect 4216 114212 4220 114268
rect 4220 114212 4276 114268
rect 4276 114212 4280 114268
rect 4216 114208 4280 114212
rect 4296 114268 4360 114272
rect 4296 114212 4300 114268
rect 4300 114212 4356 114268
rect 4356 114212 4360 114268
rect 4296 114208 4360 114212
rect 4376 114268 4440 114272
rect 4376 114212 4380 114268
rect 4380 114212 4436 114268
rect 4436 114212 4440 114268
rect 4376 114208 4440 114212
rect 4456 114268 4520 114272
rect 4456 114212 4460 114268
rect 4460 114212 4516 114268
rect 4516 114212 4520 114268
rect 4456 114208 4520 114212
rect 34936 114268 35000 114272
rect 34936 114212 34940 114268
rect 34940 114212 34996 114268
rect 34996 114212 35000 114268
rect 34936 114208 35000 114212
rect 35016 114268 35080 114272
rect 35016 114212 35020 114268
rect 35020 114212 35076 114268
rect 35076 114212 35080 114268
rect 35016 114208 35080 114212
rect 35096 114268 35160 114272
rect 35096 114212 35100 114268
rect 35100 114212 35156 114268
rect 35156 114212 35160 114268
rect 35096 114208 35160 114212
rect 35176 114268 35240 114272
rect 35176 114212 35180 114268
rect 35180 114212 35236 114268
rect 35236 114212 35240 114268
rect 35176 114208 35240 114212
rect 65656 114268 65720 114272
rect 65656 114212 65660 114268
rect 65660 114212 65716 114268
rect 65716 114212 65720 114268
rect 65656 114208 65720 114212
rect 65736 114268 65800 114272
rect 65736 114212 65740 114268
rect 65740 114212 65796 114268
rect 65796 114212 65800 114268
rect 65736 114208 65800 114212
rect 65816 114268 65880 114272
rect 65816 114212 65820 114268
rect 65820 114212 65876 114268
rect 65876 114212 65880 114268
rect 65816 114208 65880 114212
rect 65896 114268 65960 114272
rect 65896 114212 65900 114268
rect 65900 114212 65956 114268
rect 65956 114212 65960 114268
rect 65896 114208 65960 114212
rect 96376 114268 96440 114272
rect 96376 114212 96380 114268
rect 96380 114212 96436 114268
rect 96436 114212 96440 114268
rect 96376 114208 96440 114212
rect 96456 114268 96520 114272
rect 96456 114212 96460 114268
rect 96460 114212 96516 114268
rect 96516 114212 96520 114268
rect 96456 114208 96520 114212
rect 96536 114268 96600 114272
rect 96536 114212 96540 114268
rect 96540 114212 96596 114268
rect 96596 114212 96600 114268
rect 96536 114208 96600 114212
rect 96616 114268 96680 114272
rect 96616 114212 96620 114268
rect 96620 114212 96676 114268
rect 96676 114212 96680 114268
rect 96616 114208 96680 114212
rect 127096 114268 127160 114272
rect 127096 114212 127100 114268
rect 127100 114212 127156 114268
rect 127156 114212 127160 114268
rect 127096 114208 127160 114212
rect 127176 114268 127240 114272
rect 127176 114212 127180 114268
rect 127180 114212 127236 114268
rect 127236 114212 127240 114268
rect 127176 114208 127240 114212
rect 127256 114268 127320 114272
rect 127256 114212 127260 114268
rect 127260 114212 127316 114268
rect 127316 114212 127320 114268
rect 127256 114208 127320 114212
rect 127336 114268 127400 114272
rect 127336 114212 127340 114268
rect 127340 114212 127396 114268
rect 127396 114212 127400 114268
rect 127336 114208 127400 114212
rect 157816 114268 157880 114272
rect 157816 114212 157820 114268
rect 157820 114212 157876 114268
rect 157876 114212 157880 114268
rect 157816 114208 157880 114212
rect 157896 114268 157960 114272
rect 157896 114212 157900 114268
rect 157900 114212 157956 114268
rect 157956 114212 157960 114268
rect 157896 114208 157960 114212
rect 157976 114268 158040 114272
rect 157976 114212 157980 114268
rect 157980 114212 158036 114268
rect 158036 114212 158040 114268
rect 157976 114208 158040 114212
rect 158056 114268 158120 114272
rect 158056 114212 158060 114268
rect 158060 114212 158116 114268
rect 158116 114212 158120 114268
rect 158056 114208 158120 114212
rect 19576 113724 19640 113728
rect 19576 113668 19580 113724
rect 19580 113668 19636 113724
rect 19636 113668 19640 113724
rect 19576 113664 19640 113668
rect 19656 113724 19720 113728
rect 19656 113668 19660 113724
rect 19660 113668 19716 113724
rect 19716 113668 19720 113724
rect 19656 113664 19720 113668
rect 19736 113724 19800 113728
rect 19736 113668 19740 113724
rect 19740 113668 19796 113724
rect 19796 113668 19800 113724
rect 19736 113664 19800 113668
rect 19816 113724 19880 113728
rect 19816 113668 19820 113724
rect 19820 113668 19876 113724
rect 19876 113668 19880 113724
rect 19816 113664 19880 113668
rect 50296 113724 50360 113728
rect 50296 113668 50300 113724
rect 50300 113668 50356 113724
rect 50356 113668 50360 113724
rect 50296 113664 50360 113668
rect 50376 113724 50440 113728
rect 50376 113668 50380 113724
rect 50380 113668 50436 113724
rect 50436 113668 50440 113724
rect 50376 113664 50440 113668
rect 50456 113724 50520 113728
rect 50456 113668 50460 113724
rect 50460 113668 50516 113724
rect 50516 113668 50520 113724
rect 50456 113664 50520 113668
rect 50536 113724 50600 113728
rect 50536 113668 50540 113724
rect 50540 113668 50596 113724
rect 50596 113668 50600 113724
rect 50536 113664 50600 113668
rect 81016 113724 81080 113728
rect 81016 113668 81020 113724
rect 81020 113668 81076 113724
rect 81076 113668 81080 113724
rect 81016 113664 81080 113668
rect 81096 113724 81160 113728
rect 81096 113668 81100 113724
rect 81100 113668 81156 113724
rect 81156 113668 81160 113724
rect 81096 113664 81160 113668
rect 81176 113724 81240 113728
rect 81176 113668 81180 113724
rect 81180 113668 81236 113724
rect 81236 113668 81240 113724
rect 81176 113664 81240 113668
rect 81256 113724 81320 113728
rect 81256 113668 81260 113724
rect 81260 113668 81316 113724
rect 81316 113668 81320 113724
rect 81256 113664 81320 113668
rect 111736 113724 111800 113728
rect 111736 113668 111740 113724
rect 111740 113668 111796 113724
rect 111796 113668 111800 113724
rect 111736 113664 111800 113668
rect 111816 113724 111880 113728
rect 111816 113668 111820 113724
rect 111820 113668 111876 113724
rect 111876 113668 111880 113724
rect 111816 113664 111880 113668
rect 111896 113724 111960 113728
rect 111896 113668 111900 113724
rect 111900 113668 111956 113724
rect 111956 113668 111960 113724
rect 111896 113664 111960 113668
rect 111976 113724 112040 113728
rect 111976 113668 111980 113724
rect 111980 113668 112036 113724
rect 112036 113668 112040 113724
rect 111976 113664 112040 113668
rect 142456 113724 142520 113728
rect 142456 113668 142460 113724
rect 142460 113668 142516 113724
rect 142516 113668 142520 113724
rect 142456 113664 142520 113668
rect 142536 113724 142600 113728
rect 142536 113668 142540 113724
rect 142540 113668 142596 113724
rect 142596 113668 142600 113724
rect 142536 113664 142600 113668
rect 142616 113724 142680 113728
rect 142616 113668 142620 113724
rect 142620 113668 142676 113724
rect 142676 113668 142680 113724
rect 142616 113664 142680 113668
rect 142696 113724 142760 113728
rect 142696 113668 142700 113724
rect 142700 113668 142756 113724
rect 142756 113668 142760 113724
rect 142696 113664 142760 113668
rect 173176 113724 173240 113728
rect 173176 113668 173180 113724
rect 173180 113668 173236 113724
rect 173236 113668 173240 113724
rect 173176 113664 173240 113668
rect 173256 113724 173320 113728
rect 173256 113668 173260 113724
rect 173260 113668 173316 113724
rect 173316 113668 173320 113724
rect 173256 113664 173320 113668
rect 173336 113724 173400 113728
rect 173336 113668 173340 113724
rect 173340 113668 173396 113724
rect 173396 113668 173400 113724
rect 173336 113664 173400 113668
rect 173416 113724 173480 113728
rect 173416 113668 173420 113724
rect 173420 113668 173476 113724
rect 173476 113668 173480 113724
rect 173416 113664 173480 113668
rect 4216 113180 4280 113184
rect 4216 113124 4220 113180
rect 4220 113124 4276 113180
rect 4276 113124 4280 113180
rect 4216 113120 4280 113124
rect 4296 113180 4360 113184
rect 4296 113124 4300 113180
rect 4300 113124 4356 113180
rect 4356 113124 4360 113180
rect 4296 113120 4360 113124
rect 4376 113180 4440 113184
rect 4376 113124 4380 113180
rect 4380 113124 4436 113180
rect 4436 113124 4440 113180
rect 4376 113120 4440 113124
rect 4456 113180 4520 113184
rect 4456 113124 4460 113180
rect 4460 113124 4516 113180
rect 4516 113124 4520 113180
rect 4456 113120 4520 113124
rect 34936 113180 35000 113184
rect 34936 113124 34940 113180
rect 34940 113124 34996 113180
rect 34996 113124 35000 113180
rect 34936 113120 35000 113124
rect 35016 113180 35080 113184
rect 35016 113124 35020 113180
rect 35020 113124 35076 113180
rect 35076 113124 35080 113180
rect 35016 113120 35080 113124
rect 35096 113180 35160 113184
rect 35096 113124 35100 113180
rect 35100 113124 35156 113180
rect 35156 113124 35160 113180
rect 35096 113120 35160 113124
rect 35176 113180 35240 113184
rect 35176 113124 35180 113180
rect 35180 113124 35236 113180
rect 35236 113124 35240 113180
rect 35176 113120 35240 113124
rect 65656 113180 65720 113184
rect 65656 113124 65660 113180
rect 65660 113124 65716 113180
rect 65716 113124 65720 113180
rect 65656 113120 65720 113124
rect 65736 113180 65800 113184
rect 65736 113124 65740 113180
rect 65740 113124 65796 113180
rect 65796 113124 65800 113180
rect 65736 113120 65800 113124
rect 65816 113180 65880 113184
rect 65816 113124 65820 113180
rect 65820 113124 65876 113180
rect 65876 113124 65880 113180
rect 65816 113120 65880 113124
rect 65896 113180 65960 113184
rect 65896 113124 65900 113180
rect 65900 113124 65956 113180
rect 65956 113124 65960 113180
rect 65896 113120 65960 113124
rect 96376 113180 96440 113184
rect 96376 113124 96380 113180
rect 96380 113124 96436 113180
rect 96436 113124 96440 113180
rect 96376 113120 96440 113124
rect 96456 113180 96520 113184
rect 96456 113124 96460 113180
rect 96460 113124 96516 113180
rect 96516 113124 96520 113180
rect 96456 113120 96520 113124
rect 96536 113180 96600 113184
rect 96536 113124 96540 113180
rect 96540 113124 96596 113180
rect 96596 113124 96600 113180
rect 96536 113120 96600 113124
rect 96616 113180 96680 113184
rect 96616 113124 96620 113180
rect 96620 113124 96676 113180
rect 96676 113124 96680 113180
rect 96616 113120 96680 113124
rect 127096 113180 127160 113184
rect 127096 113124 127100 113180
rect 127100 113124 127156 113180
rect 127156 113124 127160 113180
rect 127096 113120 127160 113124
rect 127176 113180 127240 113184
rect 127176 113124 127180 113180
rect 127180 113124 127236 113180
rect 127236 113124 127240 113180
rect 127176 113120 127240 113124
rect 127256 113180 127320 113184
rect 127256 113124 127260 113180
rect 127260 113124 127316 113180
rect 127316 113124 127320 113180
rect 127256 113120 127320 113124
rect 127336 113180 127400 113184
rect 127336 113124 127340 113180
rect 127340 113124 127396 113180
rect 127396 113124 127400 113180
rect 127336 113120 127400 113124
rect 157816 113180 157880 113184
rect 157816 113124 157820 113180
rect 157820 113124 157876 113180
rect 157876 113124 157880 113180
rect 157816 113120 157880 113124
rect 157896 113180 157960 113184
rect 157896 113124 157900 113180
rect 157900 113124 157956 113180
rect 157956 113124 157960 113180
rect 157896 113120 157960 113124
rect 157976 113180 158040 113184
rect 157976 113124 157980 113180
rect 157980 113124 158036 113180
rect 158036 113124 158040 113180
rect 157976 113120 158040 113124
rect 158056 113180 158120 113184
rect 158056 113124 158060 113180
rect 158060 113124 158116 113180
rect 158116 113124 158120 113180
rect 158056 113120 158120 113124
rect 19576 112636 19640 112640
rect 19576 112580 19580 112636
rect 19580 112580 19636 112636
rect 19636 112580 19640 112636
rect 19576 112576 19640 112580
rect 19656 112636 19720 112640
rect 19656 112580 19660 112636
rect 19660 112580 19716 112636
rect 19716 112580 19720 112636
rect 19656 112576 19720 112580
rect 19736 112636 19800 112640
rect 19736 112580 19740 112636
rect 19740 112580 19796 112636
rect 19796 112580 19800 112636
rect 19736 112576 19800 112580
rect 19816 112636 19880 112640
rect 19816 112580 19820 112636
rect 19820 112580 19876 112636
rect 19876 112580 19880 112636
rect 19816 112576 19880 112580
rect 50296 112636 50360 112640
rect 50296 112580 50300 112636
rect 50300 112580 50356 112636
rect 50356 112580 50360 112636
rect 50296 112576 50360 112580
rect 50376 112636 50440 112640
rect 50376 112580 50380 112636
rect 50380 112580 50436 112636
rect 50436 112580 50440 112636
rect 50376 112576 50440 112580
rect 50456 112636 50520 112640
rect 50456 112580 50460 112636
rect 50460 112580 50516 112636
rect 50516 112580 50520 112636
rect 50456 112576 50520 112580
rect 50536 112636 50600 112640
rect 50536 112580 50540 112636
rect 50540 112580 50596 112636
rect 50596 112580 50600 112636
rect 50536 112576 50600 112580
rect 81016 112636 81080 112640
rect 81016 112580 81020 112636
rect 81020 112580 81076 112636
rect 81076 112580 81080 112636
rect 81016 112576 81080 112580
rect 81096 112636 81160 112640
rect 81096 112580 81100 112636
rect 81100 112580 81156 112636
rect 81156 112580 81160 112636
rect 81096 112576 81160 112580
rect 81176 112636 81240 112640
rect 81176 112580 81180 112636
rect 81180 112580 81236 112636
rect 81236 112580 81240 112636
rect 81176 112576 81240 112580
rect 81256 112636 81320 112640
rect 81256 112580 81260 112636
rect 81260 112580 81316 112636
rect 81316 112580 81320 112636
rect 81256 112576 81320 112580
rect 111736 112636 111800 112640
rect 111736 112580 111740 112636
rect 111740 112580 111796 112636
rect 111796 112580 111800 112636
rect 111736 112576 111800 112580
rect 111816 112636 111880 112640
rect 111816 112580 111820 112636
rect 111820 112580 111876 112636
rect 111876 112580 111880 112636
rect 111816 112576 111880 112580
rect 111896 112636 111960 112640
rect 111896 112580 111900 112636
rect 111900 112580 111956 112636
rect 111956 112580 111960 112636
rect 111896 112576 111960 112580
rect 111976 112636 112040 112640
rect 111976 112580 111980 112636
rect 111980 112580 112036 112636
rect 112036 112580 112040 112636
rect 111976 112576 112040 112580
rect 142456 112636 142520 112640
rect 142456 112580 142460 112636
rect 142460 112580 142516 112636
rect 142516 112580 142520 112636
rect 142456 112576 142520 112580
rect 142536 112636 142600 112640
rect 142536 112580 142540 112636
rect 142540 112580 142596 112636
rect 142596 112580 142600 112636
rect 142536 112576 142600 112580
rect 142616 112636 142680 112640
rect 142616 112580 142620 112636
rect 142620 112580 142676 112636
rect 142676 112580 142680 112636
rect 142616 112576 142680 112580
rect 142696 112636 142760 112640
rect 142696 112580 142700 112636
rect 142700 112580 142756 112636
rect 142756 112580 142760 112636
rect 142696 112576 142760 112580
rect 173176 112636 173240 112640
rect 173176 112580 173180 112636
rect 173180 112580 173236 112636
rect 173236 112580 173240 112636
rect 173176 112576 173240 112580
rect 173256 112636 173320 112640
rect 173256 112580 173260 112636
rect 173260 112580 173316 112636
rect 173316 112580 173320 112636
rect 173256 112576 173320 112580
rect 173336 112636 173400 112640
rect 173336 112580 173340 112636
rect 173340 112580 173396 112636
rect 173396 112580 173400 112636
rect 173336 112576 173400 112580
rect 173416 112636 173480 112640
rect 173416 112580 173420 112636
rect 173420 112580 173476 112636
rect 173476 112580 173480 112636
rect 173416 112576 173480 112580
rect 4216 112092 4280 112096
rect 4216 112036 4220 112092
rect 4220 112036 4276 112092
rect 4276 112036 4280 112092
rect 4216 112032 4280 112036
rect 4296 112092 4360 112096
rect 4296 112036 4300 112092
rect 4300 112036 4356 112092
rect 4356 112036 4360 112092
rect 4296 112032 4360 112036
rect 4376 112092 4440 112096
rect 4376 112036 4380 112092
rect 4380 112036 4436 112092
rect 4436 112036 4440 112092
rect 4376 112032 4440 112036
rect 4456 112092 4520 112096
rect 4456 112036 4460 112092
rect 4460 112036 4516 112092
rect 4516 112036 4520 112092
rect 4456 112032 4520 112036
rect 34936 112092 35000 112096
rect 34936 112036 34940 112092
rect 34940 112036 34996 112092
rect 34996 112036 35000 112092
rect 34936 112032 35000 112036
rect 35016 112092 35080 112096
rect 35016 112036 35020 112092
rect 35020 112036 35076 112092
rect 35076 112036 35080 112092
rect 35016 112032 35080 112036
rect 35096 112092 35160 112096
rect 35096 112036 35100 112092
rect 35100 112036 35156 112092
rect 35156 112036 35160 112092
rect 35096 112032 35160 112036
rect 35176 112092 35240 112096
rect 35176 112036 35180 112092
rect 35180 112036 35236 112092
rect 35236 112036 35240 112092
rect 35176 112032 35240 112036
rect 65656 112092 65720 112096
rect 65656 112036 65660 112092
rect 65660 112036 65716 112092
rect 65716 112036 65720 112092
rect 65656 112032 65720 112036
rect 65736 112092 65800 112096
rect 65736 112036 65740 112092
rect 65740 112036 65796 112092
rect 65796 112036 65800 112092
rect 65736 112032 65800 112036
rect 65816 112092 65880 112096
rect 65816 112036 65820 112092
rect 65820 112036 65876 112092
rect 65876 112036 65880 112092
rect 65816 112032 65880 112036
rect 65896 112092 65960 112096
rect 65896 112036 65900 112092
rect 65900 112036 65956 112092
rect 65956 112036 65960 112092
rect 65896 112032 65960 112036
rect 96376 112092 96440 112096
rect 96376 112036 96380 112092
rect 96380 112036 96436 112092
rect 96436 112036 96440 112092
rect 96376 112032 96440 112036
rect 96456 112092 96520 112096
rect 96456 112036 96460 112092
rect 96460 112036 96516 112092
rect 96516 112036 96520 112092
rect 96456 112032 96520 112036
rect 96536 112092 96600 112096
rect 96536 112036 96540 112092
rect 96540 112036 96596 112092
rect 96596 112036 96600 112092
rect 96536 112032 96600 112036
rect 96616 112092 96680 112096
rect 96616 112036 96620 112092
rect 96620 112036 96676 112092
rect 96676 112036 96680 112092
rect 96616 112032 96680 112036
rect 127096 112092 127160 112096
rect 127096 112036 127100 112092
rect 127100 112036 127156 112092
rect 127156 112036 127160 112092
rect 127096 112032 127160 112036
rect 127176 112092 127240 112096
rect 127176 112036 127180 112092
rect 127180 112036 127236 112092
rect 127236 112036 127240 112092
rect 127176 112032 127240 112036
rect 127256 112092 127320 112096
rect 127256 112036 127260 112092
rect 127260 112036 127316 112092
rect 127316 112036 127320 112092
rect 127256 112032 127320 112036
rect 127336 112092 127400 112096
rect 127336 112036 127340 112092
rect 127340 112036 127396 112092
rect 127396 112036 127400 112092
rect 127336 112032 127400 112036
rect 157816 112092 157880 112096
rect 157816 112036 157820 112092
rect 157820 112036 157876 112092
rect 157876 112036 157880 112092
rect 157816 112032 157880 112036
rect 157896 112092 157960 112096
rect 157896 112036 157900 112092
rect 157900 112036 157956 112092
rect 157956 112036 157960 112092
rect 157896 112032 157960 112036
rect 157976 112092 158040 112096
rect 157976 112036 157980 112092
rect 157980 112036 158036 112092
rect 158036 112036 158040 112092
rect 157976 112032 158040 112036
rect 158056 112092 158120 112096
rect 158056 112036 158060 112092
rect 158060 112036 158116 112092
rect 158116 112036 158120 112092
rect 158056 112032 158120 112036
rect 19576 111548 19640 111552
rect 19576 111492 19580 111548
rect 19580 111492 19636 111548
rect 19636 111492 19640 111548
rect 19576 111488 19640 111492
rect 19656 111548 19720 111552
rect 19656 111492 19660 111548
rect 19660 111492 19716 111548
rect 19716 111492 19720 111548
rect 19656 111488 19720 111492
rect 19736 111548 19800 111552
rect 19736 111492 19740 111548
rect 19740 111492 19796 111548
rect 19796 111492 19800 111548
rect 19736 111488 19800 111492
rect 19816 111548 19880 111552
rect 19816 111492 19820 111548
rect 19820 111492 19876 111548
rect 19876 111492 19880 111548
rect 19816 111488 19880 111492
rect 50296 111548 50360 111552
rect 50296 111492 50300 111548
rect 50300 111492 50356 111548
rect 50356 111492 50360 111548
rect 50296 111488 50360 111492
rect 50376 111548 50440 111552
rect 50376 111492 50380 111548
rect 50380 111492 50436 111548
rect 50436 111492 50440 111548
rect 50376 111488 50440 111492
rect 50456 111548 50520 111552
rect 50456 111492 50460 111548
rect 50460 111492 50516 111548
rect 50516 111492 50520 111548
rect 50456 111488 50520 111492
rect 50536 111548 50600 111552
rect 50536 111492 50540 111548
rect 50540 111492 50596 111548
rect 50596 111492 50600 111548
rect 50536 111488 50600 111492
rect 81016 111548 81080 111552
rect 81016 111492 81020 111548
rect 81020 111492 81076 111548
rect 81076 111492 81080 111548
rect 81016 111488 81080 111492
rect 81096 111548 81160 111552
rect 81096 111492 81100 111548
rect 81100 111492 81156 111548
rect 81156 111492 81160 111548
rect 81096 111488 81160 111492
rect 81176 111548 81240 111552
rect 81176 111492 81180 111548
rect 81180 111492 81236 111548
rect 81236 111492 81240 111548
rect 81176 111488 81240 111492
rect 81256 111548 81320 111552
rect 81256 111492 81260 111548
rect 81260 111492 81316 111548
rect 81316 111492 81320 111548
rect 81256 111488 81320 111492
rect 111736 111548 111800 111552
rect 111736 111492 111740 111548
rect 111740 111492 111796 111548
rect 111796 111492 111800 111548
rect 111736 111488 111800 111492
rect 111816 111548 111880 111552
rect 111816 111492 111820 111548
rect 111820 111492 111876 111548
rect 111876 111492 111880 111548
rect 111816 111488 111880 111492
rect 111896 111548 111960 111552
rect 111896 111492 111900 111548
rect 111900 111492 111956 111548
rect 111956 111492 111960 111548
rect 111896 111488 111960 111492
rect 111976 111548 112040 111552
rect 111976 111492 111980 111548
rect 111980 111492 112036 111548
rect 112036 111492 112040 111548
rect 111976 111488 112040 111492
rect 142456 111548 142520 111552
rect 142456 111492 142460 111548
rect 142460 111492 142516 111548
rect 142516 111492 142520 111548
rect 142456 111488 142520 111492
rect 142536 111548 142600 111552
rect 142536 111492 142540 111548
rect 142540 111492 142596 111548
rect 142596 111492 142600 111548
rect 142536 111488 142600 111492
rect 142616 111548 142680 111552
rect 142616 111492 142620 111548
rect 142620 111492 142676 111548
rect 142676 111492 142680 111548
rect 142616 111488 142680 111492
rect 142696 111548 142760 111552
rect 142696 111492 142700 111548
rect 142700 111492 142756 111548
rect 142756 111492 142760 111548
rect 142696 111488 142760 111492
rect 173176 111548 173240 111552
rect 173176 111492 173180 111548
rect 173180 111492 173236 111548
rect 173236 111492 173240 111548
rect 173176 111488 173240 111492
rect 173256 111548 173320 111552
rect 173256 111492 173260 111548
rect 173260 111492 173316 111548
rect 173316 111492 173320 111548
rect 173256 111488 173320 111492
rect 173336 111548 173400 111552
rect 173336 111492 173340 111548
rect 173340 111492 173396 111548
rect 173396 111492 173400 111548
rect 173336 111488 173400 111492
rect 173416 111548 173480 111552
rect 173416 111492 173420 111548
rect 173420 111492 173476 111548
rect 173476 111492 173480 111548
rect 173416 111488 173480 111492
rect 4216 111004 4280 111008
rect 4216 110948 4220 111004
rect 4220 110948 4276 111004
rect 4276 110948 4280 111004
rect 4216 110944 4280 110948
rect 4296 111004 4360 111008
rect 4296 110948 4300 111004
rect 4300 110948 4356 111004
rect 4356 110948 4360 111004
rect 4296 110944 4360 110948
rect 4376 111004 4440 111008
rect 4376 110948 4380 111004
rect 4380 110948 4436 111004
rect 4436 110948 4440 111004
rect 4376 110944 4440 110948
rect 4456 111004 4520 111008
rect 4456 110948 4460 111004
rect 4460 110948 4516 111004
rect 4516 110948 4520 111004
rect 4456 110944 4520 110948
rect 34936 111004 35000 111008
rect 34936 110948 34940 111004
rect 34940 110948 34996 111004
rect 34996 110948 35000 111004
rect 34936 110944 35000 110948
rect 35016 111004 35080 111008
rect 35016 110948 35020 111004
rect 35020 110948 35076 111004
rect 35076 110948 35080 111004
rect 35016 110944 35080 110948
rect 35096 111004 35160 111008
rect 35096 110948 35100 111004
rect 35100 110948 35156 111004
rect 35156 110948 35160 111004
rect 35096 110944 35160 110948
rect 35176 111004 35240 111008
rect 35176 110948 35180 111004
rect 35180 110948 35236 111004
rect 35236 110948 35240 111004
rect 35176 110944 35240 110948
rect 65656 111004 65720 111008
rect 65656 110948 65660 111004
rect 65660 110948 65716 111004
rect 65716 110948 65720 111004
rect 65656 110944 65720 110948
rect 65736 111004 65800 111008
rect 65736 110948 65740 111004
rect 65740 110948 65796 111004
rect 65796 110948 65800 111004
rect 65736 110944 65800 110948
rect 65816 111004 65880 111008
rect 65816 110948 65820 111004
rect 65820 110948 65876 111004
rect 65876 110948 65880 111004
rect 65816 110944 65880 110948
rect 65896 111004 65960 111008
rect 65896 110948 65900 111004
rect 65900 110948 65956 111004
rect 65956 110948 65960 111004
rect 65896 110944 65960 110948
rect 96376 111004 96440 111008
rect 96376 110948 96380 111004
rect 96380 110948 96436 111004
rect 96436 110948 96440 111004
rect 96376 110944 96440 110948
rect 96456 111004 96520 111008
rect 96456 110948 96460 111004
rect 96460 110948 96516 111004
rect 96516 110948 96520 111004
rect 96456 110944 96520 110948
rect 96536 111004 96600 111008
rect 96536 110948 96540 111004
rect 96540 110948 96596 111004
rect 96596 110948 96600 111004
rect 96536 110944 96600 110948
rect 96616 111004 96680 111008
rect 96616 110948 96620 111004
rect 96620 110948 96676 111004
rect 96676 110948 96680 111004
rect 96616 110944 96680 110948
rect 127096 111004 127160 111008
rect 127096 110948 127100 111004
rect 127100 110948 127156 111004
rect 127156 110948 127160 111004
rect 127096 110944 127160 110948
rect 127176 111004 127240 111008
rect 127176 110948 127180 111004
rect 127180 110948 127236 111004
rect 127236 110948 127240 111004
rect 127176 110944 127240 110948
rect 127256 111004 127320 111008
rect 127256 110948 127260 111004
rect 127260 110948 127316 111004
rect 127316 110948 127320 111004
rect 127256 110944 127320 110948
rect 127336 111004 127400 111008
rect 127336 110948 127340 111004
rect 127340 110948 127396 111004
rect 127396 110948 127400 111004
rect 127336 110944 127400 110948
rect 157816 111004 157880 111008
rect 157816 110948 157820 111004
rect 157820 110948 157876 111004
rect 157876 110948 157880 111004
rect 157816 110944 157880 110948
rect 157896 111004 157960 111008
rect 157896 110948 157900 111004
rect 157900 110948 157956 111004
rect 157956 110948 157960 111004
rect 157896 110944 157960 110948
rect 157976 111004 158040 111008
rect 157976 110948 157980 111004
rect 157980 110948 158036 111004
rect 158036 110948 158040 111004
rect 157976 110944 158040 110948
rect 158056 111004 158120 111008
rect 158056 110948 158060 111004
rect 158060 110948 158116 111004
rect 158116 110948 158120 111004
rect 158056 110944 158120 110948
rect 19576 110460 19640 110464
rect 19576 110404 19580 110460
rect 19580 110404 19636 110460
rect 19636 110404 19640 110460
rect 19576 110400 19640 110404
rect 19656 110460 19720 110464
rect 19656 110404 19660 110460
rect 19660 110404 19716 110460
rect 19716 110404 19720 110460
rect 19656 110400 19720 110404
rect 19736 110460 19800 110464
rect 19736 110404 19740 110460
rect 19740 110404 19796 110460
rect 19796 110404 19800 110460
rect 19736 110400 19800 110404
rect 19816 110460 19880 110464
rect 19816 110404 19820 110460
rect 19820 110404 19876 110460
rect 19876 110404 19880 110460
rect 19816 110400 19880 110404
rect 50296 110460 50360 110464
rect 50296 110404 50300 110460
rect 50300 110404 50356 110460
rect 50356 110404 50360 110460
rect 50296 110400 50360 110404
rect 50376 110460 50440 110464
rect 50376 110404 50380 110460
rect 50380 110404 50436 110460
rect 50436 110404 50440 110460
rect 50376 110400 50440 110404
rect 50456 110460 50520 110464
rect 50456 110404 50460 110460
rect 50460 110404 50516 110460
rect 50516 110404 50520 110460
rect 50456 110400 50520 110404
rect 50536 110460 50600 110464
rect 50536 110404 50540 110460
rect 50540 110404 50596 110460
rect 50596 110404 50600 110460
rect 50536 110400 50600 110404
rect 81016 110460 81080 110464
rect 81016 110404 81020 110460
rect 81020 110404 81076 110460
rect 81076 110404 81080 110460
rect 81016 110400 81080 110404
rect 81096 110460 81160 110464
rect 81096 110404 81100 110460
rect 81100 110404 81156 110460
rect 81156 110404 81160 110460
rect 81096 110400 81160 110404
rect 81176 110460 81240 110464
rect 81176 110404 81180 110460
rect 81180 110404 81236 110460
rect 81236 110404 81240 110460
rect 81176 110400 81240 110404
rect 81256 110460 81320 110464
rect 81256 110404 81260 110460
rect 81260 110404 81316 110460
rect 81316 110404 81320 110460
rect 81256 110400 81320 110404
rect 111736 110460 111800 110464
rect 111736 110404 111740 110460
rect 111740 110404 111796 110460
rect 111796 110404 111800 110460
rect 111736 110400 111800 110404
rect 111816 110460 111880 110464
rect 111816 110404 111820 110460
rect 111820 110404 111876 110460
rect 111876 110404 111880 110460
rect 111816 110400 111880 110404
rect 111896 110460 111960 110464
rect 111896 110404 111900 110460
rect 111900 110404 111956 110460
rect 111956 110404 111960 110460
rect 111896 110400 111960 110404
rect 111976 110460 112040 110464
rect 111976 110404 111980 110460
rect 111980 110404 112036 110460
rect 112036 110404 112040 110460
rect 111976 110400 112040 110404
rect 142456 110460 142520 110464
rect 142456 110404 142460 110460
rect 142460 110404 142516 110460
rect 142516 110404 142520 110460
rect 142456 110400 142520 110404
rect 142536 110460 142600 110464
rect 142536 110404 142540 110460
rect 142540 110404 142596 110460
rect 142596 110404 142600 110460
rect 142536 110400 142600 110404
rect 142616 110460 142680 110464
rect 142616 110404 142620 110460
rect 142620 110404 142676 110460
rect 142676 110404 142680 110460
rect 142616 110400 142680 110404
rect 142696 110460 142760 110464
rect 142696 110404 142700 110460
rect 142700 110404 142756 110460
rect 142756 110404 142760 110460
rect 142696 110400 142760 110404
rect 173176 110460 173240 110464
rect 173176 110404 173180 110460
rect 173180 110404 173236 110460
rect 173236 110404 173240 110460
rect 173176 110400 173240 110404
rect 173256 110460 173320 110464
rect 173256 110404 173260 110460
rect 173260 110404 173316 110460
rect 173316 110404 173320 110460
rect 173256 110400 173320 110404
rect 173336 110460 173400 110464
rect 173336 110404 173340 110460
rect 173340 110404 173396 110460
rect 173396 110404 173400 110460
rect 173336 110400 173400 110404
rect 173416 110460 173480 110464
rect 173416 110404 173420 110460
rect 173420 110404 173476 110460
rect 173476 110404 173480 110460
rect 173416 110400 173480 110404
rect 4216 109916 4280 109920
rect 4216 109860 4220 109916
rect 4220 109860 4276 109916
rect 4276 109860 4280 109916
rect 4216 109856 4280 109860
rect 4296 109916 4360 109920
rect 4296 109860 4300 109916
rect 4300 109860 4356 109916
rect 4356 109860 4360 109916
rect 4296 109856 4360 109860
rect 4376 109916 4440 109920
rect 4376 109860 4380 109916
rect 4380 109860 4436 109916
rect 4436 109860 4440 109916
rect 4376 109856 4440 109860
rect 4456 109916 4520 109920
rect 4456 109860 4460 109916
rect 4460 109860 4516 109916
rect 4516 109860 4520 109916
rect 4456 109856 4520 109860
rect 34936 109916 35000 109920
rect 34936 109860 34940 109916
rect 34940 109860 34996 109916
rect 34996 109860 35000 109916
rect 34936 109856 35000 109860
rect 35016 109916 35080 109920
rect 35016 109860 35020 109916
rect 35020 109860 35076 109916
rect 35076 109860 35080 109916
rect 35016 109856 35080 109860
rect 35096 109916 35160 109920
rect 35096 109860 35100 109916
rect 35100 109860 35156 109916
rect 35156 109860 35160 109916
rect 35096 109856 35160 109860
rect 35176 109916 35240 109920
rect 35176 109860 35180 109916
rect 35180 109860 35236 109916
rect 35236 109860 35240 109916
rect 35176 109856 35240 109860
rect 65656 109916 65720 109920
rect 65656 109860 65660 109916
rect 65660 109860 65716 109916
rect 65716 109860 65720 109916
rect 65656 109856 65720 109860
rect 65736 109916 65800 109920
rect 65736 109860 65740 109916
rect 65740 109860 65796 109916
rect 65796 109860 65800 109916
rect 65736 109856 65800 109860
rect 65816 109916 65880 109920
rect 65816 109860 65820 109916
rect 65820 109860 65876 109916
rect 65876 109860 65880 109916
rect 65816 109856 65880 109860
rect 65896 109916 65960 109920
rect 65896 109860 65900 109916
rect 65900 109860 65956 109916
rect 65956 109860 65960 109916
rect 65896 109856 65960 109860
rect 96376 109916 96440 109920
rect 96376 109860 96380 109916
rect 96380 109860 96436 109916
rect 96436 109860 96440 109916
rect 96376 109856 96440 109860
rect 96456 109916 96520 109920
rect 96456 109860 96460 109916
rect 96460 109860 96516 109916
rect 96516 109860 96520 109916
rect 96456 109856 96520 109860
rect 96536 109916 96600 109920
rect 96536 109860 96540 109916
rect 96540 109860 96596 109916
rect 96596 109860 96600 109916
rect 96536 109856 96600 109860
rect 96616 109916 96680 109920
rect 96616 109860 96620 109916
rect 96620 109860 96676 109916
rect 96676 109860 96680 109916
rect 96616 109856 96680 109860
rect 127096 109916 127160 109920
rect 127096 109860 127100 109916
rect 127100 109860 127156 109916
rect 127156 109860 127160 109916
rect 127096 109856 127160 109860
rect 127176 109916 127240 109920
rect 127176 109860 127180 109916
rect 127180 109860 127236 109916
rect 127236 109860 127240 109916
rect 127176 109856 127240 109860
rect 127256 109916 127320 109920
rect 127256 109860 127260 109916
rect 127260 109860 127316 109916
rect 127316 109860 127320 109916
rect 127256 109856 127320 109860
rect 127336 109916 127400 109920
rect 127336 109860 127340 109916
rect 127340 109860 127396 109916
rect 127396 109860 127400 109916
rect 127336 109856 127400 109860
rect 157816 109916 157880 109920
rect 157816 109860 157820 109916
rect 157820 109860 157876 109916
rect 157876 109860 157880 109916
rect 157816 109856 157880 109860
rect 157896 109916 157960 109920
rect 157896 109860 157900 109916
rect 157900 109860 157956 109916
rect 157956 109860 157960 109916
rect 157896 109856 157960 109860
rect 157976 109916 158040 109920
rect 157976 109860 157980 109916
rect 157980 109860 158036 109916
rect 158036 109860 158040 109916
rect 157976 109856 158040 109860
rect 158056 109916 158120 109920
rect 158056 109860 158060 109916
rect 158060 109860 158116 109916
rect 158116 109860 158120 109916
rect 158056 109856 158120 109860
rect 19576 109372 19640 109376
rect 19576 109316 19580 109372
rect 19580 109316 19636 109372
rect 19636 109316 19640 109372
rect 19576 109312 19640 109316
rect 19656 109372 19720 109376
rect 19656 109316 19660 109372
rect 19660 109316 19716 109372
rect 19716 109316 19720 109372
rect 19656 109312 19720 109316
rect 19736 109372 19800 109376
rect 19736 109316 19740 109372
rect 19740 109316 19796 109372
rect 19796 109316 19800 109372
rect 19736 109312 19800 109316
rect 19816 109372 19880 109376
rect 19816 109316 19820 109372
rect 19820 109316 19876 109372
rect 19876 109316 19880 109372
rect 19816 109312 19880 109316
rect 50296 109372 50360 109376
rect 50296 109316 50300 109372
rect 50300 109316 50356 109372
rect 50356 109316 50360 109372
rect 50296 109312 50360 109316
rect 50376 109372 50440 109376
rect 50376 109316 50380 109372
rect 50380 109316 50436 109372
rect 50436 109316 50440 109372
rect 50376 109312 50440 109316
rect 50456 109372 50520 109376
rect 50456 109316 50460 109372
rect 50460 109316 50516 109372
rect 50516 109316 50520 109372
rect 50456 109312 50520 109316
rect 50536 109372 50600 109376
rect 50536 109316 50540 109372
rect 50540 109316 50596 109372
rect 50596 109316 50600 109372
rect 50536 109312 50600 109316
rect 81016 109372 81080 109376
rect 81016 109316 81020 109372
rect 81020 109316 81076 109372
rect 81076 109316 81080 109372
rect 81016 109312 81080 109316
rect 81096 109372 81160 109376
rect 81096 109316 81100 109372
rect 81100 109316 81156 109372
rect 81156 109316 81160 109372
rect 81096 109312 81160 109316
rect 81176 109372 81240 109376
rect 81176 109316 81180 109372
rect 81180 109316 81236 109372
rect 81236 109316 81240 109372
rect 81176 109312 81240 109316
rect 81256 109372 81320 109376
rect 81256 109316 81260 109372
rect 81260 109316 81316 109372
rect 81316 109316 81320 109372
rect 81256 109312 81320 109316
rect 111736 109372 111800 109376
rect 111736 109316 111740 109372
rect 111740 109316 111796 109372
rect 111796 109316 111800 109372
rect 111736 109312 111800 109316
rect 111816 109372 111880 109376
rect 111816 109316 111820 109372
rect 111820 109316 111876 109372
rect 111876 109316 111880 109372
rect 111816 109312 111880 109316
rect 111896 109372 111960 109376
rect 111896 109316 111900 109372
rect 111900 109316 111956 109372
rect 111956 109316 111960 109372
rect 111896 109312 111960 109316
rect 111976 109372 112040 109376
rect 111976 109316 111980 109372
rect 111980 109316 112036 109372
rect 112036 109316 112040 109372
rect 111976 109312 112040 109316
rect 142456 109372 142520 109376
rect 142456 109316 142460 109372
rect 142460 109316 142516 109372
rect 142516 109316 142520 109372
rect 142456 109312 142520 109316
rect 142536 109372 142600 109376
rect 142536 109316 142540 109372
rect 142540 109316 142596 109372
rect 142596 109316 142600 109372
rect 142536 109312 142600 109316
rect 142616 109372 142680 109376
rect 142616 109316 142620 109372
rect 142620 109316 142676 109372
rect 142676 109316 142680 109372
rect 142616 109312 142680 109316
rect 142696 109372 142760 109376
rect 142696 109316 142700 109372
rect 142700 109316 142756 109372
rect 142756 109316 142760 109372
rect 142696 109312 142760 109316
rect 173176 109372 173240 109376
rect 173176 109316 173180 109372
rect 173180 109316 173236 109372
rect 173236 109316 173240 109372
rect 173176 109312 173240 109316
rect 173256 109372 173320 109376
rect 173256 109316 173260 109372
rect 173260 109316 173316 109372
rect 173316 109316 173320 109372
rect 173256 109312 173320 109316
rect 173336 109372 173400 109376
rect 173336 109316 173340 109372
rect 173340 109316 173396 109372
rect 173396 109316 173400 109372
rect 173336 109312 173400 109316
rect 173416 109372 173480 109376
rect 173416 109316 173420 109372
rect 173420 109316 173476 109372
rect 173476 109316 173480 109372
rect 173416 109312 173480 109316
rect 4216 108828 4280 108832
rect 4216 108772 4220 108828
rect 4220 108772 4276 108828
rect 4276 108772 4280 108828
rect 4216 108768 4280 108772
rect 4296 108828 4360 108832
rect 4296 108772 4300 108828
rect 4300 108772 4356 108828
rect 4356 108772 4360 108828
rect 4296 108768 4360 108772
rect 4376 108828 4440 108832
rect 4376 108772 4380 108828
rect 4380 108772 4436 108828
rect 4436 108772 4440 108828
rect 4376 108768 4440 108772
rect 4456 108828 4520 108832
rect 4456 108772 4460 108828
rect 4460 108772 4516 108828
rect 4516 108772 4520 108828
rect 4456 108768 4520 108772
rect 34936 108828 35000 108832
rect 34936 108772 34940 108828
rect 34940 108772 34996 108828
rect 34996 108772 35000 108828
rect 34936 108768 35000 108772
rect 35016 108828 35080 108832
rect 35016 108772 35020 108828
rect 35020 108772 35076 108828
rect 35076 108772 35080 108828
rect 35016 108768 35080 108772
rect 35096 108828 35160 108832
rect 35096 108772 35100 108828
rect 35100 108772 35156 108828
rect 35156 108772 35160 108828
rect 35096 108768 35160 108772
rect 35176 108828 35240 108832
rect 35176 108772 35180 108828
rect 35180 108772 35236 108828
rect 35236 108772 35240 108828
rect 35176 108768 35240 108772
rect 65656 108828 65720 108832
rect 65656 108772 65660 108828
rect 65660 108772 65716 108828
rect 65716 108772 65720 108828
rect 65656 108768 65720 108772
rect 65736 108828 65800 108832
rect 65736 108772 65740 108828
rect 65740 108772 65796 108828
rect 65796 108772 65800 108828
rect 65736 108768 65800 108772
rect 65816 108828 65880 108832
rect 65816 108772 65820 108828
rect 65820 108772 65876 108828
rect 65876 108772 65880 108828
rect 65816 108768 65880 108772
rect 65896 108828 65960 108832
rect 65896 108772 65900 108828
rect 65900 108772 65956 108828
rect 65956 108772 65960 108828
rect 65896 108768 65960 108772
rect 96376 108828 96440 108832
rect 96376 108772 96380 108828
rect 96380 108772 96436 108828
rect 96436 108772 96440 108828
rect 96376 108768 96440 108772
rect 96456 108828 96520 108832
rect 96456 108772 96460 108828
rect 96460 108772 96516 108828
rect 96516 108772 96520 108828
rect 96456 108768 96520 108772
rect 96536 108828 96600 108832
rect 96536 108772 96540 108828
rect 96540 108772 96596 108828
rect 96596 108772 96600 108828
rect 96536 108768 96600 108772
rect 96616 108828 96680 108832
rect 96616 108772 96620 108828
rect 96620 108772 96676 108828
rect 96676 108772 96680 108828
rect 96616 108768 96680 108772
rect 127096 108828 127160 108832
rect 127096 108772 127100 108828
rect 127100 108772 127156 108828
rect 127156 108772 127160 108828
rect 127096 108768 127160 108772
rect 127176 108828 127240 108832
rect 127176 108772 127180 108828
rect 127180 108772 127236 108828
rect 127236 108772 127240 108828
rect 127176 108768 127240 108772
rect 127256 108828 127320 108832
rect 127256 108772 127260 108828
rect 127260 108772 127316 108828
rect 127316 108772 127320 108828
rect 127256 108768 127320 108772
rect 127336 108828 127400 108832
rect 127336 108772 127340 108828
rect 127340 108772 127396 108828
rect 127396 108772 127400 108828
rect 127336 108768 127400 108772
rect 157816 108828 157880 108832
rect 157816 108772 157820 108828
rect 157820 108772 157876 108828
rect 157876 108772 157880 108828
rect 157816 108768 157880 108772
rect 157896 108828 157960 108832
rect 157896 108772 157900 108828
rect 157900 108772 157956 108828
rect 157956 108772 157960 108828
rect 157896 108768 157960 108772
rect 157976 108828 158040 108832
rect 157976 108772 157980 108828
rect 157980 108772 158036 108828
rect 158036 108772 158040 108828
rect 157976 108768 158040 108772
rect 158056 108828 158120 108832
rect 158056 108772 158060 108828
rect 158060 108772 158116 108828
rect 158116 108772 158120 108828
rect 158056 108768 158120 108772
rect 19576 108284 19640 108288
rect 19576 108228 19580 108284
rect 19580 108228 19636 108284
rect 19636 108228 19640 108284
rect 19576 108224 19640 108228
rect 19656 108284 19720 108288
rect 19656 108228 19660 108284
rect 19660 108228 19716 108284
rect 19716 108228 19720 108284
rect 19656 108224 19720 108228
rect 19736 108284 19800 108288
rect 19736 108228 19740 108284
rect 19740 108228 19796 108284
rect 19796 108228 19800 108284
rect 19736 108224 19800 108228
rect 19816 108284 19880 108288
rect 19816 108228 19820 108284
rect 19820 108228 19876 108284
rect 19876 108228 19880 108284
rect 19816 108224 19880 108228
rect 50296 108284 50360 108288
rect 50296 108228 50300 108284
rect 50300 108228 50356 108284
rect 50356 108228 50360 108284
rect 50296 108224 50360 108228
rect 50376 108284 50440 108288
rect 50376 108228 50380 108284
rect 50380 108228 50436 108284
rect 50436 108228 50440 108284
rect 50376 108224 50440 108228
rect 50456 108284 50520 108288
rect 50456 108228 50460 108284
rect 50460 108228 50516 108284
rect 50516 108228 50520 108284
rect 50456 108224 50520 108228
rect 50536 108284 50600 108288
rect 50536 108228 50540 108284
rect 50540 108228 50596 108284
rect 50596 108228 50600 108284
rect 50536 108224 50600 108228
rect 81016 108284 81080 108288
rect 81016 108228 81020 108284
rect 81020 108228 81076 108284
rect 81076 108228 81080 108284
rect 81016 108224 81080 108228
rect 81096 108284 81160 108288
rect 81096 108228 81100 108284
rect 81100 108228 81156 108284
rect 81156 108228 81160 108284
rect 81096 108224 81160 108228
rect 81176 108284 81240 108288
rect 81176 108228 81180 108284
rect 81180 108228 81236 108284
rect 81236 108228 81240 108284
rect 81176 108224 81240 108228
rect 81256 108284 81320 108288
rect 81256 108228 81260 108284
rect 81260 108228 81316 108284
rect 81316 108228 81320 108284
rect 81256 108224 81320 108228
rect 111736 108284 111800 108288
rect 111736 108228 111740 108284
rect 111740 108228 111796 108284
rect 111796 108228 111800 108284
rect 111736 108224 111800 108228
rect 111816 108284 111880 108288
rect 111816 108228 111820 108284
rect 111820 108228 111876 108284
rect 111876 108228 111880 108284
rect 111816 108224 111880 108228
rect 111896 108284 111960 108288
rect 111896 108228 111900 108284
rect 111900 108228 111956 108284
rect 111956 108228 111960 108284
rect 111896 108224 111960 108228
rect 111976 108284 112040 108288
rect 111976 108228 111980 108284
rect 111980 108228 112036 108284
rect 112036 108228 112040 108284
rect 111976 108224 112040 108228
rect 142456 108284 142520 108288
rect 142456 108228 142460 108284
rect 142460 108228 142516 108284
rect 142516 108228 142520 108284
rect 142456 108224 142520 108228
rect 142536 108284 142600 108288
rect 142536 108228 142540 108284
rect 142540 108228 142596 108284
rect 142596 108228 142600 108284
rect 142536 108224 142600 108228
rect 142616 108284 142680 108288
rect 142616 108228 142620 108284
rect 142620 108228 142676 108284
rect 142676 108228 142680 108284
rect 142616 108224 142680 108228
rect 142696 108284 142760 108288
rect 142696 108228 142700 108284
rect 142700 108228 142756 108284
rect 142756 108228 142760 108284
rect 142696 108224 142760 108228
rect 173176 108284 173240 108288
rect 173176 108228 173180 108284
rect 173180 108228 173236 108284
rect 173236 108228 173240 108284
rect 173176 108224 173240 108228
rect 173256 108284 173320 108288
rect 173256 108228 173260 108284
rect 173260 108228 173316 108284
rect 173316 108228 173320 108284
rect 173256 108224 173320 108228
rect 173336 108284 173400 108288
rect 173336 108228 173340 108284
rect 173340 108228 173396 108284
rect 173396 108228 173400 108284
rect 173336 108224 173400 108228
rect 173416 108284 173480 108288
rect 173416 108228 173420 108284
rect 173420 108228 173476 108284
rect 173476 108228 173480 108284
rect 173416 108224 173480 108228
rect 4216 107740 4280 107744
rect 4216 107684 4220 107740
rect 4220 107684 4276 107740
rect 4276 107684 4280 107740
rect 4216 107680 4280 107684
rect 4296 107740 4360 107744
rect 4296 107684 4300 107740
rect 4300 107684 4356 107740
rect 4356 107684 4360 107740
rect 4296 107680 4360 107684
rect 4376 107740 4440 107744
rect 4376 107684 4380 107740
rect 4380 107684 4436 107740
rect 4436 107684 4440 107740
rect 4376 107680 4440 107684
rect 4456 107740 4520 107744
rect 4456 107684 4460 107740
rect 4460 107684 4516 107740
rect 4516 107684 4520 107740
rect 4456 107680 4520 107684
rect 34936 107740 35000 107744
rect 34936 107684 34940 107740
rect 34940 107684 34996 107740
rect 34996 107684 35000 107740
rect 34936 107680 35000 107684
rect 35016 107740 35080 107744
rect 35016 107684 35020 107740
rect 35020 107684 35076 107740
rect 35076 107684 35080 107740
rect 35016 107680 35080 107684
rect 35096 107740 35160 107744
rect 35096 107684 35100 107740
rect 35100 107684 35156 107740
rect 35156 107684 35160 107740
rect 35096 107680 35160 107684
rect 35176 107740 35240 107744
rect 35176 107684 35180 107740
rect 35180 107684 35236 107740
rect 35236 107684 35240 107740
rect 35176 107680 35240 107684
rect 65656 107740 65720 107744
rect 65656 107684 65660 107740
rect 65660 107684 65716 107740
rect 65716 107684 65720 107740
rect 65656 107680 65720 107684
rect 65736 107740 65800 107744
rect 65736 107684 65740 107740
rect 65740 107684 65796 107740
rect 65796 107684 65800 107740
rect 65736 107680 65800 107684
rect 65816 107740 65880 107744
rect 65816 107684 65820 107740
rect 65820 107684 65876 107740
rect 65876 107684 65880 107740
rect 65816 107680 65880 107684
rect 65896 107740 65960 107744
rect 65896 107684 65900 107740
rect 65900 107684 65956 107740
rect 65956 107684 65960 107740
rect 65896 107680 65960 107684
rect 96376 107740 96440 107744
rect 96376 107684 96380 107740
rect 96380 107684 96436 107740
rect 96436 107684 96440 107740
rect 96376 107680 96440 107684
rect 96456 107740 96520 107744
rect 96456 107684 96460 107740
rect 96460 107684 96516 107740
rect 96516 107684 96520 107740
rect 96456 107680 96520 107684
rect 96536 107740 96600 107744
rect 96536 107684 96540 107740
rect 96540 107684 96596 107740
rect 96596 107684 96600 107740
rect 96536 107680 96600 107684
rect 96616 107740 96680 107744
rect 96616 107684 96620 107740
rect 96620 107684 96676 107740
rect 96676 107684 96680 107740
rect 96616 107680 96680 107684
rect 127096 107740 127160 107744
rect 127096 107684 127100 107740
rect 127100 107684 127156 107740
rect 127156 107684 127160 107740
rect 127096 107680 127160 107684
rect 127176 107740 127240 107744
rect 127176 107684 127180 107740
rect 127180 107684 127236 107740
rect 127236 107684 127240 107740
rect 127176 107680 127240 107684
rect 127256 107740 127320 107744
rect 127256 107684 127260 107740
rect 127260 107684 127316 107740
rect 127316 107684 127320 107740
rect 127256 107680 127320 107684
rect 127336 107740 127400 107744
rect 127336 107684 127340 107740
rect 127340 107684 127396 107740
rect 127396 107684 127400 107740
rect 127336 107680 127400 107684
rect 157816 107740 157880 107744
rect 157816 107684 157820 107740
rect 157820 107684 157876 107740
rect 157876 107684 157880 107740
rect 157816 107680 157880 107684
rect 157896 107740 157960 107744
rect 157896 107684 157900 107740
rect 157900 107684 157956 107740
rect 157956 107684 157960 107740
rect 157896 107680 157960 107684
rect 157976 107740 158040 107744
rect 157976 107684 157980 107740
rect 157980 107684 158036 107740
rect 158036 107684 158040 107740
rect 157976 107680 158040 107684
rect 158056 107740 158120 107744
rect 158056 107684 158060 107740
rect 158060 107684 158116 107740
rect 158116 107684 158120 107740
rect 158056 107680 158120 107684
rect 19576 107196 19640 107200
rect 19576 107140 19580 107196
rect 19580 107140 19636 107196
rect 19636 107140 19640 107196
rect 19576 107136 19640 107140
rect 19656 107196 19720 107200
rect 19656 107140 19660 107196
rect 19660 107140 19716 107196
rect 19716 107140 19720 107196
rect 19656 107136 19720 107140
rect 19736 107196 19800 107200
rect 19736 107140 19740 107196
rect 19740 107140 19796 107196
rect 19796 107140 19800 107196
rect 19736 107136 19800 107140
rect 19816 107196 19880 107200
rect 19816 107140 19820 107196
rect 19820 107140 19876 107196
rect 19876 107140 19880 107196
rect 19816 107136 19880 107140
rect 50296 107196 50360 107200
rect 50296 107140 50300 107196
rect 50300 107140 50356 107196
rect 50356 107140 50360 107196
rect 50296 107136 50360 107140
rect 50376 107196 50440 107200
rect 50376 107140 50380 107196
rect 50380 107140 50436 107196
rect 50436 107140 50440 107196
rect 50376 107136 50440 107140
rect 50456 107196 50520 107200
rect 50456 107140 50460 107196
rect 50460 107140 50516 107196
rect 50516 107140 50520 107196
rect 50456 107136 50520 107140
rect 50536 107196 50600 107200
rect 50536 107140 50540 107196
rect 50540 107140 50596 107196
rect 50596 107140 50600 107196
rect 50536 107136 50600 107140
rect 81016 107196 81080 107200
rect 81016 107140 81020 107196
rect 81020 107140 81076 107196
rect 81076 107140 81080 107196
rect 81016 107136 81080 107140
rect 81096 107196 81160 107200
rect 81096 107140 81100 107196
rect 81100 107140 81156 107196
rect 81156 107140 81160 107196
rect 81096 107136 81160 107140
rect 81176 107196 81240 107200
rect 81176 107140 81180 107196
rect 81180 107140 81236 107196
rect 81236 107140 81240 107196
rect 81176 107136 81240 107140
rect 81256 107196 81320 107200
rect 81256 107140 81260 107196
rect 81260 107140 81316 107196
rect 81316 107140 81320 107196
rect 81256 107136 81320 107140
rect 111736 107196 111800 107200
rect 111736 107140 111740 107196
rect 111740 107140 111796 107196
rect 111796 107140 111800 107196
rect 111736 107136 111800 107140
rect 111816 107196 111880 107200
rect 111816 107140 111820 107196
rect 111820 107140 111876 107196
rect 111876 107140 111880 107196
rect 111816 107136 111880 107140
rect 111896 107196 111960 107200
rect 111896 107140 111900 107196
rect 111900 107140 111956 107196
rect 111956 107140 111960 107196
rect 111896 107136 111960 107140
rect 111976 107196 112040 107200
rect 111976 107140 111980 107196
rect 111980 107140 112036 107196
rect 112036 107140 112040 107196
rect 111976 107136 112040 107140
rect 142456 107196 142520 107200
rect 142456 107140 142460 107196
rect 142460 107140 142516 107196
rect 142516 107140 142520 107196
rect 142456 107136 142520 107140
rect 142536 107196 142600 107200
rect 142536 107140 142540 107196
rect 142540 107140 142596 107196
rect 142596 107140 142600 107196
rect 142536 107136 142600 107140
rect 142616 107196 142680 107200
rect 142616 107140 142620 107196
rect 142620 107140 142676 107196
rect 142676 107140 142680 107196
rect 142616 107136 142680 107140
rect 142696 107196 142760 107200
rect 142696 107140 142700 107196
rect 142700 107140 142756 107196
rect 142756 107140 142760 107196
rect 142696 107136 142760 107140
rect 173176 107196 173240 107200
rect 173176 107140 173180 107196
rect 173180 107140 173236 107196
rect 173236 107140 173240 107196
rect 173176 107136 173240 107140
rect 173256 107196 173320 107200
rect 173256 107140 173260 107196
rect 173260 107140 173316 107196
rect 173316 107140 173320 107196
rect 173256 107136 173320 107140
rect 173336 107196 173400 107200
rect 173336 107140 173340 107196
rect 173340 107140 173396 107196
rect 173396 107140 173400 107196
rect 173336 107136 173400 107140
rect 173416 107196 173480 107200
rect 173416 107140 173420 107196
rect 173420 107140 173476 107196
rect 173476 107140 173480 107196
rect 173416 107136 173480 107140
rect 4216 106652 4280 106656
rect 4216 106596 4220 106652
rect 4220 106596 4276 106652
rect 4276 106596 4280 106652
rect 4216 106592 4280 106596
rect 4296 106652 4360 106656
rect 4296 106596 4300 106652
rect 4300 106596 4356 106652
rect 4356 106596 4360 106652
rect 4296 106592 4360 106596
rect 4376 106652 4440 106656
rect 4376 106596 4380 106652
rect 4380 106596 4436 106652
rect 4436 106596 4440 106652
rect 4376 106592 4440 106596
rect 4456 106652 4520 106656
rect 4456 106596 4460 106652
rect 4460 106596 4516 106652
rect 4516 106596 4520 106652
rect 4456 106592 4520 106596
rect 34936 106652 35000 106656
rect 34936 106596 34940 106652
rect 34940 106596 34996 106652
rect 34996 106596 35000 106652
rect 34936 106592 35000 106596
rect 35016 106652 35080 106656
rect 35016 106596 35020 106652
rect 35020 106596 35076 106652
rect 35076 106596 35080 106652
rect 35016 106592 35080 106596
rect 35096 106652 35160 106656
rect 35096 106596 35100 106652
rect 35100 106596 35156 106652
rect 35156 106596 35160 106652
rect 35096 106592 35160 106596
rect 35176 106652 35240 106656
rect 35176 106596 35180 106652
rect 35180 106596 35236 106652
rect 35236 106596 35240 106652
rect 35176 106592 35240 106596
rect 65656 106652 65720 106656
rect 65656 106596 65660 106652
rect 65660 106596 65716 106652
rect 65716 106596 65720 106652
rect 65656 106592 65720 106596
rect 65736 106652 65800 106656
rect 65736 106596 65740 106652
rect 65740 106596 65796 106652
rect 65796 106596 65800 106652
rect 65736 106592 65800 106596
rect 65816 106652 65880 106656
rect 65816 106596 65820 106652
rect 65820 106596 65876 106652
rect 65876 106596 65880 106652
rect 65816 106592 65880 106596
rect 65896 106652 65960 106656
rect 65896 106596 65900 106652
rect 65900 106596 65956 106652
rect 65956 106596 65960 106652
rect 65896 106592 65960 106596
rect 96376 106652 96440 106656
rect 96376 106596 96380 106652
rect 96380 106596 96436 106652
rect 96436 106596 96440 106652
rect 96376 106592 96440 106596
rect 96456 106652 96520 106656
rect 96456 106596 96460 106652
rect 96460 106596 96516 106652
rect 96516 106596 96520 106652
rect 96456 106592 96520 106596
rect 96536 106652 96600 106656
rect 96536 106596 96540 106652
rect 96540 106596 96596 106652
rect 96596 106596 96600 106652
rect 96536 106592 96600 106596
rect 96616 106652 96680 106656
rect 96616 106596 96620 106652
rect 96620 106596 96676 106652
rect 96676 106596 96680 106652
rect 96616 106592 96680 106596
rect 127096 106652 127160 106656
rect 127096 106596 127100 106652
rect 127100 106596 127156 106652
rect 127156 106596 127160 106652
rect 127096 106592 127160 106596
rect 127176 106652 127240 106656
rect 127176 106596 127180 106652
rect 127180 106596 127236 106652
rect 127236 106596 127240 106652
rect 127176 106592 127240 106596
rect 127256 106652 127320 106656
rect 127256 106596 127260 106652
rect 127260 106596 127316 106652
rect 127316 106596 127320 106652
rect 127256 106592 127320 106596
rect 127336 106652 127400 106656
rect 127336 106596 127340 106652
rect 127340 106596 127396 106652
rect 127396 106596 127400 106652
rect 127336 106592 127400 106596
rect 157816 106652 157880 106656
rect 157816 106596 157820 106652
rect 157820 106596 157876 106652
rect 157876 106596 157880 106652
rect 157816 106592 157880 106596
rect 157896 106652 157960 106656
rect 157896 106596 157900 106652
rect 157900 106596 157956 106652
rect 157956 106596 157960 106652
rect 157896 106592 157960 106596
rect 157976 106652 158040 106656
rect 157976 106596 157980 106652
rect 157980 106596 158036 106652
rect 158036 106596 158040 106652
rect 157976 106592 158040 106596
rect 158056 106652 158120 106656
rect 158056 106596 158060 106652
rect 158060 106596 158116 106652
rect 158116 106596 158120 106652
rect 158056 106592 158120 106596
rect 19576 106108 19640 106112
rect 19576 106052 19580 106108
rect 19580 106052 19636 106108
rect 19636 106052 19640 106108
rect 19576 106048 19640 106052
rect 19656 106108 19720 106112
rect 19656 106052 19660 106108
rect 19660 106052 19716 106108
rect 19716 106052 19720 106108
rect 19656 106048 19720 106052
rect 19736 106108 19800 106112
rect 19736 106052 19740 106108
rect 19740 106052 19796 106108
rect 19796 106052 19800 106108
rect 19736 106048 19800 106052
rect 19816 106108 19880 106112
rect 19816 106052 19820 106108
rect 19820 106052 19876 106108
rect 19876 106052 19880 106108
rect 19816 106048 19880 106052
rect 50296 106108 50360 106112
rect 50296 106052 50300 106108
rect 50300 106052 50356 106108
rect 50356 106052 50360 106108
rect 50296 106048 50360 106052
rect 50376 106108 50440 106112
rect 50376 106052 50380 106108
rect 50380 106052 50436 106108
rect 50436 106052 50440 106108
rect 50376 106048 50440 106052
rect 50456 106108 50520 106112
rect 50456 106052 50460 106108
rect 50460 106052 50516 106108
rect 50516 106052 50520 106108
rect 50456 106048 50520 106052
rect 50536 106108 50600 106112
rect 50536 106052 50540 106108
rect 50540 106052 50596 106108
rect 50596 106052 50600 106108
rect 50536 106048 50600 106052
rect 81016 106108 81080 106112
rect 81016 106052 81020 106108
rect 81020 106052 81076 106108
rect 81076 106052 81080 106108
rect 81016 106048 81080 106052
rect 81096 106108 81160 106112
rect 81096 106052 81100 106108
rect 81100 106052 81156 106108
rect 81156 106052 81160 106108
rect 81096 106048 81160 106052
rect 81176 106108 81240 106112
rect 81176 106052 81180 106108
rect 81180 106052 81236 106108
rect 81236 106052 81240 106108
rect 81176 106048 81240 106052
rect 81256 106108 81320 106112
rect 81256 106052 81260 106108
rect 81260 106052 81316 106108
rect 81316 106052 81320 106108
rect 81256 106048 81320 106052
rect 111736 106108 111800 106112
rect 111736 106052 111740 106108
rect 111740 106052 111796 106108
rect 111796 106052 111800 106108
rect 111736 106048 111800 106052
rect 111816 106108 111880 106112
rect 111816 106052 111820 106108
rect 111820 106052 111876 106108
rect 111876 106052 111880 106108
rect 111816 106048 111880 106052
rect 111896 106108 111960 106112
rect 111896 106052 111900 106108
rect 111900 106052 111956 106108
rect 111956 106052 111960 106108
rect 111896 106048 111960 106052
rect 111976 106108 112040 106112
rect 111976 106052 111980 106108
rect 111980 106052 112036 106108
rect 112036 106052 112040 106108
rect 111976 106048 112040 106052
rect 142456 106108 142520 106112
rect 142456 106052 142460 106108
rect 142460 106052 142516 106108
rect 142516 106052 142520 106108
rect 142456 106048 142520 106052
rect 142536 106108 142600 106112
rect 142536 106052 142540 106108
rect 142540 106052 142596 106108
rect 142596 106052 142600 106108
rect 142536 106048 142600 106052
rect 142616 106108 142680 106112
rect 142616 106052 142620 106108
rect 142620 106052 142676 106108
rect 142676 106052 142680 106108
rect 142616 106048 142680 106052
rect 142696 106108 142760 106112
rect 142696 106052 142700 106108
rect 142700 106052 142756 106108
rect 142756 106052 142760 106108
rect 142696 106048 142760 106052
rect 173176 106108 173240 106112
rect 173176 106052 173180 106108
rect 173180 106052 173236 106108
rect 173236 106052 173240 106108
rect 173176 106048 173240 106052
rect 173256 106108 173320 106112
rect 173256 106052 173260 106108
rect 173260 106052 173316 106108
rect 173316 106052 173320 106108
rect 173256 106048 173320 106052
rect 173336 106108 173400 106112
rect 173336 106052 173340 106108
rect 173340 106052 173396 106108
rect 173396 106052 173400 106108
rect 173336 106048 173400 106052
rect 173416 106108 173480 106112
rect 173416 106052 173420 106108
rect 173420 106052 173476 106108
rect 173476 106052 173480 106108
rect 173416 106048 173480 106052
rect 4216 105564 4280 105568
rect 4216 105508 4220 105564
rect 4220 105508 4276 105564
rect 4276 105508 4280 105564
rect 4216 105504 4280 105508
rect 4296 105564 4360 105568
rect 4296 105508 4300 105564
rect 4300 105508 4356 105564
rect 4356 105508 4360 105564
rect 4296 105504 4360 105508
rect 4376 105564 4440 105568
rect 4376 105508 4380 105564
rect 4380 105508 4436 105564
rect 4436 105508 4440 105564
rect 4376 105504 4440 105508
rect 4456 105564 4520 105568
rect 4456 105508 4460 105564
rect 4460 105508 4516 105564
rect 4516 105508 4520 105564
rect 4456 105504 4520 105508
rect 34936 105564 35000 105568
rect 34936 105508 34940 105564
rect 34940 105508 34996 105564
rect 34996 105508 35000 105564
rect 34936 105504 35000 105508
rect 35016 105564 35080 105568
rect 35016 105508 35020 105564
rect 35020 105508 35076 105564
rect 35076 105508 35080 105564
rect 35016 105504 35080 105508
rect 35096 105564 35160 105568
rect 35096 105508 35100 105564
rect 35100 105508 35156 105564
rect 35156 105508 35160 105564
rect 35096 105504 35160 105508
rect 35176 105564 35240 105568
rect 35176 105508 35180 105564
rect 35180 105508 35236 105564
rect 35236 105508 35240 105564
rect 35176 105504 35240 105508
rect 65656 105564 65720 105568
rect 65656 105508 65660 105564
rect 65660 105508 65716 105564
rect 65716 105508 65720 105564
rect 65656 105504 65720 105508
rect 65736 105564 65800 105568
rect 65736 105508 65740 105564
rect 65740 105508 65796 105564
rect 65796 105508 65800 105564
rect 65736 105504 65800 105508
rect 65816 105564 65880 105568
rect 65816 105508 65820 105564
rect 65820 105508 65876 105564
rect 65876 105508 65880 105564
rect 65816 105504 65880 105508
rect 65896 105564 65960 105568
rect 65896 105508 65900 105564
rect 65900 105508 65956 105564
rect 65956 105508 65960 105564
rect 65896 105504 65960 105508
rect 96376 105564 96440 105568
rect 96376 105508 96380 105564
rect 96380 105508 96436 105564
rect 96436 105508 96440 105564
rect 96376 105504 96440 105508
rect 96456 105564 96520 105568
rect 96456 105508 96460 105564
rect 96460 105508 96516 105564
rect 96516 105508 96520 105564
rect 96456 105504 96520 105508
rect 96536 105564 96600 105568
rect 96536 105508 96540 105564
rect 96540 105508 96596 105564
rect 96596 105508 96600 105564
rect 96536 105504 96600 105508
rect 96616 105564 96680 105568
rect 96616 105508 96620 105564
rect 96620 105508 96676 105564
rect 96676 105508 96680 105564
rect 96616 105504 96680 105508
rect 127096 105564 127160 105568
rect 127096 105508 127100 105564
rect 127100 105508 127156 105564
rect 127156 105508 127160 105564
rect 127096 105504 127160 105508
rect 127176 105564 127240 105568
rect 127176 105508 127180 105564
rect 127180 105508 127236 105564
rect 127236 105508 127240 105564
rect 127176 105504 127240 105508
rect 127256 105564 127320 105568
rect 127256 105508 127260 105564
rect 127260 105508 127316 105564
rect 127316 105508 127320 105564
rect 127256 105504 127320 105508
rect 127336 105564 127400 105568
rect 127336 105508 127340 105564
rect 127340 105508 127396 105564
rect 127396 105508 127400 105564
rect 127336 105504 127400 105508
rect 157816 105564 157880 105568
rect 157816 105508 157820 105564
rect 157820 105508 157876 105564
rect 157876 105508 157880 105564
rect 157816 105504 157880 105508
rect 157896 105564 157960 105568
rect 157896 105508 157900 105564
rect 157900 105508 157956 105564
rect 157956 105508 157960 105564
rect 157896 105504 157960 105508
rect 157976 105564 158040 105568
rect 157976 105508 157980 105564
rect 157980 105508 158036 105564
rect 158036 105508 158040 105564
rect 157976 105504 158040 105508
rect 158056 105564 158120 105568
rect 158056 105508 158060 105564
rect 158060 105508 158116 105564
rect 158116 105508 158120 105564
rect 158056 105504 158120 105508
rect 19576 105020 19640 105024
rect 19576 104964 19580 105020
rect 19580 104964 19636 105020
rect 19636 104964 19640 105020
rect 19576 104960 19640 104964
rect 19656 105020 19720 105024
rect 19656 104964 19660 105020
rect 19660 104964 19716 105020
rect 19716 104964 19720 105020
rect 19656 104960 19720 104964
rect 19736 105020 19800 105024
rect 19736 104964 19740 105020
rect 19740 104964 19796 105020
rect 19796 104964 19800 105020
rect 19736 104960 19800 104964
rect 19816 105020 19880 105024
rect 19816 104964 19820 105020
rect 19820 104964 19876 105020
rect 19876 104964 19880 105020
rect 19816 104960 19880 104964
rect 50296 105020 50360 105024
rect 50296 104964 50300 105020
rect 50300 104964 50356 105020
rect 50356 104964 50360 105020
rect 50296 104960 50360 104964
rect 50376 105020 50440 105024
rect 50376 104964 50380 105020
rect 50380 104964 50436 105020
rect 50436 104964 50440 105020
rect 50376 104960 50440 104964
rect 50456 105020 50520 105024
rect 50456 104964 50460 105020
rect 50460 104964 50516 105020
rect 50516 104964 50520 105020
rect 50456 104960 50520 104964
rect 50536 105020 50600 105024
rect 50536 104964 50540 105020
rect 50540 104964 50596 105020
rect 50596 104964 50600 105020
rect 50536 104960 50600 104964
rect 81016 105020 81080 105024
rect 81016 104964 81020 105020
rect 81020 104964 81076 105020
rect 81076 104964 81080 105020
rect 81016 104960 81080 104964
rect 81096 105020 81160 105024
rect 81096 104964 81100 105020
rect 81100 104964 81156 105020
rect 81156 104964 81160 105020
rect 81096 104960 81160 104964
rect 81176 105020 81240 105024
rect 81176 104964 81180 105020
rect 81180 104964 81236 105020
rect 81236 104964 81240 105020
rect 81176 104960 81240 104964
rect 81256 105020 81320 105024
rect 81256 104964 81260 105020
rect 81260 104964 81316 105020
rect 81316 104964 81320 105020
rect 81256 104960 81320 104964
rect 111736 105020 111800 105024
rect 111736 104964 111740 105020
rect 111740 104964 111796 105020
rect 111796 104964 111800 105020
rect 111736 104960 111800 104964
rect 111816 105020 111880 105024
rect 111816 104964 111820 105020
rect 111820 104964 111876 105020
rect 111876 104964 111880 105020
rect 111816 104960 111880 104964
rect 111896 105020 111960 105024
rect 111896 104964 111900 105020
rect 111900 104964 111956 105020
rect 111956 104964 111960 105020
rect 111896 104960 111960 104964
rect 111976 105020 112040 105024
rect 111976 104964 111980 105020
rect 111980 104964 112036 105020
rect 112036 104964 112040 105020
rect 111976 104960 112040 104964
rect 142456 105020 142520 105024
rect 142456 104964 142460 105020
rect 142460 104964 142516 105020
rect 142516 104964 142520 105020
rect 142456 104960 142520 104964
rect 142536 105020 142600 105024
rect 142536 104964 142540 105020
rect 142540 104964 142596 105020
rect 142596 104964 142600 105020
rect 142536 104960 142600 104964
rect 142616 105020 142680 105024
rect 142616 104964 142620 105020
rect 142620 104964 142676 105020
rect 142676 104964 142680 105020
rect 142616 104960 142680 104964
rect 142696 105020 142760 105024
rect 142696 104964 142700 105020
rect 142700 104964 142756 105020
rect 142756 104964 142760 105020
rect 142696 104960 142760 104964
rect 173176 105020 173240 105024
rect 173176 104964 173180 105020
rect 173180 104964 173236 105020
rect 173236 104964 173240 105020
rect 173176 104960 173240 104964
rect 173256 105020 173320 105024
rect 173256 104964 173260 105020
rect 173260 104964 173316 105020
rect 173316 104964 173320 105020
rect 173256 104960 173320 104964
rect 173336 105020 173400 105024
rect 173336 104964 173340 105020
rect 173340 104964 173396 105020
rect 173396 104964 173400 105020
rect 173336 104960 173400 104964
rect 173416 105020 173480 105024
rect 173416 104964 173420 105020
rect 173420 104964 173476 105020
rect 173476 104964 173480 105020
rect 173416 104960 173480 104964
rect 4216 104476 4280 104480
rect 4216 104420 4220 104476
rect 4220 104420 4276 104476
rect 4276 104420 4280 104476
rect 4216 104416 4280 104420
rect 4296 104476 4360 104480
rect 4296 104420 4300 104476
rect 4300 104420 4356 104476
rect 4356 104420 4360 104476
rect 4296 104416 4360 104420
rect 4376 104476 4440 104480
rect 4376 104420 4380 104476
rect 4380 104420 4436 104476
rect 4436 104420 4440 104476
rect 4376 104416 4440 104420
rect 4456 104476 4520 104480
rect 4456 104420 4460 104476
rect 4460 104420 4516 104476
rect 4516 104420 4520 104476
rect 4456 104416 4520 104420
rect 34936 104476 35000 104480
rect 34936 104420 34940 104476
rect 34940 104420 34996 104476
rect 34996 104420 35000 104476
rect 34936 104416 35000 104420
rect 35016 104476 35080 104480
rect 35016 104420 35020 104476
rect 35020 104420 35076 104476
rect 35076 104420 35080 104476
rect 35016 104416 35080 104420
rect 35096 104476 35160 104480
rect 35096 104420 35100 104476
rect 35100 104420 35156 104476
rect 35156 104420 35160 104476
rect 35096 104416 35160 104420
rect 35176 104476 35240 104480
rect 35176 104420 35180 104476
rect 35180 104420 35236 104476
rect 35236 104420 35240 104476
rect 35176 104416 35240 104420
rect 65656 104476 65720 104480
rect 65656 104420 65660 104476
rect 65660 104420 65716 104476
rect 65716 104420 65720 104476
rect 65656 104416 65720 104420
rect 65736 104476 65800 104480
rect 65736 104420 65740 104476
rect 65740 104420 65796 104476
rect 65796 104420 65800 104476
rect 65736 104416 65800 104420
rect 65816 104476 65880 104480
rect 65816 104420 65820 104476
rect 65820 104420 65876 104476
rect 65876 104420 65880 104476
rect 65816 104416 65880 104420
rect 65896 104476 65960 104480
rect 65896 104420 65900 104476
rect 65900 104420 65956 104476
rect 65956 104420 65960 104476
rect 65896 104416 65960 104420
rect 96376 104476 96440 104480
rect 96376 104420 96380 104476
rect 96380 104420 96436 104476
rect 96436 104420 96440 104476
rect 96376 104416 96440 104420
rect 96456 104476 96520 104480
rect 96456 104420 96460 104476
rect 96460 104420 96516 104476
rect 96516 104420 96520 104476
rect 96456 104416 96520 104420
rect 96536 104476 96600 104480
rect 96536 104420 96540 104476
rect 96540 104420 96596 104476
rect 96596 104420 96600 104476
rect 96536 104416 96600 104420
rect 96616 104476 96680 104480
rect 96616 104420 96620 104476
rect 96620 104420 96676 104476
rect 96676 104420 96680 104476
rect 96616 104416 96680 104420
rect 127096 104476 127160 104480
rect 127096 104420 127100 104476
rect 127100 104420 127156 104476
rect 127156 104420 127160 104476
rect 127096 104416 127160 104420
rect 127176 104476 127240 104480
rect 127176 104420 127180 104476
rect 127180 104420 127236 104476
rect 127236 104420 127240 104476
rect 127176 104416 127240 104420
rect 127256 104476 127320 104480
rect 127256 104420 127260 104476
rect 127260 104420 127316 104476
rect 127316 104420 127320 104476
rect 127256 104416 127320 104420
rect 127336 104476 127400 104480
rect 127336 104420 127340 104476
rect 127340 104420 127396 104476
rect 127396 104420 127400 104476
rect 127336 104416 127400 104420
rect 157816 104476 157880 104480
rect 157816 104420 157820 104476
rect 157820 104420 157876 104476
rect 157876 104420 157880 104476
rect 157816 104416 157880 104420
rect 157896 104476 157960 104480
rect 157896 104420 157900 104476
rect 157900 104420 157956 104476
rect 157956 104420 157960 104476
rect 157896 104416 157960 104420
rect 157976 104476 158040 104480
rect 157976 104420 157980 104476
rect 157980 104420 158036 104476
rect 158036 104420 158040 104476
rect 157976 104416 158040 104420
rect 158056 104476 158120 104480
rect 158056 104420 158060 104476
rect 158060 104420 158116 104476
rect 158116 104420 158120 104476
rect 158056 104416 158120 104420
rect 19576 103932 19640 103936
rect 19576 103876 19580 103932
rect 19580 103876 19636 103932
rect 19636 103876 19640 103932
rect 19576 103872 19640 103876
rect 19656 103932 19720 103936
rect 19656 103876 19660 103932
rect 19660 103876 19716 103932
rect 19716 103876 19720 103932
rect 19656 103872 19720 103876
rect 19736 103932 19800 103936
rect 19736 103876 19740 103932
rect 19740 103876 19796 103932
rect 19796 103876 19800 103932
rect 19736 103872 19800 103876
rect 19816 103932 19880 103936
rect 19816 103876 19820 103932
rect 19820 103876 19876 103932
rect 19876 103876 19880 103932
rect 19816 103872 19880 103876
rect 50296 103932 50360 103936
rect 50296 103876 50300 103932
rect 50300 103876 50356 103932
rect 50356 103876 50360 103932
rect 50296 103872 50360 103876
rect 50376 103932 50440 103936
rect 50376 103876 50380 103932
rect 50380 103876 50436 103932
rect 50436 103876 50440 103932
rect 50376 103872 50440 103876
rect 50456 103932 50520 103936
rect 50456 103876 50460 103932
rect 50460 103876 50516 103932
rect 50516 103876 50520 103932
rect 50456 103872 50520 103876
rect 50536 103932 50600 103936
rect 50536 103876 50540 103932
rect 50540 103876 50596 103932
rect 50596 103876 50600 103932
rect 50536 103872 50600 103876
rect 81016 103932 81080 103936
rect 81016 103876 81020 103932
rect 81020 103876 81076 103932
rect 81076 103876 81080 103932
rect 81016 103872 81080 103876
rect 81096 103932 81160 103936
rect 81096 103876 81100 103932
rect 81100 103876 81156 103932
rect 81156 103876 81160 103932
rect 81096 103872 81160 103876
rect 81176 103932 81240 103936
rect 81176 103876 81180 103932
rect 81180 103876 81236 103932
rect 81236 103876 81240 103932
rect 81176 103872 81240 103876
rect 81256 103932 81320 103936
rect 81256 103876 81260 103932
rect 81260 103876 81316 103932
rect 81316 103876 81320 103932
rect 81256 103872 81320 103876
rect 111736 103932 111800 103936
rect 111736 103876 111740 103932
rect 111740 103876 111796 103932
rect 111796 103876 111800 103932
rect 111736 103872 111800 103876
rect 111816 103932 111880 103936
rect 111816 103876 111820 103932
rect 111820 103876 111876 103932
rect 111876 103876 111880 103932
rect 111816 103872 111880 103876
rect 111896 103932 111960 103936
rect 111896 103876 111900 103932
rect 111900 103876 111956 103932
rect 111956 103876 111960 103932
rect 111896 103872 111960 103876
rect 111976 103932 112040 103936
rect 111976 103876 111980 103932
rect 111980 103876 112036 103932
rect 112036 103876 112040 103932
rect 111976 103872 112040 103876
rect 142456 103932 142520 103936
rect 142456 103876 142460 103932
rect 142460 103876 142516 103932
rect 142516 103876 142520 103932
rect 142456 103872 142520 103876
rect 142536 103932 142600 103936
rect 142536 103876 142540 103932
rect 142540 103876 142596 103932
rect 142596 103876 142600 103932
rect 142536 103872 142600 103876
rect 142616 103932 142680 103936
rect 142616 103876 142620 103932
rect 142620 103876 142676 103932
rect 142676 103876 142680 103932
rect 142616 103872 142680 103876
rect 142696 103932 142760 103936
rect 142696 103876 142700 103932
rect 142700 103876 142756 103932
rect 142756 103876 142760 103932
rect 142696 103872 142760 103876
rect 173176 103932 173240 103936
rect 173176 103876 173180 103932
rect 173180 103876 173236 103932
rect 173236 103876 173240 103932
rect 173176 103872 173240 103876
rect 173256 103932 173320 103936
rect 173256 103876 173260 103932
rect 173260 103876 173316 103932
rect 173316 103876 173320 103932
rect 173256 103872 173320 103876
rect 173336 103932 173400 103936
rect 173336 103876 173340 103932
rect 173340 103876 173396 103932
rect 173396 103876 173400 103932
rect 173336 103872 173400 103876
rect 173416 103932 173480 103936
rect 173416 103876 173420 103932
rect 173420 103876 173476 103932
rect 173476 103876 173480 103932
rect 173416 103872 173480 103876
rect 4216 103388 4280 103392
rect 4216 103332 4220 103388
rect 4220 103332 4276 103388
rect 4276 103332 4280 103388
rect 4216 103328 4280 103332
rect 4296 103388 4360 103392
rect 4296 103332 4300 103388
rect 4300 103332 4356 103388
rect 4356 103332 4360 103388
rect 4296 103328 4360 103332
rect 4376 103388 4440 103392
rect 4376 103332 4380 103388
rect 4380 103332 4436 103388
rect 4436 103332 4440 103388
rect 4376 103328 4440 103332
rect 4456 103388 4520 103392
rect 4456 103332 4460 103388
rect 4460 103332 4516 103388
rect 4516 103332 4520 103388
rect 4456 103328 4520 103332
rect 34936 103388 35000 103392
rect 34936 103332 34940 103388
rect 34940 103332 34996 103388
rect 34996 103332 35000 103388
rect 34936 103328 35000 103332
rect 35016 103388 35080 103392
rect 35016 103332 35020 103388
rect 35020 103332 35076 103388
rect 35076 103332 35080 103388
rect 35016 103328 35080 103332
rect 35096 103388 35160 103392
rect 35096 103332 35100 103388
rect 35100 103332 35156 103388
rect 35156 103332 35160 103388
rect 35096 103328 35160 103332
rect 35176 103388 35240 103392
rect 35176 103332 35180 103388
rect 35180 103332 35236 103388
rect 35236 103332 35240 103388
rect 35176 103328 35240 103332
rect 65656 103388 65720 103392
rect 65656 103332 65660 103388
rect 65660 103332 65716 103388
rect 65716 103332 65720 103388
rect 65656 103328 65720 103332
rect 65736 103388 65800 103392
rect 65736 103332 65740 103388
rect 65740 103332 65796 103388
rect 65796 103332 65800 103388
rect 65736 103328 65800 103332
rect 65816 103388 65880 103392
rect 65816 103332 65820 103388
rect 65820 103332 65876 103388
rect 65876 103332 65880 103388
rect 65816 103328 65880 103332
rect 65896 103388 65960 103392
rect 65896 103332 65900 103388
rect 65900 103332 65956 103388
rect 65956 103332 65960 103388
rect 65896 103328 65960 103332
rect 96376 103388 96440 103392
rect 96376 103332 96380 103388
rect 96380 103332 96436 103388
rect 96436 103332 96440 103388
rect 96376 103328 96440 103332
rect 96456 103388 96520 103392
rect 96456 103332 96460 103388
rect 96460 103332 96516 103388
rect 96516 103332 96520 103388
rect 96456 103328 96520 103332
rect 96536 103388 96600 103392
rect 96536 103332 96540 103388
rect 96540 103332 96596 103388
rect 96596 103332 96600 103388
rect 96536 103328 96600 103332
rect 96616 103388 96680 103392
rect 96616 103332 96620 103388
rect 96620 103332 96676 103388
rect 96676 103332 96680 103388
rect 96616 103328 96680 103332
rect 127096 103388 127160 103392
rect 127096 103332 127100 103388
rect 127100 103332 127156 103388
rect 127156 103332 127160 103388
rect 127096 103328 127160 103332
rect 127176 103388 127240 103392
rect 127176 103332 127180 103388
rect 127180 103332 127236 103388
rect 127236 103332 127240 103388
rect 127176 103328 127240 103332
rect 127256 103388 127320 103392
rect 127256 103332 127260 103388
rect 127260 103332 127316 103388
rect 127316 103332 127320 103388
rect 127256 103328 127320 103332
rect 127336 103388 127400 103392
rect 127336 103332 127340 103388
rect 127340 103332 127396 103388
rect 127396 103332 127400 103388
rect 127336 103328 127400 103332
rect 157816 103388 157880 103392
rect 157816 103332 157820 103388
rect 157820 103332 157876 103388
rect 157876 103332 157880 103388
rect 157816 103328 157880 103332
rect 157896 103388 157960 103392
rect 157896 103332 157900 103388
rect 157900 103332 157956 103388
rect 157956 103332 157960 103388
rect 157896 103328 157960 103332
rect 157976 103388 158040 103392
rect 157976 103332 157980 103388
rect 157980 103332 158036 103388
rect 158036 103332 158040 103388
rect 157976 103328 158040 103332
rect 158056 103388 158120 103392
rect 158056 103332 158060 103388
rect 158060 103332 158116 103388
rect 158116 103332 158120 103388
rect 158056 103328 158120 103332
rect 19576 102844 19640 102848
rect 19576 102788 19580 102844
rect 19580 102788 19636 102844
rect 19636 102788 19640 102844
rect 19576 102784 19640 102788
rect 19656 102844 19720 102848
rect 19656 102788 19660 102844
rect 19660 102788 19716 102844
rect 19716 102788 19720 102844
rect 19656 102784 19720 102788
rect 19736 102844 19800 102848
rect 19736 102788 19740 102844
rect 19740 102788 19796 102844
rect 19796 102788 19800 102844
rect 19736 102784 19800 102788
rect 19816 102844 19880 102848
rect 19816 102788 19820 102844
rect 19820 102788 19876 102844
rect 19876 102788 19880 102844
rect 19816 102784 19880 102788
rect 50296 102844 50360 102848
rect 50296 102788 50300 102844
rect 50300 102788 50356 102844
rect 50356 102788 50360 102844
rect 50296 102784 50360 102788
rect 50376 102844 50440 102848
rect 50376 102788 50380 102844
rect 50380 102788 50436 102844
rect 50436 102788 50440 102844
rect 50376 102784 50440 102788
rect 50456 102844 50520 102848
rect 50456 102788 50460 102844
rect 50460 102788 50516 102844
rect 50516 102788 50520 102844
rect 50456 102784 50520 102788
rect 50536 102844 50600 102848
rect 50536 102788 50540 102844
rect 50540 102788 50596 102844
rect 50596 102788 50600 102844
rect 50536 102784 50600 102788
rect 81016 102844 81080 102848
rect 81016 102788 81020 102844
rect 81020 102788 81076 102844
rect 81076 102788 81080 102844
rect 81016 102784 81080 102788
rect 81096 102844 81160 102848
rect 81096 102788 81100 102844
rect 81100 102788 81156 102844
rect 81156 102788 81160 102844
rect 81096 102784 81160 102788
rect 81176 102844 81240 102848
rect 81176 102788 81180 102844
rect 81180 102788 81236 102844
rect 81236 102788 81240 102844
rect 81176 102784 81240 102788
rect 81256 102844 81320 102848
rect 81256 102788 81260 102844
rect 81260 102788 81316 102844
rect 81316 102788 81320 102844
rect 81256 102784 81320 102788
rect 111736 102844 111800 102848
rect 111736 102788 111740 102844
rect 111740 102788 111796 102844
rect 111796 102788 111800 102844
rect 111736 102784 111800 102788
rect 111816 102844 111880 102848
rect 111816 102788 111820 102844
rect 111820 102788 111876 102844
rect 111876 102788 111880 102844
rect 111816 102784 111880 102788
rect 111896 102844 111960 102848
rect 111896 102788 111900 102844
rect 111900 102788 111956 102844
rect 111956 102788 111960 102844
rect 111896 102784 111960 102788
rect 111976 102844 112040 102848
rect 111976 102788 111980 102844
rect 111980 102788 112036 102844
rect 112036 102788 112040 102844
rect 111976 102784 112040 102788
rect 142456 102844 142520 102848
rect 142456 102788 142460 102844
rect 142460 102788 142516 102844
rect 142516 102788 142520 102844
rect 142456 102784 142520 102788
rect 142536 102844 142600 102848
rect 142536 102788 142540 102844
rect 142540 102788 142596 102844
rect 142596 102788 142600 102844
rect 142536 102784 142600 102788
rect 142616 102844 142680 102848
rect 142616 102788 142620 102844
rect 142620 102788 142676 102844
rect 142676 102788 142680 102844
rect 142616 102784 142680 102788
rect 142696 102844 142760 102848
rect 142696 102788 142700 102844
rect 142700 102788 142756 102844
rect 142756 102788 142760 102844
rect 142696 102784 142760 102788
rect 173176 102844 173240 102848
rect 173176 102788 173180 102844
rect 173180 102788 173236 102844
rect 173236 102788 173240 102844
rect 173176 102784 173240 102788
rect 173256 102844 173320 102848
rect 173256 102788 173260 102844
rect 173260 102788 173316 102844
rect 173316 102788 173320 102844
rect 173256 102784 173320 102788
rect 173336 102844 173400 102848
rect 173336 102788 173340 102844
rect 173340 102788 173396 102844
rect 173396 102788 173400 102844
rect 173336 102784 173400 102788
rect 173416 102844 173480 102848
rect 173416 102788 173420 102844
rect 173420 102788 173476 102844
rect 173476 102788 173480 102844
rect 173416 102784 173480 102788
rect 4216 102300 4280 102304
rect 4216 102244 4220 102300
rect 4220 102244 4276 102300
rect 4276 102244 4280 102300
rect 4216 102240 4280 102244
rect 4296 102300 4360 102304
rect 4296 102244 4300 102300
rect 4300 102244 4356 102300
rect 4356 102244 4360 102300
rect 4296 102240 4360 102244
rect 4376 102300 4440 102304
rect 4376 102244 4380 102300
rect 4380 102244 4436 102300
rect 4436 102244 4440 102300
rect 4376 102240 4440 102244
rect 4456 102300 4520 102304
rect 4456 102244 4460 102300
rect 4460 102244 4516 102300
rect 4516 102244 4520 102300
rect 4456 102240 4520 102244
rect 34936 102300 35000 102304
rect 34936 102244 34940 102300
rect 34940 102244 34996 102300
rect 34996 102244 35000 102300
rect 34936 102240 35000 102244
rect 35016 102300 35080 102304
rect 35016 102244 35020 102300
rect 35020 102244 35076 102300
rect 35076 102244 35080 102300
rect 35016 102240 35080 102244
rect 35096 102300 35160 102304
rect 35096 102244 35100 102300
rect 35100 102244 35156 102300
rect 35156 102244 35160 102300
rect 35096 102240 35160 102244
rect 35176 102300 35240 102304
rect 35176 102244 35180 102300
rect 35180 102244 35236 102300
rect 35236 102244 35240 102300
rect 35176 102240 35240 102244
rect 65656 102300 65720 102304
rect 65656 102244 65660 102300
rect 65660 102244 65716 102300
rect 65716 102244 65720 102300
rect 65656 102240 65720 102244
rect 65736 102300 65800 102304
rect 65736 102244 65740 102300
rect 65740 102244 65796 102300
rect 65796 102244 65800 102300
rect 65736 102240 65800 102244
rect 65816 102300 65880 102304
rect 65816 102244 65820 102300
rect 65820 102244 65876 102300
rect 65876 102244 65880 102300
rect 65816 102240 65880 102244
rect 65896 102300 65960 102304
rect 65896 102244 65900 102300
rect 65900 102244 65956 102300
rect 65956 102244 65960 102300
rect 65896 102240 65960 102244
rect 96376 102300 96440 102304
rect 96376 102244 96380 102300
rect 96380 102244 96436 102300
rect 96436 102244 96440 102300
rect 96376 102240 96440 102244
rect 96456 102300 96520 102304
rect 96456 102244 96460 102300
rect 96460 102244 96516 102300
rect 96516 102244 96520 102300
rect 96456 102240 96520 102244
rect 96536 102300 96600 102304
rect 96536 102244 96540 102300
rect 96540 102244 96596 102300
rect 96596 102244 96600 102300
rect 96536 102240 96600 102244
rect 96616 102300 96680 102304
rect 96616 102244 96620 102300
rect 96620 102244 96676 102300
rect 96676 102244 96680 102300
rect 96616 102240 96680 102244
rect 127096 102300 127160 102304
rect 127096 102244 127100 102300
rect 127100 102244 127156 102300
rect 127156 102244 127160 102300
rect 127096 102240 127160 102244
rect 127176 102300 127240 102304
rect 127176 102244 127180 102300
rect 127180 102244 127236 102300
rect 127236 102244 127240 102300
rect 127176 102240 127240 102244
rect 127256 102300 127320 102304
rect 127256 102244 127260 102300
rect 127260 102244 127316 102300
rect 127316 102244 127320 102300
rect 127256 102240 127320 102244
rect 127336 102300 127400 102304
rect 127336 102244 127340 102300
rect 127340 102244 127396 102300
rect 127396 102244 127400 102300
rect 127336 102240 127400 102244
rect 157816 102300 157880 102304
rect 157816 102244 157820 102300
rect 157820 102244 157876 102300
rect 157876 102244 157880 102300
rect 157816 102240 157880 102244
rect 157896 102300 157960 102304
rect 157896 102244 157900 102300
rect 157900 102244 157956 102300
rect 157956 102244 157960 102300
rect 157896 102240 157960 102244
rect 157976 102300 158040 102304
rect 157976 102244 157980 102300
rect 157980 102244 158036 102300
rect 158036 102244 158040 102300
rect 157976 102240 158040 102244
rect 158056 102300 158120 102304
rect 158056 102244 158060 102300
rect 158060 102244 158116 102300
rect 158116 102244 158120 102300
rect 158056 102240 158120 102244
rect 19576 101756 19640 101760
rect 19576 101700 19580 101756
rect 19580 101700 19636 101756
rect 19636 101700 19640 101756
rect 19576 101696 19640 101700
rect 19656 101756 19720 101760
rect 19656 101700 19660 101756
rect 19660 101700 19716 101756
rect 19716 101700 19720 101756
rect 19656 101696 19720 101700
rect 19736 101756 19800 101760
rect 19736 101700 19740 101756
rect 19740 101700 19796 101756
rect 19796 101700 19800 101756
rect 19736 101696 19800 101700
rect 19816 101756 19880 101760
rect 19816 101700 19820 101756
rect 19820 101700 19876 101756
rect 19876 101700 19880 101756
rect 19816 101696 19880 101700
rect 50296 101756 50360 101760
rect 50296 101700 50300 101756
rect 50300 101700 50356 101756
rect 50356 101700 50360 101756
rect 50296 101696 50360 101700
rect 50376 101756 50440 101760
rect 50376 101700 50380 101756
rect 50380 101700 50436 101756
rect 50436 101700 50440 101756
rect 50376 101696 50440 101700
rect 50456 101756 50520 101760
rect 50456 101700 50460 101756
rect 50460 101700 50516 101756
rect 50516 101700 50520 101756
rect 50456 101696 50520 101700
rect 50536 101756 50600 101760
rect 50536 101700 50540 101756
rect 50540 101700 50596 101756
rect 50596 101700 50600 101756
rect 50536 101696 50600 101700
rect 81016 101756 81080 101760
rect 81016 101700 81020 101756
rect 81020 101700 81076 101756
rect 81076 101700 81080 101756
rect 81016 101696 81080 101700
rect 81096 101756 81160 101760
rect 81096 101700 81100 101756
rect 81100 101700 81156 101756
rect 81156 101700 81160 101756
rect 81096 101696 81160 101700
rect 81176 101756 81240 101760
rect 81176 101700 81180 101756
rect 81180 101700 81236 101756
rect 81236 101700 81240 101756
rect 81176 101696 81240 101700
rect 81256 101756 81320 101760
rect 81256 101700 81260 101756
rect 81260 101700 81316 101756
rect 81316 101700 81320 101756
rect 81256 101696 81320 101700
rect 111736 101756 111800 101760
rect 111736 101700 111740 101756
rect 111740 101700 111796 101756
rect 111796 101700 111800 101756
rect 111736 101696 111800 101700
rect 111816 101756 111880 101760
rect 111816 101700 111820 101756
rect 111820 101700 111876 101756
rect 111876 101700 111880 101756
rect 111816 101696 111880 101700
rect 111896 101756 111960 101760
rect 111896 101700 111900 101756
rect 111900 101700 111956 101756
rect 111956 101700 111960 101756
rect 111896 101696 111960 101700
rect 111976 101756 112040 101760
rect 111976 101700 111980 101756
rect 111980 101700 112036 101756
rect 112036 101700 112040 101756
rect 111976 101696 112040 101700
rect 142456 101756 142520 101760
rect 142456 101700 142460 101756
rect 142460 101700 142516 101756
rect 142516 101700 142520 101756
rect 142456 101696 142520 101700
rect 142536 101756 142600 101760
rect 142536 101700 142540 101756
rect 142540 101700 142596 101756
rect 142596 101700 142600 101756
rect 142536 101696 142600 101700
rect 142616 101756 142680 101760
rect 142616 101700 142620 101756
rect 142620 101700 142676 101756
rect 142676 101700 142680 101756
rect 142616 101696 142680 101700
rect 142696 101756 142760 101760
rect 142696 101700 142700 101756
rect 142700 101700 142756 101756
rect 142756 101700 142760 101756
rect 142696 101696 142760 101700
rect 173176 101756 173240 101760
rect 173176 101700 173180 101756
rect 173180 101700 173236 101756
rect 173236 101700 173240 101756
rect 173176 101696 173240 101700
rect 173256 101756 173320 101760
rect 173256 101700 173260 101756
rect 173260 101700 173316 101756
rect 173316 101700 173320 101756
rect 173256 101696 173320 101700
rect 173336 101756 173400 101760
rect 173336 101700 173340 101756
rect 173340 101700 173396 101756
rect 173396 101700 173400 101756
rect 173336 101696 173400 101700
rect 173416 101756 173480 101760
rect 173416 101700 173420 101756
rect 173420 101700 173476 101756
rect 173476 101700 173480 101756
rect 173416 101696 173480 101700
rect 4216 101212 4280 101216
rect 4216 101156 4220 101212
rect 4220 101156 4276 101212
rect 4276 101156 4280 101212
rect 4216 101152 4280 101156
rect 4296 101212 4360 101216
rect 4296 101156 4300 101212
rect 4300 101156 4356 101212
rect 4356 101156 4360 101212
rect 4296 101152 4360 101156
rect 4376 101212 4440 101216
rect 4376 101156 4380 101212
rect 4380 101156 4436 101212
rect 4436 101156 4440 101212
rect 4376 101152 4440 101156
rect 4456 101212 4520 101216
rect 4456 101156 4460 101212
rect 4460 101156 4516 101212
rect 4516 101156 4520 101212
rect 4456 101152 4520 101156
rect 34936 101212 35000 101216
rect 34936 101156 34940 101212
rect 34940 101156 34996 101212
rect 34996 101156 35000 101212
rect 34936 101152 35000 101156
rect 35016 101212 35080 101216
rect 35016 101156 35020 101212
rect 35020 101156 35076 101212
rect 35076 101156 35080 101212
rect 35016 101152 35080 101156
rect 35096 101212 35160 101216
rect 35096 101156 35100 101212
rect 35100 101156 35156 101212
rect 35156 101156 35160 101212
rect 35096 101152 35160 101156
rect 35176 101212 35240 101216
rect 35176 101156 35180 101212
rect 35180 101156 35236 101212
rect 35236 101156 35240 101212
rect 35176 101152 35240 101156
rect 65656 101212 65720 101216
rect 65656 101156 65660 101212
rect 65660 101156 65716 101212
rect 65716 101156 65720 101212
rect 65656 101152 65720 101156
rect 65736 101212 65800 101216
rect 65736 101156 65740 101212
rect 65740 101156 65796 101212
rect 65796 101156 65800 101212
rect 65736 101152 65800 101156
rect 65816 101212 65880 101216
rect 65816 101156 65820 101212
rect 65820 101156 65876 101212
rect 65876 101156 65880 101212
rect 65816 101152 65880 101156
rect 65896 101212 65960 101216
rect 65896 101156 65900 101212
rect 65900 101156 65956 101212
rect 65956 101156 65960 101212
rect 65896 101152 65960 101156
rect 96376 101212 96440 101216
rect 96376 101156 96380 101212
rect 96380 101156 96436 101212
rect 96436 101156 96440 101212
rect 96376 101152 96440 101156
rect 96456 101212 96520 101216
rect 96456 101156 96460 101212
rect 96460 101156 96516 101212
rect 96516 101156 96520 101212
rect 96456 101152 96520 101156
rect 96536 101212 96600 101216
rect 96536 101156 96540 101212
rect 96540 101156 96596 101212
rect 96596 101156 96600 101212
rect 96536 101152 96600 101156
rect 96616 101212 96680 101216
rect 96616 101156 96620 101212
rect 96620 101156 96676 101212
rect 96676 101156 96680 101212
rect 96616 101152 96680 101156
rect 127096 101212 127160 101216
rect 127096 101156 127100 101212
rect 127100 101156 127156 101212
rect 127156 101156 127160 101212
rect 127096 101152 127160 101156
rect 127176 101212 127240 101216
rect 127176 101156 127180 101212
rect 127180 101156 127236 101212
rect 127236 101156 127240 101212
rect 127176 101152 127240 101156
rect 127256 101212 127320 101216
rect 127256 101156 127260 101212
rect 127260 101156 127316 101212
rect 127316 101156 127320 101212
rect 127256 101152 127320 101156
rect 127336 101212 127400 101216
rect 127336 101156 127340 101212
rect 127340 101156 127396 101212
rect 127396 101156 127400 101212
rect 127336 101152 127400 101156
rect 157816 101212 157880 101216
rect 157816 101156 157820 101212
rect 157820 101156 157876 101212
rect 157876 101156 157880 101212
rect 157816 101152 157880 101156
rect 157896 101212 157960 101216
rect 157896 101156 157900 101212
rect 157900 101156 157956 101212
rect 157956 101156 157960 101212
rect 157896 101152 157960 101156
rect 157976 101212 158040 101216
rect 157976 101156 157980 101212
rect 157980 101156 158036 101212
rect 158036 101156 158040 101212
rect 157976 101152 158040 101156
rect 158056 101212 158120 101216
rect 158056 101156 158060 101212
rect 158060 101156 158116 101212
rect 158116 101156 158120 101212
rect 158056 101152 158120 101156
rect 19576 100668 19640 100672
rect 19576 100612 19580 100668
rect 19580 100612 19636 100668
rect 19636 100612 19640 100668
rect 19576 100608 19640 100612
rect 19656 100668 19720 100672
rect 19656 100612 19660 100668
rect 19660 100612 19716 100668
rect 19716 100612 19720 100668
rect 19656 100608 19720 100612
rect 19736 100668 19800 100672
rect 19736 100612 19740 100668
rect 19740 100612 19796 100668
rect 19796 100612 19800 100668
rect 19736 100608 19800 100612
rect 19816 100668 19880 100672
rect 19816 100612 19820 100668
rect 19820 100612 19876 100668
rect 19876 100612 19880 100668
rect 19816 100608 19880 100612
rect 50296 100668 50360 100672
rect 50296 100612 50300 100668
rect 50300 100612 50356 100668
rect 50356 100612 50360 100668
rect 50296 100608 50360 100612
rect 50376 100668 50440 100672
rect 50376 100612 50380 100668
rect 50380 100612 50436 100668
rect 50436 100612 50440 100668
rect 50376 100608 50440 100612
rect 50456 100668 50520 100672
rect 50456 100612 50460 100668
rect 50460 100612 50516 100668
rect 50516 100612 50520 100668
rect 50456 100608 50520 100612
rect 50536 100668 50600 100672
rect 50536 100612 50540 100668
rect 50540 100612 50596 100668
rect 50596 100612 50600 100668
rect 50536 100608 50600 100612
rect 81016 100668 81080 100672
rect 81016 100612 81020 100668
rect 81020 100612 81076 100668
rect 81076 100612 81080 100668
rect 81016 100608 81080 100612
rect 81096 100668 81160 100672
rect 81096 100612 81100 100668
rect 81100 100612 81156 100668
rect 81156 100612 81160 100668
rect 81096 100608 81160 100612
rect 81176 100668 81240 100672
rect 81176 100612 81180 100668
rect 81180 100612 81236 100668
rect 81236 100612 81240 100668
rect 81176 100608 81240 100612
rect 81256 100668 81320 100672
rect 81256 100612 81260 100668
rect 81260 100612 81316 100668
rect 81316 100612 81320 100668
rect 81256 100608 81320 100612
rect 111736 100668 111800 100672
rect 111736 100612 111740 100668
rect 111740 100612 111796 100668
rect 111796 100612 111800 100668
rect 111736 100608 111800 100612
rect 111816 100668 111880 100672
rect 111816 100612 111820 100668
rect 111820 100612 111876 100668
rect 111876 100612 111880 100668
rect 111816 100608 111880 100612
rect 111896 100668 111960 100672
rect 111896 100612 111900 100668
rect 111900 100612 111956 100668
rect 111956 100612 111960 100668
rect 111896 100608 111960 100612
rect 111976 100668 112040 100672
rect 111976 100612 111980 100668
rect 111980 100612 112036 100668
rect 112036 100612 112040 100668
rect 111976 100608 112040 100612
rect 142456 100668 142520 100672
rect 142456 100612 142460 100668
rect 142460 100612 142516 100668
rect 142516 100612 142520 100668
rect 142456 100608 142520 100612
rect 142536 100668 142600 100672
rect 142536 100612 142540 100668
rect 142540 100612 142596 100668
rect 142596 100612 142600 100668
rect 142536 100608 142600 100612
rect 142616 100668 142680 100672
rect 142616 100612 142620 100668
rect 142620 100612 142676 100668
rect 142676 100612 142680 100668
rect 142616 100608 142680 100612
rect 142696 100668 142760 100672
rect 142696 100612 142700 100668
rect 142700 100612 142756 100668
rect 142756 100612 142760 100668
rect 142696 100608 142760 100612
rect 173176 100668 173240 100672
rect 173176 100612 173180 100668
rect 173180 100612 173236 100668
rect 173236 100612 173240 100668
rect 173176 100608 173240 100612
rect 173256 100668 173320 100672
rect 173256 100612 173260 100668
rect 173260 100612 173316 100668
rect 173316 100612 173320 100668
rect 173256 100608 173320 100612
rect 173336 100668 173400 100672
rect 173336 100612 173340 100668
rect 173340 100612 173396 100668
rect 173396 100612 173400 100668
rect 173336 100608 173400 100612
rect 173416 100668 173480 100672
rect 173416 100612 173420 100668
rect 173420 100612 173476 100668
rect 173476 100612 173480 100668
rect 173416 100608 173480 100612
rect 4216 100124 4280 100128
rect 4216 100068 4220 100124
rect 4220 100068 4276 100124
rect 4276 100068 4280 100124
rect 4216 100064 4280 100068
rect 4296 100124 4360 100128
rect 4296 100068 4300 100124
rect 4300 100068 4356 100124
rect 4356 100068 4360 100124
rect 4296 100064 4360 100068
rect 4376 100124 4440 100128
rect 4376 100068 4380 100124
rect 4380 100068 4436 100124
rect 4436 100068 4440 100124
rect 4376 100064 4440 100068
rect 4456 100124 4520 100128
rect 4456 100068 4460 100124
rect 4460 100068 4516 100124
rect 4516 100068 4520 100124
rect 4456 100064 4520 100068
rect 34936 100124 35000 100128
rect 34936 100068 34940 100124
rect 34940 100068 34996 100124
rect 34996 100068 35000 100124
rect 34936 100064 35000 100068
rect 35016 100124 35080 100128
rect 35016 100068 35020 100124
rect 35020 100068 35076 100124
rect 35076 100068 35080 100124
rect 35016 100064 35080 100068
rect 35096 100124 35160 100128
rect 35096 100068 35100 100124
rect 35100 100068 35156 100124
rect 35156 100068 35160 100124
rect 35096 100064 35160 100068
rect 35176 100124 35240 100128
rect 35176 100068 35180 100124
rect 35180 100068 35236 100124
rect 35236 100068 35240 100124
rect 35176 100064 35240 100068
rect 65656 100124 65720 100128
rect 65656 100068 65660 100124
rect 65660 100068 65716 100124
rect 65716 100068 65720 100124
rect 65656 100064 65720 100068
rect 65736 100124 65800 100128
rect 65736 100068 65740 100124
rect 65740 100068 65796 100124
rect 65796 100068 65800 100124
rect 65736 100064 65800 100068
rect 65816 100124 65880 100128
rect 65816 100068 65820 100124
rect 65820 100068 65876 100124
rect 65876 100068 65880 100124
rect 65816 100064 65880 100068
rect 65896 100124 65960 100128
rect 65896 100068 65900 100124
rect 65900 100068 65956 100124
rect 65956 100068 65960 100124
rect 65896 100064 65960 100068
rect 96376 100124 96440 100128
rect 96376 100068 96380 100124
rect 96380 100068 96436 100124
rect 96436 100068 96440 100124
rect 96376 100064 96440 100068
rect 96456 100124 96520 100128
rect 96456 100068 96460 100124
rect 96460 100068 96516 100124
rect 96516 100068 96520 100124
rect 96456 100064 96520 100068
rect 96536 100124 96600 100128
rect 96536 100068 96540 100124
rect 96540 100068 96596 100124
rect 96596 100068 96600 100124
rect 96536 100064 96600 100068
rect 96616 100124 96680 100128
rect 96616 100068 96620 100124
rect 96620 100068 96676 100124
rect 96676 100068 96680 100124
rect 96616 100064 96680 100068
rect 127096 100124 127160 100128
rect 127096 100068 127100 100124
rect 127100 100068 127156 100124
rect 127156 100068 127160 100124
rect 127096 100064 127160 100068
rect 127176 100124 127240 100128
rect 127176 100068 127180 100124
rect 127180 100068 127236 100124
rect 127236 100068 127240 100124
rect 127176 100064 127240 100068
rect 127256 100124 127320 100128
rect 127256 100068 127260 100124
rect 127260 100068 127316 100124
rect 127316 100068 127320 100124
rect 127256 100064 127320 100068
rect 127336 100124 127400 100128
rect 127336 100068 127340 100124
rect 127340 100068 127396 100124
rect 127396 100068 127400 100124
rect 127336 100064 127400 100068
rect 157816 100124 157880 100128
rect 157816 100068 157820 100124
rect 157820 100068 157876 100124
rect 157876 100068 157880 100124
rect 157816 100064 157880 100068
rect 157896 100124 157960 100128
rect 157896 100068 157900 100124
rect 157900 100068 157956 100124
rect 157956 100068 157960 100124
rect 157896 100064 157960 100068
rect 157976 100124 158040 100128
rect 157976 100068 157980 100124
rect 157980 100068 158036 100124
rect 158036 100068 158040 100124
rect 157976 100064 158040 100068
rect 158056 100124 158120 100128
rect 158056 100068 158060 100124
rect 158060 100068 158116 100124
rect 158116 100068 158120 100124
rect 158056 100064 158120 100068
rect 19576 99580 19640 99584
rect 19576 99524 19580 99580
rect 19580 99524 19636 99580
rect 19636 99524 19640 99580
rect 19576 99520 19640 99524
rect 19656 99580 19720 99584
rect 19656 99524 19660 99580
rect 19660 99524 19716 99580
rect 19716 99524 19720 99580
rect 19656 99520 19720 99524
rect 19736 99580 19800 99584
rect 19736 99524 19740 99580
rect 19740 99524 19796 99580
rect 19796 99524 19800 99580
rect 19736 99520 19800 99524
rect 19816 99580 19880 99584
rect 19816 99524 19820 99580
rect 19820 99524 19876 99580
rect 19876 99524 19880 99580
rect 19816 99520 19880 99524
rect 50296 99580 50360 99584
rect 50296 99524 50300 99580
rect 50300 99524 50356 99580
rect 50356 99524 50360 99580
rect 50296 99520 50360 99524
rect 50376 99580 50440 99584
rect 50376 99524 50380 99580
rect 50380 99524 50436 99580
rect 50436 99524 50440 99580
rect 50376 99520 50440 99524
rect 50456 99580 50520 99584
rect 50456 99524 50460 99580
rect 50460 99524 50516 99580
rect 50516 99524 50520 99580
rect 50456 99520 50520 99524
rect 50536 99580 50600 99584
rect 50536 99524 50540 99580
rect 50540 99524 50596 99580
rect 50596 99524 50600 99580
rect 50536 99520 50600 99524
rect 81016 99580 81080 99584
rect 81016 99524 81020 99580
rect 81020 99524 81076 99580
rect 81076 99524 81080 99580
rect 81016 99520 81080 99524
rect 81096 99580 81160 99584
rect 81096 99524 81100 99580
rect 81100 99524 81156 99580
rect 81156 99524 81160 99580
rect 81096 99520 81160 99524
rect 81176 99580 81240 99584
rect 81176 99524 81180 99580
rect 81180 99524 81236 99580
rect 81236 99524 81240 99580
rect 81176 99520 81240 99524
rect 81256 99580 81320 99584
rect 81256 99524 81260 99580
rect 81260 99524 81316 99580
rect 81316 99524 81320 99580
rect 81256 99520 81320 99524
rect 111736 99580 111800 99584
rect 111736 99524 111740 99580
rect 111740 99524 111796 99580
rect 111796 99524 111800 99580
rect 111736 99520 111800 99524
rect 111816 99580 111880 99584
rect 111816 99524 111820 99580
rect 111820 99524 111876 99580
rect 111876 99524 111880 99580
rect 111816 99520 111880 99524
rect 111896 99580 111960 99584
rect 111896 99524 111900 99580
rect 111900 99524 111956 99580
rect 111956 99524 111960 99580
rect 111896 99520 111960 99524
rect 111976 99580 112040 99584
rect 111976 99524 111980 99580
rect 111980 99524 112036 99580
rect 112036 99524 112040 99580
rect 111976 99520 112040 99524
rect 142456 99580 142520 99584
rect 142456 99524 142460 99580
rect 142460 99524 142516 99580
rect 142516 99524 142520 99580
rect 142456 99520 142520 99524
rect 142536 99580 142600 99584
rect 142536 99524 142540 99580
rect 142540 99524 142596 99580
rect 142596 99524 142600 99580
rect 142536 99520 142600 99524
rect 142616 99580 142680 99584
rect 142616 99524 142620 99580
rect 142620 99524 142676 99580
rect 142676 99524 142680 99580
rect 142616 99520 142680 99524
rect 142696 99580 142760 99584
rect 142696 99524 142700 99580
rect 142700 99524 142756 99580
rect 142756 99524 142760 99580
rect 142696 99520 142760 99524
rect 173176 99580 173240 99584
rect 173176 99524 173180 99580
rect 173180 99524 173236 99580
rect 173236 99524 173240 99580
rect 173176 99520 173240 99524
rect 173256 99580 173320 99584
rect 173256 99524 173260 99580
rect 173260 99524 173316 99580
rect 173316 99524 173320 99580
rect 173256 99520 173320 99524
rect 173336 99580 173400 99584
rect 173336 99524 173340 99580
rect 173340 99524 173396 99580
rect 173396 99524 173400 99580
rect 173336 99520 173400 99524
rect 173416 99580 173480 99584
rect 173416 99524 173420 99580
rect 173420 99524 173476 99580
rect 173476 99524 173480 99580
rect 173416 99520 173480 99524
rect 4216 99036 4280 99040
rect 4216 98980 4220 99036
rect 4220 98980 4276 99036
rect 4276 98980 4280 99036
rect 4216 98976 4280 98980
rect 4296 99036 4360 99040
rect 4296 98980 4300 99036
rect 4300 98980 4356 99036
rect 4356 98980 4360 99036
rect 4296 98976 4360 98980
rect 4376 99036 4440 99040
rect 4376 98980 4380 99036
rect 4380 98980 4436 99036
rect 4436 98980 4440 99036
rect 4376 98976 4440 98980
rect 4456 99036 4520 99040
rect 4456 98980 4460 99036
rect 4460 98980 4516 99036
rect 4516 98980 4520 99036
rect 4456 98976 4520 98980
rect 34936 99036 35000 99040
rect 34936 98980 34940 99036
rect 34940 98980 34996 99036
rect 34996 98980 35000 99036
rect 34936 98976 35000 98980
rect 35016 99036 35080 99040
rect 35016 98980 35020 99036
rect 35020 98980 35076 99036
rect 35076 98980 35080 99036
rect 35016 98976 35080 98980
rect 35096 99036 35160 99040
rect 35096 98980 35100 99036
rect 35100 98980 35156 99036
rect 35156 98980 35160 99036
rect 35096 98976 35160 98980
rect 35176 99036 35240 99040
rect 35176 98980 35180 99036
rect 35180 98980 35236 99036
rect 35236 98980 35240 99036
rect 35176 98976 35240 98980
rect 65656 99036 65720 99040
rect 65656 98980 65660 99036
rect 65660 98980 65716 99036
rect 65716 98980 65720 99036
rect 65656 98976 65720 98980
rect 65736 99036 65800 99040
rect 65736 98980 65740 99036
rect 65740 98980 65796 99036
rect 65796 98980 65800 99036
rect 65736 98976 65800 98980
rect 65816 99036 65880 99040
rect 65816 98980 65820 99036
rect 65820 98980 65876 99036
rect 65876 98980 65880 99036
rect 65816 98976 65880 98980
rect 65896 99036 65960 99040
rect 65896 98980 65900 99036
rect 65900 98980 65956 99036
rect 65956 98980 65960 99036
rect 65896 98976 65960 98980
rect 96376 99036 96440 99040
rect 96376 98980 96380 99036
rect 96380 98980 96436 99036
rect 96436 98980 96440 99036
rect 96376 98976 96440 98980
rect 96456 99036 96520 99040
rect 96456 98980 96460 99036
rect 96460 98980 96516 99036
rect 96516 98980 96520 99036
rect 96456 98976 96520 98980
rect 96536 99036 96600 99040
rect 96536 98980 96540 99036
rect 96540 98980 96596 99036
rect 96596 98980 96600 99036
rect 96536 98976 96600 98980
rect 96616 99036 96680 99040
rect 96616 98980 96620 99036
rect 96620 98980 96676 99036
rect 96676 98980 96680 99036
rect 96616 98976 96680 98980
rect 127096 99036 127160 99040
rect 127096 98980 127100 99036
rect 127100 98980 127156 99036
rect 127156 98980 127160 99036
rect 127096 98976 127160 98980
rect 127176 99036 127240 99040
rect 127176 98980 127180 99036
rect 127180 98980 127236 99036
rect 127236 98980 127240 99036
rect 127176 98976 127240 98980
rect 127256 99036 127320 99040
rect 127256 98980 127260 99036
rect 127260 98980 127316 99036
rect 127316 98980 127320 99036
rect 127256 98976 127320 98980
rect 127336 99036 127400 99040
rect 127336 98980 127340 99036
rect 127340 98980 127396 99036
rect 127396 98980 127400 99036
rect 127336 98976 127400 98980
rect 157816 99036 157880 99040
rect 157816 98980 157820 99036
rect 157820 98980 157876 99036
rect 157876 98980 157880 99036
rect 157816 98976 157880 98980
rect 157896 99036 157960 99040
rect 157896 98980 157900 99036
rect 157900 98980 157956 99036
rect 157956 98980 157960 99036
rect 157896 98976 157960 98980
rect 157976 99036 158040 99040
rect 157976 98980 157980 99036
rect 157980 98980 158036 99036
rect 158036 98980 158040 99036
rect 157976 98976 158040 98980
rect 158056 99036 158120 99040
rect 158056 98980 158060 99036
rect 158060 98980 158116 99036
rect 158116 98980 158120 99036
rect 158056 98976 158120 98980
rect 19576 98492 19640 98496
rect 19576 98436 19580 98492
rect 19580 98436 19636 98492
rect 19636 98436 19640 98492
rect 19576 98432 19640 98436
rect 19656 98492 19720 98496
rect 19656 98436 19660 98492
rect 19660 98436 19716 98492
rect 19716 98436 19720 98492
rect 19656 98432 19720 98436
rect 19736 98492 19800 98496
rect 19736 98436 19740 98492
rect 19740 98436 19796 98492
rect 19796 98436 19800 98492
rect 19736 98432 19800 98436
rect 19816 98492 19880 98496
rect 19816 98436 19820 98492
rect 19820 98436 19876 98492
rect 19876 98436 19880 98492
rect 19816 98432 19880 98436
rect 50296 98492 50360 98496
rect 50296 98436 50300 98492
rect 50300 98436 50356 98492
rect 50356 98436 50360 98492
rect 50296 98432 50360 98436
rect 50376 98492 50440 98496
rect 50376 98436 50380 98492
rect 50380 98436 50436 98492
rect 50436 98436 50440 98492
rect 50376 98432 50440 98436
rect 50456 98492 50520 98496
rect 50456 98436 50460 98492
rect 50460 98436 50516 98492
rect 50516 98436 50520 98492
rect 50456 98432 50520 98436
rect 50536 98492 50600 98496
rect 50536 98436 50540 98492
rect 50540 98436 50596 98492
rect 50596 98436 50600 98492
rect 50536 98432 50600 98436
rect 81016 98492 81080 98496
rect 81016 98436 81020 98492
rect 81020 98436 81076 98492
rect 81076 98436 81080 98492
rect 81016 98432 81080 98436
rect 81096 98492 81160 98496
rect 81096 98436 81100 98492
rect 81100 98436 81156 98492
rect 81156 98436 81160 98492
rect 81096 98432 81160 98436
rect 81176 98492 81240 98496
rect 81176 98436 81180 98492
rect 81180 98436 81236 98492
rect 81236 98436 81240 98492
rect 81176 98432 81240 98436
rect 81256 98492 81320 98496
rect 81256 98436 81260 98492
rect 81260 98436 81316 98492
rect 81316 98436 81320 98492
rect 81256 98432 81320 98436
rect 111736 98492 111800 98496
rect 111736 98436 111740 98492
rect 111740 98436 111796 98492
rect 111796 98436 111800 98492
rect 111736 98432 111800 98436
rect 111816 98492 111880 98496
rect 111816 98436 111820 98492
rect 111820 98436 111876 98492
rect 111876 98436 111880 98492
rect 111816 98432 111880 98436
rect 111896 98492 111960 98496
rect 111896 98436 111900 98492
rect 111900 98436 111956 98492
rect 111956 98436 111960 98492
rect 111896 98432 111960 98436
rect 111976 98492 112040 98496
rect 111976 98436 111980 98492
rect 111980 98436 112036 98492
rect 112036 98436 112040 98492
rect 111976 98432 112040 98436
rect 142456 98492 142520 98496
rect 142456 98436 142460 98492
rect 142460 98436 142516 98492
rect 142516 98436 142520 98492
rect 142456 98432 142520 98436
rect 142536 98492 142600 98496
rect 142536 98436 142540 98492
rect 142540 98436 142596 98492
rect 142596 98436 142600 98492
rect 142536 98432 142600 98436
rect 142616 98492 142680 98496
rect 142616 98436 142620 98492
rect 142620 98436 142676 98492
rect 142676 98436 142680 98492
rect 142616 98432 142680 98436
rect 142696 98492 142760 98496
rect 142696 98436 142700 98492
rect 142700 98436 142756 98492
rect 142756 98436 142760 98492
rect 142696 98432 142760 98436
rect 173176 98492 173240 98496
rect 173176 98436 173180 98492
rect 173180 98436 173236 98492
rect 173236 98436 173240 98492
rect 173176 98432 173240 98436
rect 173256 98492 173320 98496
rect 173256 98436 173260 98492
rect 173260 98436 173316 98492
rect 173316 98436 173320 98492
rect 173256 98432 173320 98436
rect 173336 98492 173400 98496
rect 173336 98436 173340 98492
rect 173340 98436 173396 98492
rect 173396 98436 173400 98492
rect 173336 98432 173400 98436
rect 173416 98492 173480 98496
rect 173416 98436 173420 98492
rect 173420 98436 173476 98492
rect 173476 98436 173480 98492
rect 173416 98432 173480 98436
rect 4216 97948 4280 97952
rect 4216 97892 4220 97948
rect 4220 97892 4276 97948
rect 4276 97892 4280 97948
rect 4216 97888 4280 97892
rect 4296 97948 4360 97952
rect 4296 97892 4300 97948
rect 4300 97892 4356 97948
rect 4356 97892 4360 97948
rect 4296 97888 4360 97892
rect 4376 97948 4440 97952
rect 4376 97892 4380 97948
rect 4380 97892 4436 97948
rect 4436 97892 4440 97948
rect 4376 97888 4440 97892
rect 4456 97948 4520 97952
rect 4456 97892 4460 97948
rect 4460 97892 4516 97948
rect 4516 97892 4520 97948
rect 4456 97888 4520 97892
rect 34936 97948 35000 97952
rect 34936 97892 34940 97948
rect 34940 97892 34996 97948
rect 34996 97892 35000 97948
rect 34936 97888 35000 97892
rect 35016 97948 35080 97952
rect 35016 97892 35020 97948
rect 35020 97892 35076 97948
rect 35076 97892 35080 97948
rect 35016 97888 35080 97892
rect 35096 97948 35160 97952
rect 35096 97892 35100 97948
rect 35100 97892 35156 97948
rect 35156 97892 35160 97948
rect 35096 97888 35160 97892
rect 35176 97948 35240 97952
rect 35176 97892 35180 97948
rect 35180 97892 35236 97948
rect 35236 97892 35240 97948
rect 35176 97888 35240 97892
rect 65656 97948 65720 97952
rect 65656 97892 65660 97948
rect 65660 97892 65716 97948
rect 65716 97892 65720 97948
rect 65656 97888 65720 97892
rect 65736 97948 65800 97952
rect 65736 97892 65740 97948
rect 65740 97892 65796 97948
rect 65796 97892 65800 97948
rect 65736 97888 65800 97892
rect 65816 97948 65880 97952
rect 65816 97892 65820 97948
rect 65820 97892 65876 97948
rect 65876 97892 65880 97948
rect 65816 97888 65880 97892
rect 65896 97948 65960 97952
rect 65896 97892 65900 97948
rect 65900 97892 65956 97948
rect 65956 97892 65960 97948
rect 65896 97888 65960 97892
rect 96376 97948 96440 97952
rect 96376 97892 96380 97948
rect 96380 97892 96436 97948
rect 96436 97892 96440 97948
rect 96376 97888 96440 97892
rect 96456 97948 96520 97952
rect 96456 97892 96460 97948
rect 96460 97892 96516 97948
rect 96516 97892 96520 97948
rect 96456 97888 96520 97892
rect 96536 97948 96600 97952
rect 96536 97892 96540 97948
rect 96540 97892 96596 97948
rect 96596 97892 96600 97948
rect 96536 97888 96600 97892
rect 96616 97948 96680 97952
rect 96616 97892 96620 97948
rect 96620 97892 96676 97948
rect 96676 97892 96680 97948
rect 96616 97888 96680 97892
rect 127096 97948 127160 97952
rect 127096 97892 127100 97948
rect 127100 97892 127156 97948
rect 127156 97892 127160 97948
rect 127096 97888 127160 97892
rect 127176 97948 127240 97952
rect 127176 97892 127180 97948
rect 127180 97892 127236 97948
rect 127236 97892 127240 97948
rect 127176 97888 127240 97892
rect 127256 97948 127320 97952
rect 127256 97892 127260 97948
rect 127260 97892 127316 97948
rect 127316 97892 127320 97948
rect 127256 97888 127320 97892
rect 127336 97948 127400 97952
rect 127336 97892 127340 97948
rect 127340 97892 127396 97948
rect 127396 97892 127400 97948
rect 127336 97888 127400 97892
rect 157816 97948 157880 97952
rect 157816 97892 157820 97948
rect 157820 97892 157876 97948
rect 157876 97892 157880 97948
rect 157816 97888 157880 97892
rect 157896 97948 157960 97952
rect 157896 97892 157900 97948
rect 157900 97892 157956 97948
rect 157956 97892 157960 97948
rect 157896 97888 157960 97892
rect 157976 97948 158040 97952
rect 157976 97892 157980 97948
rect 157980 97892 158036 97948
rect 158036 97892 158040 97948
rect 157976 97888 158040 97892
rect 158056 97948 158120 97952
rect 158056 97892 158060 97948
rect 158060 97892 158116 97948
rect 158116 97892 158120 97948
rect 158056 97888 158120 97892
rect 19576 97404 19640 97408
rect 19576 97348 19580 97404
rect 19580 97348 19636 97404
rect 19636 97348 19640 97404
rect 19576 97344 19640 97348
rect 19656 97404 19720 97408
rect 19656 97348 19660 97404
rect 19660 97348 19716 97404
rect 19716 97348 19720 97404
rect 19656 97344 19720 97348
rect 19736 97404 19800 97408
rect 19736 97348 19740 97404
rect 19740 97348 19796 97404
rect 19796 97348 19800 97404
rect 19736 97344 19800 97348
rect 19816 97404 19880 97408
rect 19816 97348 19820 97404
rect 19820 97348 19876 97404
rect 19876 97348 19880 97404
rect 19816 97344 19880 97348
rect 50296 97404 50360 97408
rect 50296 97348 50300 97404
rect 50300 97348 50356 97404
rect 50356 97348 50360 97404
rect 50296 97344 50360 97348
rect 50376 97404 50440 97408
rect 50376 97348 50380 97404
rect 50380 97348 50436 97404
rect 50436 97348 50440 97404
rect 50376 97344 50440 97348
rect 50456 97404 50520 97408
rect 50456 97348 50460 97404
rect 50460 97348 50516 97404
rect 50516 97348 50520 97404
rect 50456 97344 50520 97348
rect 50536 97404 50600 97408
rect 50536 97348 50540 97404
rect 50540 97348 50596 97404
rect 50596 97348 50600 97404
rect 50536 97344 50600 97348
rect 81016 97404 81080 97408
rect 81016 97348 81020 97404
rect 81020 97348 81076 97404
rect 81076 97348 81080 97404
rect 81016 97344 81080 97348
rect 81096 97404 81160 97408
rect 81096 97348 81100 97404
rect 81100 97348 81156 97404
rect 81156 97348 81160 97404
rect 81096 97344 81160 97348
rect 81176 97404 81240 97408
rect 81176 97348 81180 97404
rect 81180 97348 81236 97404
rect 81236 97348 81240 97404
rect 81176 97344 81240 97348
rect 81256 97404 81320 97408
rect 81256 97348 81260 97404
rect 81260 97348 81316 97404
rect 81316 97348 81320 97404
rect 81256 97344 81320 97348
rect 111736 97404 111800 97408
rect 111736 97348 111740 97404
rect 111740 97348 111796 97404
rect 111796 97348 111800 97404
rect 111736 97344 111800 97348
rect 111816 97404 111880 97408
rect 111816 97348 111820 97404
rect 111820 97348 111876 97404
rect 111876 97348 111880 97404
rect 111816 97344 111880 97348
rect 111896 97404 111960 97408
rect 111896 97348 111900 97404
rect 111900 97348 111956 97404
rect 111956 97348 111960 97404
rect 111896 97344 111960 97348
rect 111976 97404 112040 97408
rect 111976 97348 111980 97404
rect 111980 97348 112036 97404
rect 112036 97348 112040 97404
rect 111976 97344 112040 97348
rect 142456 97404 142520 97408
rect 142456 97348 142460 97404
rect 142460 97348 142516 97404
rect 142516 97348 142520 97404
rect 142456 97344 142520 97348
rect 142536 97404 142600 97408
rect 142536 97348 142540 97404
rect 142540 97348 142596 97404
rect 142596 97348 142600 97404
rect 142536 97344 142600 97348
rect 142616 97404 142680 97408
rect 142616 97348 142620 97404
rect 142620 97348 142676 97404
rect 142676 97348 142680 97404
rect 142616 97344 142680 97348
rect 142696 97404 142760 97408
rect 142696 97348 142700 97404
rect 142700 97348 142756 97404
rect 142756 97348 142760 97404
rect 142696 97344 142760 97348
rect 173176 97404 173240 97408
rect 173176 97348 173180 97404
rect 173180 97348 173236 97404
rect 173236 97348 173240 97404
rect 173176 97344 173240 97348
rect 173256 97404 173320 97408
rect 173256 97348 173260 97404
rect 173260 97348 173316 97404
rect 173316 97348 173320 97404
rect 173256 97344 173320 97348
rect 173336 97404 173400 97408
rect 173336 97348 173340 97404
rect 173340 97348 173396 97404
rect 173396 97348 173400 97404
rect 173336 97344 173400 97348
rect 173416 97404 173480 97408
rect 173416 97348 173420 97404
rect 173420 97348 173476 97404
rect 173476 97348 173480 97404
rect 173416 97344 173480 97348
rect 4216 96860 4280 96864
rect 4216 96804 4220 96860
rect 4220 96804 4276 96860
rect 4276 96804 4280 96860
rect 4216 96800 4280 96804
rect 4296 96860 4360 96864
rect 4296 96804 4300 96860
rect 4300 96804 4356 96860
rect 4356 96804 4360 96860
rect 4296 96800 4360 96804
rect 4376 96860 4440 96864
rect 4376 96804 4380 96860
rect 4380 96804 4436 96860
rect 4436 96804 4440 96860
rect 4376 96800 4440 96804
rect 4456 96860 4520 96864
rect 4456 96804 4460 96860
rect 4460 96804 4516 96860
rect 4516 96804 4520 96860
rect 4456 96800 4520 96804
rect 34936 96860 35000 96864
rect 34936 96804 34940 96860
rect 34940 96804 34996 96860
rect 34996 96804 35000 96860
rect 34936 96800 35000 96804
rect 35016 96860 35080 96864
rect 35016 96804 35020 96860
rect 35020 96804 35076 96860
rect 35076 96804 35080 96860
rect 35016 96800 35080 96804
rect 35096 96860 35160 96864
rect 35096 96804 35100 96860
rect 35100 96804 35156 96860
rect 35156 96804 35160 96860
rect 35096 96800 35160 96804
rect 35176 96860 35240 96864
rect 35176 96804 35180 96860
rect 35180 96804 35236 96860
rect 35236 96804 35240 96860
rect 35176 96800 35240 96804
rect 65656 96860 65720 96864
rect 65656 96804 65660 96860
rect 65660 96804 65716 96860
rect 65716 96804 65720 96860
rect 65656 96800 65720 96804
rect 65736 96860 65800 96864
rect 65736 96804 65740 96860
rect 65740 96804 65796 96860
rect 65796 96804 65800 96860
rect 65736 96800 65800 96804
rect 65816 96860 65880 96864
rect 65816 96804 65820 96860
rect 65820 96804 65876 96860
rect 65876 96804 65880 96860
rect 65816 96800 65880 96804
rect 65896 96860 65960 96864
rect 65896 96804 65900 96860
rect 65900 96804 65956 96860
rect 65956 96804 65960 96860
rect 65896 96800 65960 96804
rect 96376 96860 96440 96864
rect 96376 96804 96380 96860
rect 96380 96804 96436 96860
rect 96436 96804 96440 96860
rect 96376 96800 96440 96804
rect 96456 96860 96520 96864
rect 96456 96804 96460 96860
rect 96460 96804 96516 96860
rect 96516 96804 96520 96860
rect 96456 96800 96520 96804
rect 96536 96860 96600 96864
rect 96536 96804 96540 96860
rect 96540 96804 96596 96860
rect 96596 96804 96600 96860
rect 96536 96800 96600 96804
rect 96616 96860 96680 96864
rect 96616 96804 96620 96860
rect 96620 96804 96676 96860
rect 96676 96804 96680 96860
rect 96616 96800 96680 96804
rect 127096 96860 127160 96864
rect 127096 96804 127100 96860
rect 127100 96804 127156 96860
rect 127156 96804 127160 96860
rect 127096 96800 127160 96804
rect 127176 96860 127240 96864
rect 127176 96804 127180 96860
rect 127180 96804 127236 96860
rect 127236 96804 127240 96860
rect 127176 96800 127240 96804
rect 127256 96860 127320 96864
rect 127256 96804 127260 96860
rect 127260 96804 127316 96860
rect 127316 96804 127320 96860
rect 127256 96800 127320 96804
rect 127336 96860 127400 96864
rect 127336 96804 127340 96860
rect 127340 96804 127396 96860
rect 127396 96804 127400 96860
rect 127336 96800 127400 96804
rect 157816 96860 157880 96864
rect 157816 96804 157820 96860
rect 157820 96804 157876 96860
rect 157876 96804 157880 96860
rect 157816 96800 157880 96804
rect 157896 96860 157960 96864
rect 157896 96804 157900 96860
rect 157900 96804 157956 96860
rect 157956 96804 157960 96860
rect 157896 96800 157960 96804
rect 157976 96860 158040 96864
rect 157976 96804 157980 96860
rect 157980 96804 158036 96860
rect 158036 96804 158040 96860
rect 157976 96800 158040 96804
rect 158056 96860 158120 96864
rect 158056 96804 158060 96860
rect 158060 96804 158116 96860
rect 158116 96804 158120 96860
rect 158056 96800 158120 96804
rect 19576 96316 19640 96320
rect 19576 96260 19580 96316
rect 19580 96260 19636 96316
rect 19636 96260 19640 96316
rect 19576 96256 19640 96260
rect 19656 96316 19720 96320
rect 19656 96260 19660 96316
rect 19660 96260 19716 96316
rect 19716 96260 19720 96316
rect 19656 96256 19720 96260
rect 19736 96316 19800 96320
rect 19736 96260 19740 96316
rect 19740 96260 19796 96316
rect 19796 96260 19800 96316
rect 19736 96256 19800 96260
rect 19816 96316 19880 96320
rect 19816 96260 19820 96316
rect 19820 96260 19876 96316
rect 19876 96260 19880 96316
rect 19816 96256 19880 96260
rect 50296 96316 50360 96320
rect 50296 96260 50300 96316
rect 50300 96260 50356 96316
rect 50356 96260 50360 96316
rect 50296 96256 50360 96260
rect 50376 96316 50440 96320
rect 50376 96260 50380 96316
rect 50380 96260 50436 96316
rect 50436 96260 50440 96316
rect 50376 96256 50440 96260
rect 50456 96316 50520 96320
rect 50456 96260 50460 96316
rect 50460 96260 50516 96316
rect 50516 96260 50520 96316
rect 50456 96256 50520 96260
rect 50536 96316 50600 96320
rect 50536 96260 50540 96316
rect 50540 96260 50596 96316
rect 50596 96260 50600 96316
rect 50536 96256 50600 96260
rect 81016 96316 81080 96320
rect 81016 96260 81020 96316
rect 81020 96260 81076 96316
rect 81076 96260 81080 96316
rect 81016 96256 81080 96260
rect 81096 96316 81160 96320
rect 81096 96260 81100 96316
rect 81100 96260 81156 96316
rect 81156 96260 81160 96316
rect 81096 96256 81160 96260
rect 81176 96316 81240 96320
rect 81176 96260 81180 96316
rect 81180 96260 81236 96316
rect 81236 96260 81240 96316
rect 81176 96256 81240 96260
rect 81256 96316 81320 96320
rect 81256 96260 81260 96316
rect 81260 96260 81316 96316
rect 81316 96260 81320 96316
rect 81256 96256 81320 96260
rect 111736 96316 111800 96320
rect 111736 96260 111740 96316
rect 111740 96260 111796 96316
rect 111796 96260 111800 96316
rect 111736 96256 111800 96260
rect 111816 96316 111880 96320
rect 111816 96260 111820 96316
rect 111820 96260 111876 96316
rect 111876 96260 111880 96316
rect 111816 96256 111880 96260
rect 111896 96316 111960 96320
rect 111896 96260 111900 96316
rect 111900 96260 111956 96316
rect 111956 96260 111960 96316
rect 111896 96256 111960 96260
rect 111976 96316 112040 96320
rect 111976 96260 111980 96316
rect 111980 96260 112036 96316
rect 112036 96260 112040 96316
rect 111976 96256 112040 96260
rect 142456 96316 142520 96320
rect 142456 96260 142460 96316
rect 142460 96260 142516 96316
rect 142516 96260 142520 96316
rect 142456 96256 142520 96260
rect 142536 96316 142600 96320
rect 142536 96260 142540 96316
rect 142540 96260 142596 96316
rect 142596 96260 142600 96316
rect 142536 96256 142600 96260
rect 142616 96316 142680 96320
rect 142616 96260 142620 96316
rect 142620 96260 142676 96316
rect 142676 96260 142680 96316
rect 142616 96256 142680 96260
rect 142696 96316 142760 96320
rect 142696 96260 142700 96316
rect 142700 96260 142756 96316
rect 142756 96260 142760 96316
rect 142696 96256 142760 96260
rect 173176 96316 173240 96320
rect 173176 96260 173180 96316
rect 173180 96260 173236 96316
rect 173236 96260 173240 96316
rect 173176 96256 173240 96260
rect 173256 96316 173320 96320
rect 173256 96260 173260 96316
rect 173260 96260 173316 96316
rect 173316 96260 173320 96316
rect 173256 96256 173320 96260
rect 173336 96316 173400 96320
rect 173336 96260 173340 96316
rect 173340 96260 173396 96316
rect 173396 96260 173400 96316
rect 173336 96256 173400 96260
rect 173416 96316 173480 96320
rect 173416 96260 173420 96316
rect 173420 96260 173476 96316
rect 173476 96260 173480 96316
rect 173416 96256 173480 96260
rect 4216 95772 4280 95776
rect 4216 95716 4220 95772
rect 4220 95716 4276 95772
rect 4276 95716 4280 95772
rect 4216 95712 4280 95716
rect 4296 95772 4360 95776
rect 4296 95716 4300 95772
rect 4300 95716 4356 95772
rect 4356 95716 4360 95772
rect 4296 95712 4360 95716
rect 4376 95772 4440 95776
rect 4376 95716 4380 95772
rect 4380 95716 4436 95772
rect 4436 95716 4440 95772
rect 4376 95712 4440 95716
rect 4456 95772 4520 95776
rect 4456 95716 4460 95772
rect 4460 95716 4516 95772
rect 4516 95716 4520 95772
rect 4456 95712 4520 95716
rect 34936 95772 35000 95776
rect 34936 95716 34940 95772
rect 34940 95716 34996 95772
rect 34996 95716 35000 95772
rect 34936 95712 35000 95716
rect 35016 95772 35080 95776
rect 35016 95716 35020 95772
rect 35020 95716 35076 95772
rect 35076 95716 35080 95772
rect 35016 95712 35080 95716
rect 35096 95772 35160 95776
rect 35096 95716 35100 95772
rect 35100 95716 35156 95772
rect 35156 95716 35160 95772
rect 35096 95712 35160 95716
rect 35176 95772 35240 95776
rect 35176 95716 35180 95772
rect 35180 95716 35236 95772
rect 35236 95716 35240 95772
rect 35176 95712 35240 95716
rect 65656 95772 65720 95776
rect 65656 95716 65660 95772
rect 65660 95716 65716 95772
rect 65716 95716 65720 95772
rect 65656 95712 65720 95716
rect 65736 95772 65800 95776
rect 65736 95716 65740 95772
rect 65740 95716 65796 95772
rect 65796 95716 65800 95772
rect 65736 95712 65800 95716
rect 65816 95772 65880 95776
rect 65816 95716 65820 95772
rect 65820 95716 65876 95772
rect 65876 95716 65880 95772
rect 65816 95712 65880 95716
rect 65896 95772 65960 95776
rect 65896 95716 65900 95772
rect 65900 95716 65956 95772
rect 65956 95716 65960 95772
rect 65896 95712 65960 95716
rect 96376 95772 96440 95776
rect 96376 95716 96380 95772
rect 96380 95716 96436 95772
rect 96436 95716 96440 95772
rect 96376 95712 96440 95716
rect 96456 95772 96520 95776
rect 96456 95716 96460 95772
rect 96460 95716 96516 95772
rect 96516 95716 96520 95772
rect 96456 95712 96520 95716
rect 96536 95772 96600 95776
rect 96536 95716 96540 95772
rect 96540 95716 96596 95772
rect 96596 95716 96600 95772
rect 96536 95712 96600 95716
rect 96616 95772 96680 95776
rect 96616 95716 96620 95772
rect 96620 95716 96676 95772
rect 96676 95716 96680 95772
rect 96616 95712 96680 95716
rect 127096 95772 127160 95776
rect 127096 95716 127100 95772
rect 127100 95716 127156 95772
rect 127156 95716 127160 95772
rect 127096 95712 127160 95716
rect 127176 95772 127240 95776
rect 127176 95716 127180 95772
rect 127180 95716 127236 95772
rect 127236 95716 127240 95772
rect 127176 95712 127240 95716
rect 127256 95772 127320 95776
rect 127256 95716 127260 95772
rect 127260 95716 127316 95772
rect 127316 95716 127320 95772
rect 127256 95712 127320 95716
rect 127336 95772 127400 95776
rect 127336 95716 127340 95772
rect 127340 95716 127396 95772
rect 127396 95716 127400 95772
rect 127336 95712 127400 95716
rect 157816 95772 157880 95776
rect 157816 95716 157820 95772
rect 157820 95716 157876 95772
rect 157876 95716 157880 95772
rect 157816 95712 157880 95716
rect 157896 95772 157960 95776
rect 157896 95716 157900 95772
rect 157900 95716 157956 95772
rect 157956 95716 157960 95772
rect 157896 95712 157960 95716
rect 157976 95772 158040 95776
rect 157976 95716 157980 95772
rect 157980 95716 158036 95772
rect 158036 95716 158040 95772
rect 157976 95712 158040 95716
rect 158056 95772 158120 95776
rect 158056 95716 158060 95772
rect 158060 95716 158116 95772
rect 158116 95716 158120 95772
rect 158056 95712 158120 95716
rect 19576 95228 19640 95232
rect 19576 95172 19580 95228
rect 19580 95172 19636 95228
rect 19636 95172 19640 95228
rect 19576 95168 19640 95172
rect 19656 95228 19720 95232
rect 19656 95172 19660 95228
rect 19660 95172 19716 95228
rect 19716 95172 19720 95228
rect 19656 95168 19720 95172
rect 19736 95228 19800 95232
rect 19736 95172 19740 95228
rect 19740 95172 19796 95228
rect 19796 95172 19800 95228
rect 19736 95168 19800 95172
rect 19816 95228 19880 95232
rect 19816 95172 19820 95228
rect 19820 95172 19876 95228
rect 19876 95172 19880 95228
rect 19816 95168 19880 95172
rect 50296 95228 50360 95232
rect 50296 95172 50300 95228
rect 50300 95172 50356 95228
rect 50356 95172 50360 95228
rect 50296 95168 50360 95172
rect 50376 95228 50440 95232
rect 50376 95172 50380 95228
rect 50380 95172 50436 95228
rect 50436 95172 50440 95228
rect 50376 95168 50440 95172
rect 50456 95228 50520 95232
rect 50456 95172 50460 95228
rect 50460 95172 50516 95228
rect 50516 95172 50520 95228
rect 50456 95168 50520 95172
rect 50536 95228 50600 95232
rect 50536 95172 50540 95228
rect 50540 95172 50596 95228
rect 50596 95172 50600 95228
rect 50536 95168 50600 95172
rect 81016 95228 81080 95232
rect 81016 95172 81020 95228
rect 81020 95172 81076 95228
rect 81076 95172 81080 95228
rect 81016 95168 81080 95172
rect 81096 95228 81160 95232
rect 81096 95172 81100 95228
rect 81100 95172 81156 95228
rect 81156 95172 81160 95228
rect 81096 95168 81160 95172
rect 81176 95228 81240 95232
rect 81176 95172 81180 95228
rect 81180 95172 81236 95228
rect 81236 95172 81240 95228
rect 81176 95168 81240 95172
rect 81256 95228 81320 95232
rect 81256 95172 81260 95228
rect 81260 95172 81316 95228
rect 81316 95172 81320 95228
rect 81256 95168 81320 95172
rect 111736 95228 111800 95232
rect 111736 95172 111740 95228
rect 111740 95172 111796 95228
rect 111796 95172 111800 95228
rect 111736 95168 111800 95172
rect 111816 95228 111880 95232
rect 111816 95172 111820 95228
rect 111820 95172 111876 95228
rect 111876 95172 111880 95228
rect 111816 95168 111880 95172
rect 111896 95228 111960 95232
rect 111896 95172 111900 95228
rect 111900 95172 111956 95228
rect 111956 95172 111960 95228
rect 111896 95168 111960 95172
rect 111976 95228 112040 95232
rect 111976 95172 111980 95228
rect 111980 95172 112036 95228
rect 112036 95172 112040 95228
rect 111976 95168 112040 95172
rect 142456 95228 142520 95232
rect 142456 95172 142460 95228
rect 142460 95172 142516 95228
rect 142516 95172 142520 95228
rect 142456 95168 142520 95172
rect 142536 95228 142600 95232
rect 142536 95172 142540 95228
rect 142540 95172 142596 95228
rect 142596 95172 142600 95228
rect 142536 95168 142600 95172
rect 142616 95228 142680 95232
rect 142616 95172 142620 95228
rect 142620 95172 142676 95228
rect 142676 95172 142680 95228
rect 142616 95168 142680 95172
rect 142696 95228 142760 95232
rect 142696 95172 142700 95228
rect 142700 95172 142756 95228
rect 142756 95172 142760 95228
rect 142696 95168 142760 95172
rect 173176 95228 173240 95232
rect 173176 95172 173180 95228
rect 173180 95172 173236 95228
rect 173236 95172 173240 95228
rect 173176 95168 173240 95172
rect 173256 95228 173320 95232
rect 173256 95172 173260 95228
rect 173260 95172 173316 95228
rect 173316 95172 173320 95228
rect 173256 95168 173320 95172
rect 173336 95228 173400 95232
rect 173336 95172 173340 95228
rect 173340 95172 173396 95228
rect 173396 95172 173400 95228
rect 173336 95168 173400 95172
rect 173416 95228 173480 95232
rect 173416 95172 173420 95228
rect 173420 95172 173476 95228
rect 173476 95172 173480 95228
rect 173416 95168 173480 95172
rect 4216 94684 4280 94688
rect 4216 94628 4220 94684
rect 4220 94628 4276 94684
rect 4276 94628 4280 94684
rect 4216 94624 4280 94628
rect 4296 94684 4360 94688
rect 4296 94628 4300 94684
rect 4300 94628 4356 94684
rect 4356 94628 4360 94684
rect 4296 94624 4360 94628
rect 4376 94684 4440 94688
rect 4376 94628 4380 94684
rect 4380 94628 4436 94684
rect 4436 94628 4440 94684
rect 4376 94624 4440 94628
rect 4456 94684 4520 94688
rect 4456 94628 4460 94684
rect 4460 94628 4516 94684
rect 4516 94628 4520 94684
rect 4456 94624 4520 94628
rect 34936 94684 35000 94688
rect 34936 94628 34940 94684
rect 34940 94628 34996 94684
rect 34996 94628 35000 94684
rect 34936 94624 35000 94628
rect 35016 94684 35080 94688
rect 35016 94628 35020 94684
rect 35020 94628 35076 94684
rect 35076 94628 35080 94684
rect 35016 94624 35080 94628
rect 35096 94684 35160 94688
rect 35096 94628 35100 94684
rect 35100 94628 35156 94684
rect 35156 94628 35160 94684
rect 35096 94624 35160 94628
rect 35176 94684 35240 94688
rect 35176 94628 35180 94684
rect 35180 94628 35236 94684
rect 35236 94628 35240 94684
rect 35176 94624 35240 94628
rect 65656 94684 65720 94688
rect 65656 94628 65660 94684
rect 65660 94628 65716 94684
rect 65716 94628 65720 94684
rect 65656 94624 65720 94628
rect 65736 94684 65800 94688
rect 65736 94628 65740 94684
rect 65740 94628 65796 94684
rect 65796 94628 65800 94684
rect 65736 94624 65800 94628
rect 65816 94684 65880 94688
rect 65816 94628 65820 94684
rect 65820 94628 65876 94684
rect 65876 94628 65880 94684
rect 65816 94624 65880 94628
rect 65896 94684 65960 94688
rect 65896 94628 65900 94684
rect 65900 94628 65956 94684
rect 65956 94628 65960 94684
rect 65896 94624 65960 94628
rect 96376 94684 96440 94688
rect 96376 94628 96380 94684
rect 96380 94628 96436 94684
rect 96436 94628 96440 94684
rect 96376 94624 96440 94628
rect 96456 94684 96520 94688
rect 96456 94628 96460 94684
rect 96460 94628 96516 94684
rect 96516 94628 96520 94684
rect 96456 94624 96520 94628
rect 96536 94684 96600 94688
rect 96536 94628 96540 94684
rect 96540 94628 96596 94684
rect 96596 94628 96600 94684
rect 96536 94624 96600 94628
rect 96616 94684 96680 94688
rect 96616 94628 96620 94684
rect 96620 94628 96676 94684
rect 96676 94628 96680 94684
rect 96616 94624 96680 94628
rect 127096 94684 127160 94688
rect 127096 94628 127100 94684
rect 127100 94628 127156 94684
rect 127156 94628 127160 94684
rect 127096 94624 127160 94628
rect 127176 94684 127240 94688
rect 127176 94628 127180 94684
rect 127180 94628 127236 94684
rect 127236 94628 127240 94684
rect 127176 94624 127240 94628
rect 127256 94684 127320 94688
rect 127256 94628 127260 94684
rect 127260 94628 127316 94684
rect 127316 94628 127320 94684
rect 127256 94624 127320 94628
rect 127336 94684 127400 94688
rect 127336 94628 127340 94684
rect 127340 94628 127396 94684
rect 127396 94628 127400 94684
rect 127336 94624 127400 94628
rect 157816 94684 157880 94688
rect 157816 94628 157820 94684
rect 157820 94628 157876 94684
rect 157876 94628 157880 94684
rect 157816 94624 157880 94628
rect 157896 94684 157960 94688
rect 157896 94628 157900 94684
rect 157900 94628 157956 94684
rect 157956 94628 157960 94684
rect 157896 94624 157960 94628
rect 157976 94684 158040 94688
rect 157976 94628 157980 94684
rect 157980 94628 158036 94684
rect 158036 94628 158040 94684
rect 157976 94624 158040 94628
rect 158056 94684 158120 94688
rect 158056 94628 158060 94684
rect 158060 94628 158116 94684
rect 158116 94628 158120 94684
rect 158056 94624 158120 94628
rect 19576 94140 19640 94144
rect 19576 94084 19580 94140
rect 19580 94084 19636 94140
rect 19636 94084 19640 94140
rect 19576 94080 19640 94084
rect 19656 94140 19720 94144
rect 19656 94084 19660 94140
rect 19660 94084 19716 94140
rect 19716 94084 19720 94140
rect 19656 94080 19720 94084
rect 19736 94140 19800 94144
rect 19736 94084 19740 94140
rect 19740 94084 19796 94140
rect 19796 94084 19800 94140
rect 19736 94080 19800 94084
rect 19816 94140 19880 94144
rect 19816 94084 19820 94140
rect 19820 94084 19876 94140
rect 19876 94084 19880 94140
rect 19816 94080 19880 94084
rect 50296 94140 50360 94144
rect 50296 94084 50300 94140
rect 50300 94084 50356 94140
rect 50356 94084 50360 94140
rect 50296 94080 50360 94084
rect 50376 94140 50440 94144
rect 50376 94084 50380 94140
rect 50380 94084 50436 94140
rect 50436 94084 50440 94140
rect 50376 94080 50440 94084
rect 50456 94140 50520 94144
rect 50456 94084 50460 94140
rect 50460 94084 50516 94140
rect 50516 94084 50520 94140
rect 50456 94080 50520 94084
rect 50536 94140 50600 94144
rect 50536 94084 50540 94140
rect 50540 94084 50596 94140
rect 50596 94084 50600 94140
rect 50536 94080 50600 94084
rect 81016 94140 81080 94144
rect 81016 94084 81020 94140
rect 81020 94084 81076 94140
rect 81076 94084 81080 94140
rect 81016 94080 81080 94084
rect 81096 94140 81160 94144
rect 81096 94084 81100 94140
rect 81100 94084 81156 94140
rect 81156 94084 81160 94140
rect 81096 94080 81160 94084
rect 81176 94140 81240 94144
rect 81176 94084 81180 94140
rect 81180 94084 81236 94140
rect 81236 94084 81240 94140
rect 81176 94080 81240 94084
rect 81256 94140 81320 94144
rect 81256 94084 81260 94140
rect 81260 94084 81316 94140
rect 81316 94084 81320 94140
rect 81256 94080 81320 94084
rect 111736 94140 111800 94144
rect 111736 94084 111740 94140
rect 111740 94084 111796 94140
rect 111796 94084 111800 94140
rect 111736 94080 111800 94084
rect 111816 94140 111880 94144
rect 111816 94084 111820 94140
rect 111820 94084 111876 94140
rect 111876 94084 111880 94140
rect 111816 94080 111880 94084
rect 111896 94140 111960 94144
rect 111896 94084 111900 94140
rect 111900 94084 111956 94140
rect 111956 94084 111960 94140
rect 111896 94080 111960 94084
rect 111976 94140 112040 94144
rect 111976 94084 111980 94140
rect 111980 94084 112036 94140
rect 112036 94084 112040 94140
rect 111976 94080 112040 94084
rect 142456 94140 142520 94144
rect 142456 94084 142460 94140
rect 142460 94084 142516 94140
rect 142516 94084 142520 94140
rect 142456 94080 142520 94084
rect 142536 94140 142600 94144
rect 142536 94084 142540 94140
rect 142540 94084 142596 94140
rect 142596 94084 142600 94140
rect 142536 94080 142600 94084
rect 142616 94140 142680 94144
rect 142616 94084 142620 94140
rect 142620 94084 142676 94140
rect 142676 94084 142680 94140
rect 142616 94080 142680 94084
rect 142696 94140 142760 94144
rect 142696 94084 142700 94140
rect 142700 94084 142756 94140
rect 142756 94084 142760 94140
rect 142696 94080 142760 94084
rect 173176 94140 173240 94144
rect 173176 94084 173180 94140
rect 173180 94084 173236 94140
rect 173236 94084 173240 94140
rect 173176 94080 173240 94084
rect 173256 94140 173320 94144
rect 173256 94084 173260 94140
rect 173260 94084 173316 94140
rect 173316 94084 173320 94140
rect 173256 94080 173320 94084
rect 173336 94140 173400 94144
rect 173336 94084 173340 94140
rect 173340 94084 173396 94140
rect 173396 94084 173400 94140
rect 173336 94080 173400 94084
rect 173416 94140 173480 94144
rect 173416 94084 173420 94140
rect 173420 94084 173476 94140
rect 173476 94084 173480 94140
rect 173416 94080 173480 94084
rect 4216 93596 4280 93600
rect 4216 93540 4220 93596
rect 4220 93540 4276 93596
rect 4276 93540 4280 93596
rect 4216 93536 4280 93540
rect 4296 93596 4360 93600
rect 4296 93540 4300 93596
rect 4300 93540 4356 93596
rect 4356 93540 4360 93596
rect 4296 93536 4360 93540
rect 4376 93596 4440 93600
rect 4376 93540 4380 93596
rect 4380 93540 4436 93596
rect 4436 93540 4440 93596
rect 4376 93536 4440 93540
rect 4456 93596 4520 93600
rect 4456 93540 4460 93596
rect 4460 93540 4516 93596
rect 4516 93540 4520 93596
rect 4456 93536 4520 93540
rect 34936 93596 35000 93600
rect 34936 93540 34940 93596
rect 34940 93540 34996 93596
rect 34996 93540 35000 93596
rect 34936 93536 35000 93540
rect 35016 93596 35080 93600
rect 35016 93540 35020 93596
rect 35020 93540 35076 93596
rect 35076 93540 35080 93596
rect 35016 93536 35080 93540
rect 35096 93596 35160 93600
rect 35096 93540 35100 93596
rect 35100 93540 35156 93596
rect 35156 93540 35160 93596
rect 35096 93536 35160 93540
rect 35176 93596 35240 93600
rect 35176 93540 35180 93596
rect 35180 93540 35236 93596
rect 35236 93540 35240 93596
rect 35176 93536 35240 93540
rect 65656 93596 65720 93600
rect 65656 93540 65660 93596
rect 65660 93540 65716 93596
rect 65716 93540 65720 93596
rect 65656 93536 65720 93540
rect 65736 93596 65800 93600
rect 65736 93540 65740 93596
rect 65740 93540 65796 93596
rect 65796 93540 65800 93596
rect 65736 93536 65800 93540
rect 65816 93596 65880 93600
rect 65816 93540 65820 93596
rect 65820 93540 65876 93596
rect 65876 93540 65880 93596
rect 65816 93536 65880 93540
rect 65896 93596 65960 93600
rect 65896 93540 65900 93596
rect 65900 93540 65956 93596
rect 65956 93540 65960 93596
rect 65896 93536 65960 93540
rect 96376 93596 96440 93600
rect 96376 93540 96380 93596
rect 96380 93540 96436 93596
rect 96436 93540 96440 93596
rect 96376 93536 96440 93540
rect 96456 93596 96520 93600
rect 96456 93540 96460 93596
rect 96460 93540 96516 93596
rect 96516 93540 96520 93596
rect 96456 93536 96520 93540
rect 96536 93596 96600 93600
rect 96536 93540 96540 93596
rect 96540 93540 96596 93596
rect 96596 93540 96600 93596
rect 96536 93536 96600 93540
rect 96616 93596 96680 93600
rect 96616 93540 96620 93596
rect 96620 93540 96676 93596
rect 96676 93540 96680 93596
rect 96616 93536 96680 93540
rect 127096 93596 127160 93600
rect 127096 93540 127100 93596
rect 127100 93540 127156 93596
rect 127156 93540 127160 93596
rect 127096 93536 127160 93540
rect 127176 93596 127240 93600
rect 127176 93540 127180 93596
rect 127180 93540 127236 93596
rect 127236 93540 127240 93596
rect 127176 93536 127240 93540
rect 127256 93596 127320 93600
rect 127256 93540 127260 93596
rect 127260 93540 127316 93596
rect 127316 93540 127320 93596
rect 127256 93536 127320 93540
rect 127336 93596 127400 93600
rect 127336 93540 127340 93596
rect 127340 93540 127396 93596
rect 127396 93540 127400 93596
rect 127336 93536 127400 93540
rect 157816 93596 157880 93600
rect 157816 93540 157820 93596
rect 157820 93540 157876 93596
rect 157876 93540 157880 93596
rect 157816 93536 157880 93540
rect 157896 93596 157960 93600
rect 157896 93540 157900 93596
rect 157900 93540 157956 93596
rect 157956 93540 157960 93596
rect 157896 93536 157960 93540
rect 157976 93596 158040 93600
rect 157976 93540 157980 93596
rect 157980 93540 158036 93596
rect 158036 93540 158040 93596
rect 157976 93536 158040 93540
rect 158056 93596 158120 93600
rect 158056 93540 158060 93596
rect 158060 93540 158116 93596
rect 158116 93540 158120 93596
rect 158056 93536 158120 93540
rect 19576 93052 19640 93056
rect 19576 92996 19580 93052
rect 19580 92996 19636 93052
rect 19636 92996 19640 93052
rect 19576 92992 19640 92996
rect 19656 93052 19720 93056
rect 19656 92996 19660 93052
rect 19660 92996 19716 93052
rect 19716 92996 19720 93052
rect 19656 92992 19720 92996
rect 19736 93052 19800 93056
rect 19736 92996 19740 93052
rect 19740 92996 19796 93052
rect 19796 92996 19800 93052
rect 19736 92992 19800 92996
rect 19816 93052 19880 93056
rect 19816 92996 19820 93052
rect 19820 92996 19876 93052
rect 19876 92996 19880 93052
rect 19816 92992 19880 92996
rect 50296 93052 50360 93056
rect 50296 92996 50300 93052
rect 50300 92996 50356 93052
rect 50356 92996 50360 93052
rect 50296 92992 50360 92996
rect 50376 93052 50440 93056
rect 50376 92996 50380 93052
rect 50380 92996 50436 93052
rect 50436 92996 50440 93052
rect 50376 92992 50440 92996
rect 50456 93052 50520 93056
rect 50456 92996 50460 93052
rect 50460 92996 50516 93052
rect 50516 92996 50520 93052
rect 50456 92992 50520 92996
rect 50536 93052 50600 93056
rect 50536 92996 50540 93052
rect 50540 92996 50596 93052
rect 50596 92996 50600 93052
rect 50536 92992 50600 92996
rect 81016 93052 81080 93056
rect 81016 92996 81020 93052
rect 81020 92996 81076 93052
rect 81076 92996 81080 93052
rect 81016 92992 81080 92996
rect 81096 93052 81160 93056
rect 81096 92996 81100 93052
rect 81100 92996 81156 93052
rect 81156 92996 81160 93052
rect 81096 92992 81160 92996
rect 81176 93052 81240 93056
rect 81176 92996 81180 93052
rect 81180 92996 81236 93052
rect 81236 92996 81240 93052
rect 81176 92992 81240 92996
rect 81256 93052 81320 93056
rect 81256 92996 81260 93052
rect 81260 92996 81316 93052
rect 81316 92996 81320 93052
rect 81256 92992 81320 92996
rect 111736 93052 111800 93056
rect 111736 92996 111740 93052
rect 111740 92996 111796 93052
rect 111796 92996 111800 93052
rect 111736 92992 111800 92996
rect 111816 93052 111880 93056
rect 111816 92996 111820 93052
rect 111820 92996 111876 93052
rect 111876 92996 111880 93052
rect 111816 92992 111880 92996
rect 111896 93052 111960 93056
rect 111896 92996 111900 93052
rect 111900 92996 111956 93052
rect 111956 92996 111960 93052
rect 111896 92992 111960 92996
rect 111976 93052 112040 93056
rect 111976 92996 111980 93052
rect 111980 92996 112036 93052
rect 112036 92996 112040 93052
rect 111976 92992 112040 92996
rect 142456 93052 142520 93056
rect 142456 92996 142460 93052
rect 142460 92996 142516 93052
rect 142516 92996 142520 93052
rect 142456 92992 142520 92996
rect 142536 93052 142600 93056
rect 142536 92996 142540 93052
rect 142540 92996 142596 93052
rect 142596 92996 142600 93052
rect 142536 92992 142600 92996
rect 142616 93052 142680 93056
rect 142616 92996 142620 93052
rect 142620 92996 142676 93052
rect 142676 92996 142680 93052
rect 142616 92992 142680 92996
rect 142696 93052 142760 93056
rect 142696 92996 142700 93052
rect 142700 92996 142756 93052
rect 142756 92996 142760 93052
rect 142696 92992 142760 92996
rect 173176 93052 173240 93056
rect 173176 92996 173180 93052
rect 173180 92996 173236 93052
rect 173236 92996 173240 93052
rect 173176 92992 173240 92996
rect 173256 93052 173320 93056
rect 173256 92996 173260 93052
rect 173260 92996 173316 93052
rect 173316 92996 173320 93052
rect 173256 92992 173320 92996
rect 173336 93052 173400 93056
rect 173336 92996 173340 93052
rect 173340 92996 173396 93052
rect 173396 92996 173400 93052
rect 173336 92992 173400 92996
rect 173416 93052 173480 93056
rect 173416 92996 173420 93052
rect 173420 92996 173476 93052
rect 173476 92996 173480 93052
rect 173416 92992 173480 92996
rect 4216 92508 4280 92512
rect 4216 92452 4220 92508
rect 4220 92452 4276 92508
rect 4276 92452 4280 92508
rect 4216 92448 4280 92452
rect 4296 92508 4360 92512
rect 4296 92452 4300 92508
rect 4300 92452 4356 92508
rect 4356 92452 4360 92508
rect 4296 92448 4360 92452
rect 4376 92508 4440 92512
rect 4376 92452 4380 92508
rect 4380 92452 4436 92508
rect 4436 92452 4440 92508
rect 4376 92448 4440 92452
rect 4456 92508 4520 92512
rect 4456 92452 4460 92508
rect 4460 92452 4516 92508
rect 4516 92452 4520 92508
rect 4456 92448 4520 92452
rect 34936 92508 35000 92512
rect 34936 92452 34940 92508
rect 34940 92452 34996 92508
rect 34996 92452 35000 92508
rect 34936 92448 35000 92452
rect 35016 92508 35080 92512
rect 35016 92452 35020 92508
rect 35020 92452 35076 92508
rect 35076 92452 35080 92508
rect 35016 92448 35080 92452
rect 35096 92508 35160 92512
rect 35096 92452 35100 92508
rect 35100 92452 35156 92508
rect 35156 92452 35160 92508
rect 35096 92448 35160 92452
rect 35176 92508 35240 92512
rect 35176 92452 35180 92508
rect 35180 92452 35236 92508
rect 35236 92452 35240 92508
rect 35176 92448 35240 92452
rect 65656 92508 65720 92512
rect 65656 92452 65660 92508
rect 65660 92452 65716 92508
rect 65716 92452 65720 92508
rect 65656 92448 65720 92452
rect 65736 92508 65800 92512
rect 65736 92452 65740 92508
rect 65740 92452 65796 92508
rect 65796 92452 65800 92508
rect 65736 92448 65800 92452
rect 65816 92508 65880 92512
rect 65816 92452 65820 92508
rect 65820 92452 65876 92508
rect 65876 92452 65880 92508
rect 65816 92448 65880 92452
rect 65896 92508 65960 92512
rect 65896 92452 65900 92508
rect 65900 92452 65956 92508
rect 65956 92452 65960 92508
rect 65896 92448 65960 92452
rect 96376 92508 96440 92512
rect 96376 92452 96380 92508
rect 96380 92452 96436 92508
rect 96436 92452 96440 92508
rect 96376 92448 96440 92452
rect 96456 92508 96520 92512
rect 96456 92452 96460 92508
rect 96460 92452 96516 92508
rect 96516 92452 96520 92508
rect 96456 92448 96520 92452
rect 96536 92508 96600 92512
rect 96536 92452 96540 92508
rect 96540 92452 96596 92508
rect 96596 92452 96600 92508
rect 96536 92448 96600 92452
rect 96616 92508 96680 92512
rect 96616 92452 96620 92508
rect 96620 92452 96676 92508
rect 96676 92452 96680 92508
rect 96616 92448 96680 92452
rect 127096 92508 127160 92512
rect 127096 92452 127100 92508
rect 127100 92452 127156 92508
rect 127156 92452 127160 92508
rect 127096 92448 127160 92452
rect 127176 92508 127240 92512
rect 127176 92452 127180 92508
rect 127180 92452 127236 92508
rect 127236 92452 127240 92508
rect 127176 92448 127240 92452
rect 127256 92508 127320 92512
rect 127256 92452 127260 92508
rect 127260 92452 127316 92508
rect 127316 92452 127320 92508
rect 127256 92448 127320 92452
rect 127336 92508 127400 92512
rect 127336 92452 127340 92508
rect 127340 92452 127396 92508
rect 127396 92452 127400 92508
rect 127336 92448 127400 92452
rect 157816 92508 157880 92512
rect 157816 92452 157820 92508
rect 157820 92452 157876 92508
rect 157876 92452 157880 92508
rect 157816 92448 157880 92452
rect 157896 92508 157960 92512
rect 157896 92452 157900 92508
rect 157900 92452 157956 92508
rect 157956 92452 157960 92508
rect 157896 92448 157960 92452
rect 157976 92508 158040 92512
rect 157976 92452 157980 92508
rect 157980 92452 158036 92508
rect 158036 92452 158040 92508
rect 157976 92448 158040 92452
rect 158056 92508 158120 92512
rect 158056 92452 158060 92508
rect 158060 92452 158116 92508
rect 158116 92452 158120 92508
rect 158056 92448 158120 92452
rect 19576 91964 19640 91968
rect 19576 91908 19580 91964
rect 19580 91908 19636 91964
rect 19636 91908 19640 91964
rect 19576 91904 19640 91908
rect 19656 91964 19720 91968
rect 19656 91908 19660 91964
rect 19660 91908 19716 91964
rect 19716 91908 19720 91964
rect 19656 91904 19720 91908
rect 19736 91964 19800 91968
rect 19736 91908 19740 91964
rect 19740 91908 19796 91964
rect 19796 91908 19800 91964
rect 19736 91904 19800 91908
rect 19816 91964 19880 91968
rect 19816 91908 19820 91964
rect 19820 91908 19876 91964
rect 19876 91908 19880 91964
rect 19816 91904 19880 91908
rect 50296 91964 50360 91968
rect 50296 91908 50300 91964
rect 50300 91908 50356 91964
rect 50356 91908 50360 91964
rect 50296 91904 50360 91908
rect 50376 91964 50440 91968
rect 50376 91908 50380 91964
rect 50380 91908 50436 91964
rect 50436 91908 50440 91964
rect 50376 91904 50440 91908
rect 50456 91964 50520 91968
rect 50456 91908 50460 91964
rect 50460 91908 50516 91964
rect 50516 91908 50520 91964
rect 50456 91904 50520 91908
rect 50536 91964 50600 91968
rect 50536 91908 50540 91964
rect 50540 91908 50596 91964
rect 50596 91908 50600 91964
rect 50536 91904 50600 91908
rect 81016 91964 81080 91968
rect 81016 91908 81020 91964
rect 81020 91908 81076 91964
rect 81076 91908 81080 91964
rect 81016 91904 81080 91908
rect 81096 91964 81160 91968
rect 81096 91908 81100 91964
rect 81100 91908 81156 91964
rect 81156 91908 81160 91964
rect 81096 91904 81160 91908
rect 81176 91964 81240 91968
rect 81176 91908 81180 91964
rect 81180 91908 81236 91964
rect 81236 91908 81240 91964
rect 81176 91904 81240 91908
rect 81256 91964 81320 91968
rect 81256 91908 81260 91964
rect 81260 91908 81316 91964
rect 81316 91908 81320 91964
rect 81256 91904 81320 91908
rect 111736 91964 111800 91968
rect 111736 91908 111740 91964
rect 111740 91908 111796 91964
rect 111796 91908 111800 91964
rect 111736 91904 111800 91908
rect 111816 91964 111880 91968
rect 111816 91908 111820 91964
rect 111820 91908 111876 91964
rect 111876 91908 111880 91964
rect 111816 91904 111880 91908
rect 111896 91964 111960 91968
rect 111896 91908 111900 91964
rect 111900 91908 111956 91964
rect 111956 91908 111960 91964
rect 111896 91904 111960 91908
rect 111976 91964 112040 91968
rect 111976 91908 111980 91964
rect 111980 91908 112036 91964
rect 112036 91908 112040 91964
rect 111976 91904 112040 91908
rect 142456 91964 142520 91968
rect 142456 91908 142460 91964
rect 142460 91908 142516 91964
rect 142516 91908 142520 91964
rect 142456 91904 142520 91908
rect 142536 91964 142600 91968
rect 142536 91908 142540 91964
rect 142540 91908 142596 91964
rect 142596 91908 142600 91964
rect 142536 91904 142600 91908
rect 142616 91964 142680 91968
rect 142616 91908 142620 91964
rect 142620 91908 142676 91964
rect 142676 91908 142680 91964
rect 142616 91904 142680 91908
rect 142696 91964 142760 91968
rect 142696 91908 142700 91964
rect 142700 91908 142756 91964
rect 142756 91908 142760 91964
rect 142696 91904 142760 91908
rect 173176 91964 173240 91968
rect 173176 91908 173180 91964
rect 173180 91908 173236 91964
rect 173236 91908 173240 91964
rect 173176 91904 173240 91908
rect 173256 91964 173320 91968
rect 173256 91908 173260 91964
rect 173260 91908 173316 91964
rect 173316 91908 173320 91964
rect 173256 91904 173320 91908
rect 173336 91964 173400 91968
rect 173336 91908 173340 91964
rect 173340 91908 173396 91964
rect 173396 91908 173400 91964
rect 173336 91904 173400 91908
rect 173416 91964 173480 91968
rect 173416 91908 173420 91964
rect 173420 91908 173476 91964
rect 173476 91908 173480 91964
rect 173416 91904 173480 91908
rect 4216 91420 4280 91424
rect 4216 91364 4220 91420
rect 4220 91364 4276 91420
rect 4276 91364 4280 91420
rect 4216 91360 4280 91364
rect 4296 91420 4360 91424
rect 4296 91364 4300 91420
rect 4300 91364 4356 91420
rect 4356 91364 4360 91420
rect 4296 91360 4360 91364
rect 4376 91420 4440 91424
rect 4376 91364 4380 91420
rect 4380 91364 4436 91420
rect 4436 91364 4440 91420
rect 4376 91360 4440 91364
rect 4456 91420 4520 91424
rect 4456 91364 4460 91420
rect 4460 91364 4516 91420
rect 4516 91364 4520 91420
rect 4456 91360 4520 91364
rect 34936 91420 35000 91424
rect 34936 91364 34940 91420
rect 34940 91364 34996 91420
rect 34996 91364 35000 91420
rect 34936 91360 35000 91364
rect 35016 91420 35080 91424
rect 35016 91364 35020 91420
rect 35020 91364 35076 91420
rect 35076 91364 35080 91420
rect 35016 91360 35080 91364
rect 35096 91420 35160 91424
rect 35096 91364 35100 91420
rect 35100 91364 35156 91420
rect 35156 91364 35160 91420
rect 35096 91360 35160 91364
rect 35176 91420 35240 91424
rect 35176 91364 35180 91420
rect 35180 91364 35236 91420
rect 35236 91364 35240 91420
rect 35176 91360 35240 91364
rect 65656 91420 65720 91424
rect 65656 91364 65660 91420
rect 65660 91364 65716 91420
rect 65716 91364 65720 91420
rect 65656 91360 65720 91364
rect 65736 91420 65800 91424
rect 65736 91364 65740 91420
rect 65740 91364 65796 91420
rect 65796 91364 65800 91420
rect 65736 91360 65800 91364
rect 65816 91420 65880 91424
rect 65816 91364 65820 91420
rect 65820 91364 65876 91420
rect 65876 91364 65880 91420
rect 65816 91360 65880 91364
rect 65896 91420 65960 91424
rect 65896 91364 65900 91420
rect 65900 91364 65956 91420
rect 65956 91364 65960 91420
rect 65896 91360 65960 91364
rect 96376 91420 96440 91424
rect 96376 91364 96380 91420
rect 96380 91364 96436 91420
rect 96436 91364 96440 91420
rect 96376 91360 96440 91364
rect 96456 91420 96520 91424
rect 96456 91364 96460 91420
rect 96460 91364 96516 91420
rect 96516 91364 96520 91420
rect 96456 91360 96520 91364
rect 96536 91420 96600 91424
rect 96536 91364 96540 91420
rect 96540 91364 96596 91420
rect 96596 91364 96600 91420
rect 96536 91360 96600 91364
rect 96616 91420 96680 91424
rect 96616 91364 96620 91420
rect 96620 91364 96676 91420
rect 96676 91364 96680 91420
rect 96616 91360 96680 91364
rect 127096 91420 127160 91424
rect 127096 91364 127100 91420
rect 127100 91364 127156 91420
rect 127156 91364 127160 91420
rect 127096 91360 127160 91364
rect 127176 91420 127240 91424
rect 127176 91364 127180 91420
rect 127180 91364 127236 91420
rect 127236 91364 127240 91420
rect 127176 91360 127240 91364
rect 127256 91420 127320 91424
rect 127256 91364 127260 91420
rect 127260 91364 127316 91420
rect 127316 91364 127320 91420
rect 127256 91360 127320 91364
rect 127336 91420 127400 91424
rect 127336 91364 127340 91420
rect 127340 91364 127396 91420
rect 127396 91364 127400 91420
rect 127336 91360 127400 91364
rect 157816 91420 157880 91424
rect 157816 91364 157820 91420
rect 157820 91364 157876 91420
rect 157876 91364 157880 91420
rect 157816 91360 157880 91364
rect 157896 91420 157960 91424
rect 157896 91364 157900 91420
rect 157900 91364 157956 91420
rect 157956 91364 157960 91420
rect 157896 91360 157960 91364
rect 157976 91420 158040 91424
rect 157976 91364 157980 91420
rect 157980 91364 158036 91420
rect 158036 91364 158040 91420
rect 157976 91360 158040 91364
rect 158056 91420 158120 91424
rect 158056 91364 158060 91420
rect 158060 91364 158116 91420
rect 158116 91364 158120 91420
rect 158056 91360 158120 91364
rect 19576 90876 19640 90880
rect 19576 90820 19580 90876
rect 19580 90820 19636 90876
rect 19636 90820 19640 90876
rect 19576 90816 19640 90820
rect 19656 90876 19720 90880
rect 19656 90820 19660 90876
rect 19660 90820 19716 90876
rect 19716 90820 19720 90876
rect 19656 90816 19720 90820
rect 19736 90876 19800 90880
rect 19736 90820 19740 90876
rect 19740 90820 19796 90876
rect 19796 90820 19800 90876
rect 19736 90816 19800 90820
rect 19816 90876 19880 90880
rect 19816 90820 19820 90876
rect 19820 90820 19876 90876
rect 19876 90820 19880 90876
rect 19816 90816 19880 90820
rect 50296 90876 50360 90880
rect 50296 90820 50300 90876
rect 50300 90820 50356 90876
rect 50356 90820 50360 90876
rect 50296 90816 50360 90820
rect 50376 90876 50440 90880
rect 50376 90820 50380 90876
rect 50380 90820 50436 90876
rect 50436 90820 50440 90876
rect 50376 90816 50440 90820
rect 50456 90876 50520 90880
rect 50456 90820 50460 90876
rect 50460 90820 50516 90876
rect 50516 90820 50520 90876
rect 50456 90816 50520 90820
rect 50536 90876 50600 90880
rect 50536 90820 50540 90876
rect 50540 90820 50596 90876
rect 50596 90820 50600 90876
rect 50536 90816 50600 90820
rect 81016 90876 81080 90880
rect 81016 90820 81020 90876
rect 81020 90820 81076 90876
rect 81076 90820 81080 90876
rect 81016 90816 81080 90820
rect 81096 90876 81160 90880
rect 81096 90820 81100 90876
rect 81100 90820 81156 90876
rect 81156 90820 81160 90876
rect 81096 90816 81160 90820
rect 81176 90876 81240 90880
rect 81176 90820 81180 90876
rect 81180 90820 81236 90876
rect 81236 90820 81240 90876
rect 81176 90816 81240 90820
rect 81256 90876 81320 90880
rect 81256 90820 81260 90876
rect 81260 90820 81316 90876
rect 81316 90820 81320 90876
rect 81256 90816 81320 90820
rect 111736 90876 111800 90880
rect 111736 90820 111740 90876
rect 111740 90820 111796 90876
rect 111796 90820 111800 90876
rect 111736 90816 111800 90820
rect 111816 90876 111880 90880
rect 111816 90820 111820 90876
rect 111820 90820 111876 90876
rect 111876 90820 111880 90876
rect 111816 90816 111880 90820
rect 111896 90876 111960 90880
rect 111896 90820 111900 90876
rect 111900 90820 111956 90876
rect 111956 90820 111960 90876
rect 111896 90816 111960 90820
rect 111976 90876 112040 90880
rect 111976 90820 111980 90876
rect 111980 90820 112036 90876
rect 112036 90820 112040 90876
rect 111976 90816 112040 90820
rect 142456 90876 142520 90880
rect 142456 90820 142460 90876
rect 142460 90820 142516 90876
rect 142516 90820 142520 90876
rect 142456 90816 142520 90820
rect 142536 90876 142600 90880
rect 142536 90820 142540 90876
rect 142540 90820 142596 90876
rect 142596 90820 142600 90876
rect 142536 90816 142600 90820
rect 142616 90876 142680 90880
rect 142616 90820 142620 90876
rect 142620 90820 142676 90876
rect 142676 90820 142680 90876
rect 142616 90816 142680 90820
rect 142696 90876 142760 90880
rect 142696 90820 142700 90876
rect 142700 90820 142756 90876
rect 142756 90820 142760 90876
rect 142696 90816 142760 90820
rect 173176 90876 173240 90880
rect 173176 90820 173180 90876
rect 173180 90820 173236 90876
rect 173236 90820 173240 90876
rect 173176 90816 173240 90820
rect 173256 90876 173320 90880
rect 173256 90820 173260 90876
rect 173260 90820 173316 90876
rect 173316 90820 173320 90876
rect 173256 90816 173320 90820
rect 173336 90876 173400 90880
rect 173336 90820 173340 90876
rect 173340 90820 173396 90876
rect 173396 90820 173400 90876
rect 173336 90816 173400 90820
rect 173416 90876 173480 90880
rect 173416 90820 173420 90876
rect 173420 90820 173476 90876
rect 173476 90820 173480 90876
rect 173416 90816 173480 90820
rect 4216 90332 4280 90336
rect 4216 90276 4220 90332
rect 4220 90276 4276 90332
rect 4276 90276 4280 90332
rect 4216 90272 4280 90276
rect 4296 90332 4360 90336
rect 4296 90276 4300 90332
rect 4300 90276 4356 90332
rect 4356 90276 4360 90332
rect 4296 90272 4360 90276
rect 4376 90332 4440 90336
rect 4376 90276 4380 90332
rect 4380 90276 4436 90332
rect 4436 90276 4440 90332
rect 4376 90272 4440 90276
rect 4456 90332 4520 90336
rect 4456 90276 4460 90332
rect 4460 90276 4516 90332
rect 4516 90276 4520 90332
rect 4456 90272 4520 90276
rect 34936 90332 35000 90336
rect 34936 90276 34940 90332
rect 34940 90276 34996 90332
rect 34996 90276 35000 90332
rect 34936 90272 35000 90276
rect 35016 90332 35080 90336
rect 35016 90276 35020 90332
rect 35020 90276 35076 90332
rect 35076 90276 35080 90332
rect 35016 90272 35080 90276
rect 35096 90332 35160 90336
rect 35096 90276 35100 90332
rect 35100 90276 35156 90332
rect 35156 90276 35160 90332
rect 35096 90272 35160 90276
rect 35176 90332 35240 90336
rect 35176 90276 35180 90332
rect 35180 90276 35236 90332
rect 35236 90276 35240 90332
rect 35176 90272 35240 90276
rect 65656 90332 65720 90336
rect 65656 90276 65660 90332
rect 65660 90276 65716 90332
rect 65716 90276 65720 90332
rect 65656 90272 65720 90276
rect 65736 90332 65800 90336
rect 65736 90276 65740 90332
rect 65740 90276 65796 90332
rect 65796 90276 65800 90332
rect 65736 90272 65800 90276
rect 65816 90332 65880 90336
rect 65816 90276 65820 90332
rect 65820 90276 65876 90332
rect 65876 90276 65880 90332
rect 65816 90272 65880 90276
rect 65896 90332 65960 90336
rect 65896 90276 65900 90332
rect 65900 90276 65956 90332
rect 65956 90276 65960 90332
rect 65896 90272 65960 90276
rect 96376 90332 96440 90336
rect 96376 90276 96380 90332
rect 96380 90276 96436 90332
rect 96436 90276 96440 90332
rect 96376 90272 96440 90276
rect 96456 90332 96520 90336
rect 96456 90276 96460 90332
rect 96460 90276 96516 90332
rect 96516 90276 96520 90332
rect 96456 90272 96520 90276
rect 96536 90332 96600 90336
rect 96536 90276 96540 90332
rect 96540 90276 96596 90332
rect 96596 90276 96600 90332
rect 96536 90272 96600 90276
rect 96616 90332 96680 90336
rect 96616 90276 96620 90332
rect 96620 90276 96676 90332
rect 96676 90276 96680 90332
rect 96616 90272 96680 90276
rect 127096 90332 127160 90336
rect 127096 90276 127100 90332
rect 127100 90276 127156 90332
rect 127156 90276 127160 90332
rect 127096 90272 127160 90276
rect 127176 90332 127240 90336
rect 127176 90276 127180 90332
rect 127180 90276 127236 90332
rect 127236 90276 127240 90332
rect 127176 90272 127240 90276
rect 127256 90332 127320 90336
rect 127256 90276 127260 90332
rect 127260 90276 127316 90332
rect 127316 90276 127320 90332
rect 127256 90272 127320 90276
rect 127336 90332 127400 90336
rect 127336 90276 127340 90332
rect 127340 90276 127396 90332
rect 127396 90276 127400 90332
rect 127336 90272 127400 90276
rect 157816 90332 157880 90336
rect 157816 90276 157820 90332
rect 157820 90276 157876 90332
rect 157876 90276 157880 90332
rect 157816 90272 157880 90276
rect 157896 90332 157960 90336
rect 157896 90276 157900 90332
rect 157900 90276 157956 90332
rect 157956 90276 157960 90332
rect 157896 90272 157960 90276
rect 157976 90332 158040 90336
rect 157976 90276 157980 90332
rect 157980 90276 158036 90332
rect 158036 90276 158040 90332
rect 157976 90272 158040 90276
rect 158056 90332 158120 90336
rect 158056 90276 158060 90332
rect 158060 90276 158116 90332
rect 158116 90276 158120 90332
rect 158056 90272 158120 90276
rect 19576 89788 19640 89792
rect 19576 89732 19580 89788
rect 19580 89732 19636 89788
rect 19636 89732 19640 89788
rect 19576 89728 19640 89732
rect 19656 89788 19720 89792
rect 19656 89732 19660 89788
rect 19660 89732 19716 89788
rect 19716 89732 19720 89788
rect 19656 89728 19720 89732
rect 19736 89788 19800 89792
rect 19736 89732 19740 89788
rect 19740 89732 19796 89788
rect 19796 89732 19800 89788
rect 19736 89728 19800 89732
rect 19816 89788 19880 89792
rect 19816 89732 19820 89788
rect 19820 89732 19876 89788
rect 19876 89732 19880 89788
rect 19816 89728 19880 89732
rect 50296 89788 50360 89792
rect 50296 89732 50300 89788
rect 50300 89732 50356 89788
rect 50356 89732 50360 89788
rect 50296 89728 50360 89732
rect 50376 89788 50440 89792
rect 50376 89732 50380 89788
rect 50380 89732 50436 89788
rect 50436 89732 50440 89788
rect 50376 89728 50440 89732
rect 50456 89788 50520 89792
rect 50456 89732 50460 89788
rect 50460 89732 50516 89788
rect 50516 89732 50520 89788
rect 50456 89728 50520 89732
rect 50536 89788 50600 89792
rect 50536 89732 50540 89788
rect 50540 89732 50596 89788
rect 50596 89732 50600 89788
rect 50536 89728 50600 89732
rect 81016 89788 81080 89792
rect 81016 89732 81020 89788
rect 81020 89732 81076 89788
rect 81076 89732 81080 89788
rect 81016 89728 81080 89732
rect 81096 89788 81160 89792
rect 81096 89732 81100 89788
rect 81100 89732 81156 89788
rect 81156 89732 81160 89788
rect 81096 89728 81160 89732
rect 81176 89788 81240 89792
rect 81176 89732 81180 89788
rect 81180 89732 81236 89788
rect 81236 89732 81240 89788
rect 81176 89728 81240 89732
rect 81256 89788 81320 89792
rect 81256 89732 81260 89788
rect 81260 89732 81316 89788
rect 81316 89732 81320 89788
rect 81256 89728 81320 89732
rect 111736 89788 111800 89792
rect 111736 89732 111740 89788
rect 111740 89732 111796 89788
rect 111796 89732 111800 89788
rect 111736 89728 111800 89732
rect 111816 89788 111880 89792
rect 111816 89732 111820 89788
rect 111820 89732 111876 89788
rect 111876 89732 111880 89788
rect 111816 89728 111880 89732
rect 111896 89788 111960 89792
rect 111896 89732 111900 89788
rect 111900 89732 111956 89788
rect 111956 89732 111960 89788
rect 111896 89728 111960 89732
rect 111976 89788 112040 89792
rect 111976 89732 111980 89788
rect 111980 89732 112036 89788
rect 112036 89732 112040 89788
rect 111976 89728 112040 89732
rect 142456 89788 142520 89792
rect 142456 89732 142460 89788
rect 142460 89732 142516 89788
rect 142516 89732 142520 89788
rect 142456 89728 142520 89732
rect 142536 89788 142600 89792
rect 142536 89732 142540 89788
rect 142540 89732 142596 89788
rect 142596 89732 142600 89788
rect 142536 89728 142600 89732
rect 142616 89788 142680 89792
rect 142616 89732 142620 89788
rect 142620 89732 142676 89788
rect 142676 89732 142680 89788
rect 142616 89728 142680 89732
rect 142696 89788 142760 89792
rect 142696 89732 142700 89788
rect 142700 89732 142756 89788
rect 142756 89732 142760 89788
rect 142696 89728 142760 89732
rect 173176 89788 173240 89792
rect 173176 89732 173180 89788
rect 173180 89732 173236 89788
rect 173236 89732 173240 89788
rect 173176 89728 173240 89732
rect 173256 89788 173320 89792
rect 173256 89732 173260 89788
rect 173260 89732 173316 89788
rect 173316 89732 173320 89788
rect 173256 89728 173320 89732
rect 173336 89788 173400 89792
rect 173336 89732 173340 89788
rect 173340 89732 173396 89788
rect 173396 89732 173400 89788
rect 173336 89728 173400 89732
rect 173416 89788 173480 89792
rect 173416 89732 173420 89788
rect 173420 89732 173476 89788
rect 173476 89732 173480 89788
rect 173416 89728 173480 89732
rect 4216 89244 4280 89248
rect 4216 89188 4220 89244
rect 4220 89188 4276 89244
rect 4276 89188 4280 89244
rect 4216 89184 4280 89188
rect 4296 89244 4360 89248
rect 4296 89188 4300 89244
rect 4300 89188 4356 89244
rect 4356 89188 4360 89244
rect 4296 89184 4360 89188
rect 4376 89244 4440 89248
rect 4376 89188 4380 89244
rect 4380 89188 4436 89244
rect 4436 89188 4440 89244
rect 4376 89184 4440 89188
rect 4456 89244 4520 89248
rect 4456 89188 4460 89244
rect 4460 89188 4516 89244
rect 4516 89188 4520 89244
rect 4456 89184 4520 89188
rect 34936 89244 35000 89248
rect 34936 89188 34940 89244
rect 34940 89188 34996 89244
rect 34996 89188 35000 89244
rect 34936 89184 35000 89188
rect 35016 89244 35080 89248
rect 35016 89188 35020 89244
rect 35020 89188 35076 89244
rect 35076 89188 35080 89244
rect 35016 89184 35080 89188
rect 35096 89244 35160 89248
rect 35096 89188 35100 89244
rect 35100 89188 35156 89244
rect 35156 89188 35160 89244
rect 35096 89184 35160 89188
rect 35176 89244 35240 89248
rect 35176 89188 35180 89244
rect 35180 89188 35236 89244
rect 35236 89188 35240 89244
rect 35176 89184 35240 89188
rect 65656 89244 65720 89248
rect 65656 89188 65660 89244
rect 65660 89188 65716 89244
rect 65716 89188 65720 89244
rect 65656 89184 65720 89188
rect 65736 89244 65800 89248
rect 65736 89188 65740 89244
rect 65740 89188 65796 89244
rect 65796 89188 65800 89244
rect 65736 89184 65800 89188
rect 65816 89244 65880 89248
rect 65816 89188 65820 89244
rect 65820 89188 65876 89244
rect 65876 89188 65880 89244
rect 65816 89184 65880 89188
rect 65896 89244 65960 89248
rect 65896 89188 65900 89244
rect 65900 89188 65956 89244
rect 65956 89188 65960 89244
rect 65896 89184 65960 89188
rect 96376 89244 96440 89248
rect 96376 89188 96380 89244
rect 96380 89188 96436 89244
rect 96436 89188 96440 89244
rect 96376 89184 96440 89188
rect 96456 89244 96520 89248
rect 96456 89188 96460 89244
rect 96460 89188 96516 89244
rect 96516 89188 96520 89244
rect 96456 89184 96520 89188
rect 96536 89244 96600 89248
rect 96536 89188 96540 89244
rect 96540 89188 96596 89244
rect 96596 89188 96600 89244
rect 96536 89184 96600 89188
rect 96616 89244 96680 89248
rect 96616 89188 96620 89244
rect 96620 89188 96676 89244
rect 96676 89188 96680 89244
rect 96616 89184 96680 89188
rect 127096 89244 127160 89248
rect 127096 89188 127100 89244
rect 127100 89188 127156 89244
rect 127156 89188 127160 89244
rect 127096 89184 127160 89188
rect 127176 89244 127240 89248
rect 127176 89188 127180 89244
rect 127180 89188 127236 89244
rect 127236 89188 127240 89244
rect 127176 89184 127240 89188
rect 127256 89244 127320 89248
rect 127256 89188 127260 89244
rect 127260 89188 127316 89244
rect 127316 89188 127320 89244
rect 127256 89184 127320 89188
rect 127336 89244 127400 89248
rect 127336 89188 127340 89244
rect 127340 89188 127396 89244
rect 127396 89188 127400 89244
rect 127336 89184 127400 89188
rect 157816 89244 157880 89248
rect 157816 89188 157820 89244
rect 157820 89188 157876 89244
rect 157876 89188 157880 89244
rect 157816 89184 157880 89188
rect 157896 89244 157960 89248
rect 157896 89188 157900 89244
rect 157900 89188 157956 89244
rect 157956 89188 157960 89244
rect 157896 89184 157960 89188
rect 157976 89244 158040 89248
rect 157976 89188 157980 89244
rect 157980 89188 158036 89244
rect 158036 89188 158040 89244
rect 157976 89184 158040 89188
rect 158056 89244 158120 89248
rect 158056 89188 158060 89244
rect 158060 89188 158116 89244
rect 158116 89188 158120 89244
rect 158056 89184 158120 89188
rect 19576 88700 19640 88704
rect 19576 88644 19580 88700
rect 19580 88644 19636 88700
rect 19636 88644 19640 88700
rect 19576 88640 19640 88644
rect 19656 88700 19720 88704
rect 19656 88644 19660 88700
rect 19660 88644 19716 88700
rect 19716 88644 19720 88700
rect 19656 88640 19720 88644
rect 19736 88700 19800 88704
rect 19736 88644 19740 88700
rect 19740 88644 19796 88700
rect 19796 88644 19800 88700
rect 19736 88640 19800 88644
rect 19816 88700 19880 88704
rect 19816 88644 19820 88700
rect 19820 88644 19876 88700
rect 19876 88644 19880 88700
rect 19816 88640 19880 88644
rect 50296 88700 50360 88704
rect 50296 88644 50300 88700
rect 50300 88644 50356 88700
rect 50356 88644 50360 88700
rect 50296 88640 50360 88644
rect 50376 88700 50440 88704
rect 50376 88644 50380 88700
rect 50380 88644 50436 88700
rect 50436 88644 50440 88700
rect 50376 88640 50440 88644
rect 50456 88700 50520 88704
rect 50456 88644 50460 88700
rect 50460 88644 50516 88700
rect 50516 88644 50520 88700
rect 50456 88640 50520 88644
rect 50536 88700 50600 88704
rect 50536 88644 50540 88700
rect 50540 88644 50596 88700
rect 50596 88644 50600 88700
rect 50536 88640 50600 88644
rect 81016 88700 81080 88704
rect 81016 88644 81020 88700
rect 81020 88644 81076 88700
rect 81076 88644 81080 88700
rect 81016 88640 81080 88644
rect 81096 88700 81160 88704
rect 81096 88644 81100 88700
rect 81100 88644 81156 88700
rect 81156 88644 81160 88700
rect 81096 88640 81160 88644
rect 81176 88700 81240 88704
rect 81176 88644 81180 88700
rect 81180 88644 81236 88700
rect 81236 88644 81240 88700
rect 81176 88640 81240 88644
rect 81256 88700 81320 88704
rect 81256 88644 81260 88700
rect 81260 88644 81316 88700
rect 81316 88644 81320 88700
rect 81256 88640 81320 88644
rect 111736 88700 111800 88704
rect 111736 88644 111740 88700
rect 111740 88644 111796 88700
rect 111796 88644 111800 88700
rect 111736 88640 111800 88644
rect 111816 88700 111880 88704
rect 111816 88644 111820 88700
rect 111820 88644 111876 88700
rect 111876 88644 111880 88700
rect 111816 88640 111880 88644
rect 111896 88700 111960 88704
rect 111896 88644 111900 88700
rect 111900 88644 111956 88700
rect 111956 88644 111960 88700
rect 111896 88640 111960 88644
rect 111976 88700 112040 88704
rect 111976 88644 111980 88700
rect 111980 88644 112036 88700
rect 112036 88644 112040 88700
rect 111976 88640 112040 88644
rect 142456 88700 142520 88704
rect 142456 88644 142460 88700
rect 142460 88644 142516 88700
rect 142516 88644 142520 88700
rect 142456 88640 142520 88644
rect 142536 88700 142600 88704
rect 142536 88644 142540 88700
rect 142540 88644 142596 88700
rect 142596 88644 142600 88700
rect 142536 88640 142600 88644
rect 142616 88700 142680 88704
rect 142616 88644 142620 88700
rect 142620 88644 142676 88700
rect 142676 88644 142680 88700
rect 142616 88640 142680 88644
rect 142696 88700 142760 88704
rect 142696 88644 142700 88700
rect 142700 88644 142756 88700
rect 142756 88644 142760 88700
rect 142696 88640 142760 88644
rect 173176 88700 173240 88704
rect 173176 88644 173180 88700
rect 173180 88644 173236 88700
rect 173236 88644 173240 88700
rect 173176 88640 173240 88644
rect 173256 88700 173320 88704
rect 173256 88644 173260 88700
rect 173260 88644 173316 88700
rect 173316 88644 173320 88700
rect 173256 88640 173320 88644
rect 173336 88700 173400 88704
rect 173336 88644 173340 88700
rect 173340 88644 173396 88700
rect 173396 88644 173400 88700
rect 173336 88640 173400 88644
rect 173416 88700 173480 88704
rect 173416 88644 173420 88700
rect 173420 88644 173476 88700
rect 173476 88644 173480 88700
rect 173416 88640 173480 88644
rect 4216 88156 4280 88160
rect 4216 88100 4220 88156
rect 4220 88100 4276 88156
rect 4276 88100 4280 88156
rect 4216 88096 4280 88100
rect 4296 88156 4360 88160
rect 4296 88100 4300 88156
rect 4300 88100 4356 88156
rect 4356 88100 4360 88156
rect 4296 88096 4360 88100
rect 4376 88156 4440 88160
rect 4376 88100 4380 88156
rect 4380 88100 4436 88156
rect 4436 88100 4440 88156
rect 4376 88096 4440 88100
rect 4456 88156 4520 88160
rect 4456 88100 4460 88156
rect 4460 88100 4516 88156
rect 4516 88100 4520 88156
rect 4456 88096 4520 88100
rect 34936 88156 35000 88160
rect 34936 88100 34940 88156
rect 34940 88100 34996 88156
rect 34996 88100 35000 88156
rect 34936 88096 35000 88100
rect 35016 88156 35080 88160
rect 35016 88100 35020 88156
rect 35020 88100 35076 88156
rect 35076 88100 35080 88156
rect 35016 88096 35080 88100
rect 35096 88156 35160 88160
rect 35096 88100 35100 88156
rect 35100 88100 35156 88156
rect 35156 88100 35160 88156
rect 35096 88096 35160 88100
rect 35176 88156 35240 88160
rect 35176 88100 35180 88156
rect 35180 88100 35236 88156
rect 35236 88100 35240 88156
rect 35176 88096 35240 88100
rect 65656 88156 65720 88160
rect 65656 88100 65660 88156
rect 65660 88100 65716 88156
rect 65716 88100 65720 88156
rect 65656 88096 65720 88100
rect 65736 88156 65800 88160
rect 65736 88100 65740 88156
rect 65740 88100 65796 88156
rect 65796 88100 65800 88156
rect 65736 88096 65800 88100
rect 65816 88156 65880 88160
rect 65816 88100 65820 88156
rect 65820 88100 65876 88156
rect 65876 88100 65880 88156
rect 65816 88096 65880 88100
rect 65896 88156 65960 88160
rect 65896 88100 65900 88156
rect 65900 88100 65956 88156
rect 65956 88100 65960 88156
rect 65896 88096 65960 88100
rect 96376 88156 96440 88160
rect 96376 88100 96380 88156
rect 96380 88100 96436 88156
rect 96436 88100 96440 88156
rect 96376 88096 96440 88100
rect 96456 88156 96520 88160
rect 96456 88100 96460 88156
rect 96460 88100 96516 88156
rect 96516 88100 96520 88156
rect 96456 88096 96520 88100
rect 96536 88156 96600 88160
rect 96536 88100 96540 88156
rect 96540 88100 96596 88156
rect 96596 88100 96600 88156
rect 96536 88096 96600 88100
rect 96616 88156 96680 88160
rect 96616 88100 96620 88156
rect 96620 88100 96676 88156
rect 96676 88100 96680 88156
rect 96616 88096 96680 88100
rect 127096 88156 127160 88160
rect 127096 88100 127100 88156
rect 127100 88100 127156 88156
rect 127156 88100 127160 88156
rect 127096 88096 127160 88100
rect 127176 88156 127240 88160
rect 127176 88100 127180 88156
rect 127180 88100 127236 88156
rect 127236 88100 127240 88156
rect 127176 88096 127240 88100
rect 127256 88156 127320 88160
rect 127256 88100 127260 88156
rect 127260 88100 127316 88156
rect 127316 88100 127320 88156
rect 127256 88096 127320 88100
rect 127336 88156 127400 88160
rect 127336 88100 127340 88156
rect 127340 88100 127396 88156
rect 127396 88100 127400 88156
rect 127336 88096 127400 88100
rect 157816 88156 157880 88160
rect 157816 88100 157820 88156
rect 157820 88100 157876 88156
rect 157876 88100 157880 88156
rect 157816 88096 157880 88100
rect 157896 88156 157960 88160
rect 157896 88100 157900 88156
rect 157900 88100 157956 88156
rect 157956 88100 157960 88156
rect 157896 88096 157960 88100
rect 157976 88156 158040 88160
rect 157976 88100 157980 88156
rect 157980 88100 158036 88156
rect 158036 88100 158040 88156
rect 157976 88096 158040 88100
rect 158056 88156 158120 88160
rect 158056 88100 158060 88156
rect 158060 88100 158116 88156
rect 158116 88100 158120 88156
rect 158056 88096 158120 88100
rect 19576 87612 19640 87616
rect 19576 87556 19580 87612
rect 19580 87556 19636 87612
rect 19636 87556 19640 87612
rect 19576 87552 19640 87556
rect 19656 87612 19720 87616
rect 19656 87556 19660 87612
rect 19660 87556 19716 87612
rect 19716 87556 19720 87612
rect 19656 87552 19720 87556
rect 19736 87612 19800 87616
rect 19736 87556 19740 87612
rect 19740 87556 19796 87612
rect 19796 87556 19800 87612
rect 19736 87552 19800 87556
rect 19816 87612 19880 87616
rect 19816 87556 19820 87612
rect 19820 87556 19876 87612
rect 19876 87556 19880 87612
rect 19816 87552 19880 87556
rect 50296 87612 50360 87616
rect 50296 87556 50300 87612
rect 50300 87556 50356 87612
rect 50356 87556 50360 87612
rect 50296 87552 50360 87556
rect 50376 87612 50440 87616
rect 50376 87556 50380 87612
rect 50380 87556 50436 87612
rect 50436 87556 50440 87612
rect 50376 87552 50440 87556
rect 50456 87612 50520 87616
rect 50456 87556 50460 87612
rect 50460 87556 50516 87612
rect 50516 87556 50520 87612
rect 50456 87552 50520 87556
rect 50536 87612 50600 87616
rect 50536 87556 50540 87612
rect 50540 87556 50596 87612
rect 50596 87556 50600 87612
rect 50536 87552 50600 87556
rect 81016 87612 81080 87616
rect 81016 87556 81020 87612
rect 81020 87556 81076 87612
rect 81076 87556 81080 87612
rect 81016 87552 81080 87556
rect 81096 87612 81160 87616
rect 81096 87556 81100 87612
rect 81100 87556 81156 87612
rect 81156 87556 81160 87612
rect 81096 87552 81160 87556
rect 81176 87612 81240 87616
rect 81176 87556 81180 87612
rect 81180 87556 81236 87612
rect 81236 87556 81240 87612
rect 81176 87552 81240 87556
rect 81256 87612 81320 87616
rect 81256 87556 81260 87612
rect 81260 87556 81316 87612
rect 81316 87556 81320 87612
rect 81256 87552 81320 87556
rect 111736 87612 111800 87616
rect 111736 87556 111740 87612
rect 111740 87556 111796 87612
rect 111796 87556 111800 87612
rect 111736 87552 111800 87556
rect 111816 87612 111880 87616
rect 111816 87556 111820 87612
rect 111820 87556 111876 87612
rect 111876 87556 111880 87612
rect 111816 87552 111880 87556
rect 111896 87612 111960 87616
rect 111896 87556 111900 87612
rect 111900 87556 111956 87612
rect 111956 87556 111960 87612
rect 111896 87552 111960 87556
rect 111976 87612 112040 87616
rect 111976 87556 111980 87612
rect 111980 87556 112036 87612
rect 112036 87556 112040 87612
rect 111976 87552 112040 87556
rect 142456 87612 142520 87616
rect 142456 87556 142460 87612
rect 142460 87556 142516 87612
rect 142516 87556 142520 87612
rect 142456 87552 142520 87556
rect 142536 87612 142600 87616
rect 142536 87556 142540 87612
rect 142540 87556 142596 87612
rect 142596 87556 142600 87612
rect 142536 87552 142600 87556
rect 142616 87612 142680 87616
rect 142616 87556 142620 87612
rect 142620 87556 142676 87612
rect 142676 87556 142680 87612
rect 142616 87552 142680 87556
rect 142696 87612 142760 87616
rect 142696 87556 142700 87612
rect 142700 87556 142756 87612
rect 142756 87556 142760 87612
rect 142696 87552 142760 87556
rect 173176 87612 173240 87616
rect 173176 87556 173180 87612
rect 173180 87556 173236 87612
rect 173236 87556 173240 87612
rect 173176 87552 173240 87556
rect 173256 87612 173320 87616
rect 173256 87556 173260 87612
rect 173260 87556 173316 87612
rect 173316 87556 173320 87612
rect 173256 87552 173320 87556
rect 173336 87612 173400 87616
rect 173336 87556 173340 87612
rect 173340 87556 173396 87612
rect 173396 87556 173400 87612
rect 173336 87552 173400 87556
rect 173416 87612 173480 87616
rect 173416 87556 173420 87612
rect 173420 87556 173476 87612
rect 173476 87556 173480 87612
rect 173416 87552 173480 87556
rect 4216 87068 4280 87072
rect 4216 87012 4220 87068
rect 4220 87012 4276 87068
rect 4276 87012 4280 87068
rect 4216 87008 4280 87012
rect 4296 87068 4360 87072
rect 4296 87012 4300 87068
rect 4300 87012 4356 87068
rect 4356 87012 4360 87068
rect 4296 87008 4360 87012
rect 4376 87068 4440 87072
rect 4376 87012 4380 87068
rect 4380 87012 4436 87068
rect 4436 87012 4440 87068
rect 4376 87008 4440 87012
rect 4456 87068 4520 87072
rect 4456 87012 4460 87068
rect 4460 87012 4516 87068
rect 4516 87012 4520 87068
rect 4456 87008 4520 87012
rect 34936 87068 35000 87072
rect 34936 87012 34940 87068
rect 34940 87012 34996 87068
rect 34996 87012 35000 87068
rect 34936 87008 35000 87012
rect 35016 87068 35080 87072
rect 35016 87012 35020 87068
rect 35020 87012 35076 87068
rect 35076 87012 35080 87068
rect 35016 87008 35080 87012
rect 35096 87068 35160 87072
rect 35096 87012 35100 87068
rect 35100 87012 35156 87068
rect 35156 87012 35160 87068
rect 35096 87008 35160 87012
rect 35176 87068 35240 87072
rect 35176 87012 35180 87068
rect 35180 87012 35236 87068
rect 35236 87012 35240 87068
rect 35176 87008 35240 87012
rect 65656 87068 65720 87072
rect 65656 87012 65660 87068
rect 65660 87012 65716 87068
rect 65716 87012 65720 87068
rect 65656 87008 65720 87012
rect 65736 87068 65800 87072
rect 65736 87012 65740 87068
rect 65740 87012 65796 87068
rect 65796 87012 65800 87068
rect 65736 87008 65800 87012
rect 65816 87068 65880 87072
rect 65816 87012 65820 87068
rect 65820 87012 65876 87068
rect 65876 87012 65880 87068
rect 65816 87008 65880 87012
rect 65896 87068 65960 87072
rect 65896 87012 65900 87068
rect 65900 87012 65956 87068
rect 65956 87012 65960 87068
rect 65896 87008 65960 87012
rect 96376 87068 96440 87072
rect 96376 87012 96380 87068
rect 96380 87012 96436 87068
rect 96436 87012 96440 87068
rect 96376 87008 96440 87012
rect 96456 87068 96520 87072
rect 96456 87012 96460 87068
rect 96460 87012 96516 87068
rect 96516 87012 96520 87068
rect 96456 87008 96520 87012
rect 96536 87068 96600 87072
rect 96536 87012 96540 87068
rect 96540 87012 96596 87068
rect 96596 87012 96600 87068
rect 96536 87008 96600 87012
rect 96616 87068 96680 87072
rect 96616 87012 96620 87068
rect 96620 87012 96676 87068
rect 96676 87012 96680 87068
rect 96616 87008 96680 87012
rect 127096 87068 127160 87072
rect 127096 87012 127100 87068
rect 127100 87012 127156 87068
rect 127156 87012 127160 87068
rect 127096 87008 127160 87012
rect 127176 87068 127240 87072
rect 127176 87012 127180 87068
rect 127180 87012 127236 87068
rect 127236 87012 127240 87068
rect 127176 87008 127240 87012
rect 127256 87068 127320 87072
rect 127256 87012 127260 87068
rect 127260 87012 127316 87068
rect 127316 87012 127320 87068
rect 127256 87008 127320 87012
rect 127336 87068 127400 87072
rect 127336 87012 127340 87068
rect 127340 87012 127396 87068
rect 127396 87012 127400 87068
rect 127336 87008 127400 87012
rect 157816 87068 157880 87072
rect 157816 87012 157820 87068
rect 157820 87012 157876 87068
rect 157876 87012 157880 87068
rect 157816 87008 157880 87012
rect 157896 87068 157960 87072
rect 157896 87012 157900 87068
rect 157900 87012 157956 87068
rect 157956 87012 157960 87068
rect 157896 87008 157960 87012
rect 157976 87068 158040 87072
rect 157976 87012 157980 87068
rect 157980 87012 158036 87068
rect 158036 87012 158040 87068
rect 157976 87008 158040 87012
rect 158056 87068 158120 87072
rect 158056 87012 158060 87068
rect 158060 87012 158116 87068
rect 158116 87012 158120 87068
rect 158056 87008 158120 87012
rect 19576 86524 19640 86528
rect 19576 86468 19580 86524
rect 19580 86468 19636 86524
rect 19636 86468 19640 86524
rect 19576 86464 19640 86468
rect 19656 86524 19720 86528
rect 19656 86468 19660 86524
rect 19660 86468 19716 86524
rect 19716 86468 19720 86524
rect 19656 86464 19720 86468
rect 19736 86524 19800 86528
rect 19736 86468 19740 86524
rect 19740 86468 19796 86524
rect 19796 86468 19800 86524
rect 19736 86464 19800 86468
rect 19816 86524 19880 86528
rect 19816 86468 19820 86524
rect 19820 86468 19876 86524
rect 19876 86468 19880 86524
rect 19816 86464 19880 86468
rect 50296 86524 50360 86528
rect 50296 86468 50300 86524
rect 50300 86468 50356 86524
rect 50356 86468 50360 86524
rect 50296 86464 50360 86468
rect 50376 86524 50440 86528
rect 50376 86468 50380 86524
rect 50380 86468 50436 86524
rect 50436 86468 50440 86524
rect 50376 86464 50440 86468
rect 50456 86524 50520 86528
rect 50456 86468 50460 86524
rect 50460 86468 50516 86524
rect 50516 86468 50520 86524
rect 50456 86464 50520 86468
rect 50536 86524 50600 86528
rect 50536 86468 50540 86524
rect 50540 86468 50596 86524
rect 50596 86468 50600 86524
rect 50536 86464 50600 86468
rect 81016 86524 81080 86528
rect 81016 86468 81020 86524
rect 81020 86468 81076 86524
rect 81076 86468 81080 86524
rect 81016 86464 81080 86468
rect 81096 86524 81160 86528
rect 81096 86468 81100 86524
rect 81100 86468 81156 86524
rect 81156 86468 81160 86524
rect 81096 86464 81160 86468
rect 81176 86524 81240 86528
rect 81176 86468 81180 86524
rect 81180 86468 81236 86524
rect 81236 86468 81240 86524
rect 81176 86464 81240 86468
rect 81256 86524 81320 86528
rect 81256 86468 81260 86524
rect 81260 86468 81316 86524
rect 81316 86468 81320 86524
rect 81256 86464 81320 86468
rect 111736 86524 111800 86528
rect 111736 86468 111740 86524
rect 111740 86468 111796 86524
rect 111796 86468 111800 86524
rect 111736 86464 111800 86468
rect 111816 86524 111880 86528
rect 111816 86468 111820 86524
rect 111820 86468 111876 86524
rect 111876 86468 111880 86524
rect 111816 86464 111880 86468
rect 111896 86524 111960 86528
rect 111896 86468 111900 86524
rect 111900 86468 111956 86524
rect 111956 86468 111960 86524
rect 111896 86464 111960 86468
rect 111976 86524 112040 86528
rect 111976 86468 111980 86524
rect 111980 86468 112036 86524
rect 112036 86468 112040 86524
rect 111976 86464 112040 86468
rect 142456 86524 142520 86528
rect 142456 86468 142460 86524
rect 142460 86468 142516 86524
rect 142516 86468 142520 86524
rect 142456 86464 142520 86468
rect 142536 86524 142600 86528
rect 142536 86468 142540 86524
rect 142540 86468 142596 86524
rect 142596 86468 142600 86524
rect 142536 86464 142600 86468
rect 142616 86524 142680 86528
rect 142616 86468 142620 86524
rect 142620 86468 142676 86524
rect 142676 86468 142680 86524
rect 142616 86464 142680 86468
rect 142696 86524 142760 86528
rect 142696 86468 142700 86524
rect 142700 86468 142756 86524
rect 142756 86468 142760 86524
rect 142696 86464 142760 86468
rect 173176 86524 173240 86528
rect 173176 86468 173180 86524
rect 173180 86468 173236 86524
rect 173236 86468 173240 86524
rect 173176 86464 173240 86468
rect 173256 86524 173320 86528
rect 173256 86468 173260 86524
rect 173260 86468 173316 86524
rect 173316 86468 173320 86524
rect 173256 86464 173320 86468
rect 173336 86524 173400 86528
rect 173336 86468 173340 86524
rect 173340 86468 173396 86524
rect 173396 86468 173400 86524
rect 173336 86464 173400 86468
rect 173416 86524 173480 86528
rect 173416 86468 173420 86524
rect 173420 86468 173476 86524
rect 173476 86468 173480 86524
rect 173416 86464 173480 86468
rect 4216 85980 4280 85984
rect 4216 85924 4220 85980
rect 4220 85924 4276 85980
rect 4276 85924 4280 85980
rect 4216 85920 4280 85924
rect 4296 85980 4360 85984
rect 4296 85924 4300 85980
rect 4300 85924 4356 85980
rect 4356 85924 4360 85980
rect 4296 85920 4360 85924
rect 4376 85980 4440 85984
rect 4376 85924 4380 85980
rect 4380 85924 4436 85980
rect 4436 85924 4440 85980
rect 4376 85920 4440 85924
rect 4456 85980 4520 85984
rect 4456 85924 4460 85980
rect 4460 85924 4516 85980
rect 4516 85924 4520 85980
rect 4456 85920 4520 85924
rect 34936 85980 35000 85984
rect 34936 85924 34940 85980
rect 34940 85924 34996 85980
rect 34996 85924 35000 85980
rect 34936 85920 35000 85924
rect 35016 85980 35080 85984
rect 35016 85924 35020 85980
rect 35020 85924 35076 85980
rect 35076 85924 35080 85980
rect 35016 85920 35080 85924
rect 35096 85980 35160 85984
rect 35096 85924 35100 85980
rect 35100 85924 35156 85980
rect 35156 85924 35160 85980
rect 35096 85920 35160 85924
rect 35176 85980 35240 85984
rect 35176 85924 35180 85980
rect 35180 85924 35236 85980
rect 35236 85924 35240 85980
rect 35176 85920 35240 85924
rect 65656 85980 65720 85984
rect 65656 85924 65660 85980
rect 65660 85924 65716 85980
rect 65716 85924 65720 85980
rect 65656 85920 65720 85924
rect 65736 85980 65800 85984
rect 65736 85924 65740 85980
rect 65740 85924 65796 85980
rect 65796 85924 65800 85980
rect 65736 85920 65800 85924
rect 65816 85980 65880 85984
rect 65816 85924 65820 85980
rect 65820 85924 65876 85980
rect 65876 85924 65880 85980
rect 65816 85920 65880 85924
rect 65896 85980 65960 85984
rect 65896 85924 65900 85980
rect 65900 85924 65956 85980
rect 65956 85924 65960 85980
rect 65896 85920 65960 85924
rect 96376 85980 96440 85984
rect 96376 85924 96380 85980
rect 96380 85924 96436 85980
rect 96436 85924 96440 85980
rect 96376 85920 96440 85924
rect 96456 85980 96520 85984
rect 96456 85924 96460 85980
rect 96460 85924 96516 85980
rect 96516 85924 96520 85980
rect 96456 85920 96520 85924
rect 96536 85980 96600 85984
rect 96536 85924 96540 85980
rect 96540 85924 96596 85980
rect 96596 85924 96600 85980
rect 96536 85920 96600 85924
rect 96616 85980 96680 85984
rect 96616 85924 96620 85980
rect 96620 85924 96676 85980
rect 96676 85924 96680 85980
rect 96616 85920 96680 85924
rect 127096 85980 127160 85984
rect 127096 85924 127100 85980
rect 127100 85924 127156 85980
rect 127156 85924 127160 85980
rect 127096 85920 127160 85924
rect 127176 85980 127240 85984
rect 127176 85924 127180 85980
rect 127180 85924 127236 85980
rect 127236 85924 127240 85980
rect 127176 85920 127240 85924
rect 127256 85980 127320 85984
rect 127256 85924 127260 85980
rect 127260 85924 127316 85980
rect 127316 85924 127320 85980
rect 127256 85920 127320 85924
rect 127336 85980 127400 85984
rect 127336 85924 127340 85980
rect 127340 85924 127396 85980
rect 127396 85924 127400 85980
rect 127336 85920 127400 85924
rect 157816 85980 157880 85984
rect 157816 85924 157820 85980
rect 157820 85924 157876 85980
rect 157876 85924 157880 85980
rect 157816 85920 157880 85924
rect 157896 85980 157960 85984
rect 157896 85924 157900 85980
rect 157900 85924 157956 85980
rect 157956 85924 157960 85980
rect 157896 85920 157960 85924
rect 157976 85980 158040 85984
rect 157976 85924 157980 85980
rect 157980 85924 158036 85980
rect 158036 85924 158040 85980
rect 157976 85920 158040 85924
rect 158056 85980 158120 85984
rect 158056 85924 158060 85980
rect 158060 85924 158116 85980
rect 158116 85924 158120 85980
rect 158056 85920 158120 85924
rect 19576 85436 19640 85440
rect 19576 85380 19580 85436
rect 19580 85380 19636 85436
rect 19636 85380 19640 85436
rect 19576 85376 19640 85380
rect 19656 85436 19720 85440
rect 19656 85380 19660 85436
rect 19660 85380 19716 85436
rect 19716 85380 19720 85436
rect 19656 85376 19720 85380
rect 19736 85436 19800 85440
rect 19736 85380 19740 85436
rect 19740 85380 19796 85436
rect 19796 85380 19800 85436
rect 19736 85376 19800 85380
rect 19816 85436 19880 85440
rect 19816 85380 19820 85436
rect 19820 85380 19876 85436
rect 19876 85380 19880 85436
rect 19816 85376 19880 85380
rect 50296 85436 50360 85440
rect 50296 85380 50300 85436
rect 50300 85380 50356 85436
rect 50356 85380 50360 85436
rect 50296 85376 50360 85380
rect 50376 85436 50440 85440
rect 50376 85380 50380 85436
rect 50380 85380 50436 85436
rect 50436 85380 50440 85436
rect 50376 85376 50440 85380
rect 50456 85436 50520 85440
rect 50456 85380 50460 85436
rect 50460 85380 50516 85436
rect 50516 85380 50520 85436
rect 50456 85376 50520 85380
rect 50536 85436 50600 85440
rect 50536 85380 50540 85436
rect 50540 85380 50596 85436
rect 50596 85380 50600 85436
rect 50536 85376 50600 85380
rect 81016 85436 81080 85440
rect 81016 85380 81020 85436
rect 81020 85380 81076 85436
rect 81076 85380 81080 85436
rect 81016 85376 81080 85380
rect 81096 85436 81160 85440
rect 81096 85380 81100 85436
rect 81100 85380 81156 85436
rect 81156 85380 81160 85436
rect 81096 85376 81160 85380
rect 81176 85436 81240 85440
rect 81176 85380 81180 85436
rect 81180 85380 81236 85436
rect 81236 85380 81240 85436
rect 81176 85376 81240 85380
rect 81256 85436 81320 85440
rect 81256 85380 81260 85436
rect 81260 85380 81316 85436
rect 81316 85380 81320 85436
rect 81256 85376 81320 85380
rect 111736 85436 111800 85440
rect 111736 85380 111740 85436
rect 111740 85380 111796 85436
rect 111796 85380 111800 85436
rect 111736 85376 111800 85380
rect 111816 85436 111880 85440
rect 111816 85380 111820 85436
rect 111820 85380 111876 85436
rect 111876 85380 111880 85436
rect 111816 85376 111880 85380
rect 111896 85436 111960 85440
rect 111896 85380 111900 85436
rect 111900 85380 111956 85436
rect 111956 85380 111960 85436
rect 111896 85376 111960 85380
rect 111976 85436 112040 85440
rect 111976 85380 111980 85436
rect 111980 85380 112036 85436
rect 112036 85380 112040 85436
rect 111976 85376 112040 85380
rect 142456 85436 142520 85440
rect 142456 85380 142460 85436
rect 142460 85380 142516 85436
rect 142516 85380 142520 85436
rect 142456 85376 142520 85380
rect 142536 85436 142600 85440
rect 142536 85380 142540 85436
rect 142540 85380 142596 85436
rect 142596 85380 142600 85436
rect 142536 85376 142600 85380
rect 142616 85436 142680 85440
rect 142616 85380 142620 85436
rect 142620 85380 142676 85436
rect 142676 85380 142680 85436
rect 142616 85376 142680 85380
rect 142696 85436 142760 85440
rect 142696 85380 142700 85436
rect 142700 85380 142756 85436
rect 142756 85380 142760 85436
rect 142696 85376 142760 85380
rect 173176 85436 173240 85440
rect 173176 85380 173180 85436
rect 173180 85380 173236 85436
rect 173236 85380 173240 85436
rect 173176 85376 173240 85380
rect 173256 85436 173320 85440
rect 173256 85380 173260 85436
rect 173260 85380 173316 85436
rect 173316 85380 173320 85436
rect 173256 85376 173320 85380
rect 173336 85436 173400 85440
rect 173336 85380 173340 85436
rect 173340 85380 173396 85436
rect 173396 85380 173400 85436
rect 173336 85376 173400 85380
rect 173416 85436 173480 85440
rect 173416 85380 173420 85436
rect 173420 85380 173476 85436
rect 173476 85380 173480 85436
rect 173416 85376 173480 85380
rect 4216 84892 4280 84896
rect 4216 84836 4220 84892
rect 4220 84836 4276 84892
rect 4276 84836 4280 84892
rect 4216 84832 4280 84836
rect 4296 84892 4360 84896
rect 4296 84836 4300 84892
rect 4300 84836 4356 84892
rect 4356 84836 4360 84892
rect 4296 84832 4360 84836
rect 4376 84892 4440 84896
rect 4376 84836 4380 84892
rect 4380 84836 4436 84892
rect 4436 84836 4440 84892
rect 4376 84832 4440 84836
rect 4456 84892 4520 84896
rect 4456 84836 4460 84892
rect 4460 84836 4516 84892
rect 4516 84836 4520 84892
rect 4456 84832 4520 84836
rect 34936 84892 35000 84896
rect 34936 84836 34940 84892
rect 34940 84836 34996 84892
rect 34996 84836 35000 84892
rect 34936 84832 35000 84836
rect 35016 84892 35080 84896
rect 35016 84836 35020 84892
rect 35020 84836 35076 84892
rect 35076 84836 35080 84892
rect 35016 84832 35080 84836
rect 35096 84892 35160 84896
rect 35096 84836 35100 84892
rect 35100 84836 35156 84892
rect 35156 84836 35160 84892
rect 35096 84832 35160 84836
rect 35176 84892 35240 84896
rect 35176 84836 35180 84892
rect 35180 84836 35236 84892
rect 35236 84836 35240 84892
rect 35176 84832 35240 84836
rect 65656 84892 65720 84896
rect 65656 84836 65660 84892
rect 65660 84836 65716 84892
rect 65716 84836 65720 84892
rect 65656 84832 65720 84836
rect 65736 84892 65800 84896
rect 65736 84836 65740 84892
rect 65740 84836 65796 84892
rect 65796 84836 65800 84892
rect 65736 84832 65800 84836
rect 65816 84892 65880 84896
rect 65816 84836 65820 84892
rect 65820 84836 65876 84892
rect 65876 84836 65880 84892
rect 65816 84832 65880 84836
rect 65896 84892 65960 84896
rect 65896 84836 65900 84892
rect 65900 84836 65956 84892
rect 65956 84836 65960 84892
rect 65896 84832 65960 84836
rect 96376 84892 96440 84896
rect 96376 84836 96380 84892
rect 96380 84836 96436 84892
rect 96436 84836 96440 84892
rect 96376 84832 96440 84836
rect 96456 84892 96520 84896
rect 96456 84836 96460 84892
rect 96460 84836 96516 84892
rect 96516 84836 96520 84892
rect 96456 84832 96520 84836
rect 96536 84892 96600 84896
rect 96536 84836 96540 84892
rect 96540 84836 96596 84892
rect 96596 84836 96600 84892
rect 96536 84832 96600 84836
rect 96616 84892 96680 84896
rect 96616 84836 96620 84892
rect 96620 84836 96676 84892
rect 96676 84836 96680 84892
rect 96616 84832 96680 84836
rect 127096 84892 127160 84896
rect 127096 84836 127100 84892
rect 127100 84836 127156 84892
rect 127156 84836 127160 84892
rect 127096 84832 127160 84836
rect 127176 84892 127240 84896
rect 127176 84836 127180 84892
rect 127180 84836 127236 84892
rect 127236 84836 127240 84892
rect 127176 84832 127240 84836
rect 127256 84892 127320 84896
rect 127256 84836 127260 84892
rect 127260 84836 127316 84892
rect 127316 84836 127320 84892
rect 127256 84832 127320 84836
rect 127336 84892 127400 84896
rect 127336 84836 127340 84892
rect 127340 84836 127396 84892
rect 127396 84836 127400 84892
rect 127336 84832 127400 84836
rect 157816 84892 157880 84896
rect 157816 84836 157820 84892
rect 157820 84836 157876 84892
rect 157876 84836 157880 84892
rect 157816 84832 157880 84836
rect 157896 84892 157960 84896
rect 157896 84836 157900 84892
rect 157900 84836 157956 84892
rect 157956 84836 157960 84892
rect 157896 84832 157960 84836
rect 157976 84892 158040 84896
rect 157976 84836 157980 84892
rect 157980 84836 158036 84892
rect 158036 84836 158040 84892
rect 157976 84832 158040 84836
rect 158056 84892 158120 84896
rect 158056 84836 158060 84892
rect 158060 84836 158116 84892
rect 158116 84836 158120 84892
rect 158056 84832 158120 84836
rect 19576 84348 19640 84352
rect 19576 84292 19580 84348
rect 19580 84292 19636 84348
rect 19636 84292 19640 84348
rect 19576 84288 19640 84292
rect 19656 84348 19720 84352
rect 19656 84292 19660 84348
rect 19660 84292 19716 84348
rect 19716 84292 19720 84348
rect 19656 84288 19720 84292
rect 19736 84348 19800 84352
rect 19736 84292 19740 84348
rect 19740 84292 19796 84348
rect 19796 84292 19800 84348
rect 19736 84288 19800 84292
rect 19816 84348 19880 84352
rect 19816 84292 19820 84348
rect 19820 84292 19876 84348
rect 19876 84292 19880 84348
rect 19816 84288 19880 84292
rect 50296 84348 50360 84352
rect 50296 84292 50300 84348
rect 50300 84292 50356 84348
rect 50356 84292 50360 84348
rect 50296 84288 50360 84292
rect 50376 84348 50440 84352
rect 50376 84292 50380 84348
rect 50380 84292 50436 84348
rect 50436 84292 50440 84348
rect 50376 84288 50440 84292
rect 50456 84348 50520 84352
rect 50456 84292 50460 84348
rect 50460 84292 50516 84348
rect 50516 84292 50520 84348
rect 50456 84288 50520 84292
rect 50536 84348 50600 84352
rect 50536 84292 50540 84348
rect 50540 84292 50596 84348
rect 50596 84292 50600 84348
rect 50536 84288 50600 84292
rect 81016 84348 81080 84352
rect 81016 84292 81020 84348
rect 81020 84292 81076 84348
rect 81076 84292 81080 84348
rect 81016 84288 81080 84292
rect 81096 84348 81160 84352
rect 81096 84292 81100 84348
rect 81100 84292 81156 84348
rect 81156 84292 81160 84348
rect 81096 84288 81160 84292
rect 81176 84348 81240 84352
rect 81176 84292 81180 84348
rect 81180 84292 81236 84348
rect 81236 84292 81240 84348
rect 81176 84288 81240 84292
rect 81256 84348 81320 84352
rect 81256 84292 81260 84348
rect 81260 84292 81316 84348
rect 81316 84292 81320 84348
rect 81256 84288 81320 84292
rect 111736 84348 111800 84352
rect 111736 84292 111740 84348
rect 111740 84292 111796 84348
rect 111796 84292 111800 84348
rect 111736 84288 111800 84292
rect 111816 84348 111880 84352
rect 111816 84292 111820 84348
rect 111820 84292 111876 84348
rect 111876 84292 111880 84348
rect 111816 84288 111880 84292
rect 111896 84348 111960 84352
rect 111896 84292 111900 84348
rect 111900 84292 111956 84348
rect 111956 84292 111960 84348
rect 111896 84288 111960 84292
rect 111976 84348 112040 84352
rect 111976 84292 111980 84348
rect 111980 84292 112036 84348
rect 112036 84292 112040 84348
rect 111976 84288 112040 84292
rect 142456 84348 142520 84352
rect 142456 84292 142460 84348
rect 142460 84292 142516 84348
rect 142516 84292 142520 84348
rect 142456 84288 142520 84292
rect 142536 84348 142600 84352
rect 142536 84292 142540 84348
rect 142540 84292 142596 84348
rect 142596 84292 142600 84348
rect 142536 84288 142600 84292
rect 142616 84348 142680 84352
rect 142616 84292 142620 84348
rect 142620 84292 142676 84348
rect 142676 84292 142680 84348
rect 142616 84288 142680 84292
rect 142696 84348 142760 84352
rect 142696 84292 142700 84348
rect 142700 84292 142756 84348
rect 142756 84292 142760 84348
rect 142696 84288 142760 84292
rect 173176 84348 173240 84352
rect 173176 84292 173180 84348
rect 173180 84292 173236 84348
rect 173236 84292 173240 84348
rect 173176 84288 173240 84292
rect 173256 84348 173320 84352
rect 173256 84292 173260 84348
rect 173260 84292 173316 84348
rect 173316 84292 173320 84348
rect 173256 84288 173320 84292
rect 173336 84348 173400 84352
rect 173336 84292 173340 84348
rect 173340 84292 173396 84348
rect 173396 84292 173400 84348
rect 173336 84288 173400 84292
rect 173416 84348 173480 84352
rect 173416 84292 173420 84348
rect 173420 84292 173476 84348
rect 173476 84292 173480 84348
rect 173416 84288 173480 84292
rect 4216 83804 4280 83808
rect 4216 83748 4220 83804
rect 4220 83748 4276 83804
rect 4276 83748 4280 83804
rect 4216 83744 4280 83748
rect 4296 83804 4360 83808
rect 4296 83748 4300 83804
rect 4300 83748 4356 83804
rect 4356 83748 4360 83804
rect 4296 83744 4360 83748
rect 4376 83804 4440 83808
rect 4376 83748 4380 83804
rect 4380 83748 4436 83804
rect 4436 83748 4440 83804
rect 4376 83744 4440 83748
rect 4456 83804 4520 83808
rect 4456 83748 4460 83804
rect 4460 83748 4516 83804
rect 4516 83748 4520 83804
rect 4456 83744 4520 83748
rect 34936 83804 35000 83808
rect 34936 83748 34940 83804
rect 34940 83748 34996 83804
rect 34996 83748 35000 83804
rect 34936 83744 35000 83748
rect 35016 83804 35080 83808
rect 35016 83748 35020 83804
rect 35020 83748 35076 83804
rect 35076 83748 35080 83804
rect 35016 83744 35080 83748
rect 35096 83804 35160 83808
rect 35096 83748 35100 83804
rect 35100 83748 35156 83804
rect 35156 83748 35160 83804
rect 35096 83744 35160 83748
rect 35176 83804 35240 83808
rect 35176 83748 35180 83804
rect 35180 83748 35236 83804
rect 35236 83748 35240 83804
rect 35176 83744 35240 83748
rect 65656 83804 65720 83808
rect 65656 83748 65660 83804
rect 65660 83748 65716 83804
rect 65716 83748 65720 83804
rect 65656 83744 65720 83748
rect 65736 83804 65800 83808
rect 65736 83748 65740 83804
rect 65740 83748 65796 83804
rect 65796 83748 65800 83804
rect 65736 83744 65800 83748
rect 65816 83804 65880 83808
rect 65816 83748 65820 83804
rect 65820 83748 65876 83804
rect 65876 83748 65880 83804
rect 65816 83744 65880 83748
rect 65896 83804 65960 83808
rect 65896 83748 65900 83804
rect 65900 83748 65956 83804
rect 65956 83748 65960 83804
rect 65896 83744 65960 83748
rect 96376 83804 96440 83808
rect 96376 83748 96380 83804
rect 96380 83748 96436 83804
rect 96436 83748 96440 83804
rect 96376 83744 96440 83748
rect 96456 83804 96520 83808
rect 96456 83748 96460 83804
rect 96460 83748 96516 83804
rect 96516 83748 96520 83804
rect 96456 83744 96520 83748
rect 96536 83804 96600 83808
rect 96536 83748 96540 83804
rect 96540 83748 96596 83804
rect 96596 83748 96600 83804
rect 96536 83744 96600 83748
rect 96616 83804 96680 83808
rect 96616 83748 96620 83804
rect 96620 83748 96676 83804
rect 96676 83748 96680 83804
rect 96616 83744 96680 83748
rect 127096 83804 127160 83808
rect 127096 83748 127100 83804
rect 127100 83748 127156 83804
rect 127156 83748 127160 83804
rect 127096 83744 127160 83748
rect 127176 83804 127240 83808
rect 127176 83748 127180 83804
rect 127180 83748 127236 83804
rect 127236 83748 127240 83804
rect 127176 83744 127240 83748
rect 127256 83804 127320 83808
rect 127256 83748 127260 83804
rect 127260 83748 127316 83804
rect 127316 83748 127320 83804
rect 127256 83744 127320 83748
rect 127336 83804 127400 83808
rect 127336 83748 127340 83804
rect 127340 83748 127396 83804
rect 127396 83748 127400 83804
rect 127336 83744 127400 83748
rect 157816 83804 157880 83808
rect 157816 83748 157820 83804
rect 157820 83748 157876 83804
rect 157876 83748 157880 83804
rect 157816 83744 157880 83748
rect 157896 83804 157960 83808
rect 157896 83748 157900 83804
rect 157900 83748 157956 83804
rect 157956 83748 157960 83804
rect 157896 83744 157960 83748
rect 157976 83804 158040 83808
rect 157976 83748 157980 83804
rect 157980 83748 158036 83804
rect 158036 83748 158040 83804
rect 157976 83744 158040 83748
rect 158056 83804 158120 83808
rect 158056 83748 158060 83804
rect 158060 83748 158116 83804
rect 158116 83748 158120 83804
rect 158056 83744 158120 83748
rect 19576 83260 19640 83264
rect 19576 83204 19580 83260
rect 19580 83204 19636 83260
rect 19636 83204 19640 83260
rect 19576 83200 19640 83204
rect 19656 83260 19720 83264
rect 19656 83204 19660 83260
rect 19660 83204 19716 83260
rect 19716 83204 19720 83260
rect 19656 83200 19720 83204
rect 19736 83260 19800 83264
rect 19736 83204 19740 83260
rect 19740 83204 19796 83260
rect 19796 83204 19800 83260
rect 19736 83200 19800 83204
rect 19816 83260 19880 83264
rect 19816 83204 19820 83260
rect 19820 83204 19876 83260
rect 19876 83204 19880 83260
rect 19816 83200 19880 83204
rect 50296 83260 50360 83264
rect 50296 83204 50300 83260
rect 50300 83204 50356 83260
rect 50356 83204 50360 83260
rect 50296 83200 50360 83204
rect 50376 83260 50440 83264
rect 50376 83204 50380 83260
rect 50380 83204 50436 83260
rect 50436 83204 50440 83260
rect 50376 83200 50440 83204
rect 50456 83260 50520 83264
rect 50456 83204 50460 83260
rect 50460 83204 50516 83260
rect 50516 83204 50520 83260
rect 50456 83200 50520 83204
rect 50536 83260 50600 83264
rect 50536 83204 50540 83260
rect 50540 83204 50596 83260
rect 50596 83204 50600 83260
rect 50536 83200 50600 83204
rect 81016 83260 81080 83264
rect 81016 83204 81020 83260
rect 81020 83204 81076 83260
rect 81076 83204 81080 83260
rect 81016 83200 81080 83204
rect 81096 83260 81160 83264
rect 81096 83204 81100 83260
rect 81100 83204 81156 83260
rect 81156 83204 81160 83260
rect 81096 83200 81160 83204
rect 81176 83260 81240 83264
rect 81176 83204 81180 83260
rect 81180 83204 81236 83260
rect 81236 83204 81240 83260
rect 81176 83200 81240 83204
rect 81256 83260 81320 83264
rect 81256 83204 81260 83260
rect 81260 83204 81316 83260
rect 81316 83204 81320 83260
rect 81256 83200 81320 83204
rect 111736 83260 111800 83264
rect 111736 83204 111740 83260
rect 111740 83204 111796 83260
rect 111796 83204 111800 83260
rect 111736 83200 111800 83204
rect 111816 83260 111880 83264
rect 111816 83204 111820 83260
rect 111820 83204 111876 83260
rect 111876 83204 111880 83260
rect 111816 83200 111880 83204
rect 111896 83260 111960 83264
rect 111896 83204 111900 83260
rect 111900 83204 111956 83260
rect 111956 83204 111960 83260
rect 111896 83200 111960 83204
rect 111976 83260 112040 83264
rect 111976 83204 111980 83260
rect 111980 83204 112036 83260
rect 112036 83204 112040 83260
rect 111976 83200 112040 83204
rect 142456 83260 142520 83264
rect 142456 83204 142460 83260
rect 142460 83204 142516 83260
rect 142516 83204 142520 83260
rect 142456 83200 142520 83204
rect 142536 83260 142600 83264
rect 142536 83204 142540 83260
rect 142540 83204 142596 83260
rect 142596 83204 142600 83260
rect 142536 83200 142600 83204
rect 142616 83260 142680 83264
rect 142616 83204 142620 83260
rect 142620 83204 142676 83260
rect 142676 83204 142680 83260
rect 142616 83200 142680 83204
rect 142696 83260 142760 83264
rect 142696 83204 142700 83260
rect 142700 83204 142756 83260
rect 142756 83204 142760 83260
rect 142696 83200 142760 83204
rect 173176 83260 173240 83264
rect 173176 83204 173180 83260
rect 173180 83204 173236 83260
rect 173236 83204 173240 83260
rect 173176 83200 173240 83204
rect 173256 83260 173320 83264
rect 173256 83204 173260 83260
rect 173260 83204 173316 83260
rect 173316 83204 173320 83260
rect 173256 83200 173320 83204
rect 173336 83260 173400 83264
rect 173336 83204 173340 83260
rect 173340 83204 173396 83260
rect 173396 83204 173400 83260
rect 173336 83200 173400 83204
rect 173416 83260 173480 83264
rect 173416 83204 173420 83260
rect 173420 83204 173476 83260
rect 173476 83204 173480 83260
rect 173416 83200 173480 83204
rect 4216 82716 4280 82720
rect 4216 82660 4220 82716
rect 4220 82660 4276 82716
rect 4276 82660 4280 82716
rect 4216 82656 4280 82660
rect 4296 82716 4360 82720
rect 4296 82660 4300 82716
rect 4300 82660 4356 82716
rect 4356 82660 4360 82716
rect 4296 82656 4360 82660
rect 4376 82716 4440 82720
rect 4376 82660 4380 82716
rect 4380 82660 4436 82716
rect 4436 82660 4440 82716
rect 4376 82656 4440 82660
rect 4456 82716 4520 82720
rect 4456 82660 4460 82716
rect 4460 82660 4516 82716
rect 4516 82660 4520 82716
rect 4456 82656 4520 82660
rect 34936 82716 35000 82720
rect 34936 82660 34940 82716
rect 34940 82660 34996 82716
rect 34996 82660 35000 82716
rect 34936 82656 35000 82660
rect 35016 82716 35080 82720
rect 35016 82660 35020 82716
rect 35020 82660 35076 82716
rect 35076 82660 35080 82716
rect 35016 82656 35080 82660
rect 35096 82716 35160 82720
rect 35096 82660 35100 82716
rect 35100 82660 35156 82716
rect 35156 82660 35160 82716
rect 35096 82656 35160 82660
rect 35176 82716 35240 82720
rect 35176 82660 35180 82716
rect 35180 82660 35236 82716
rect 35236 82660 35240 82716
rect 35176 82656 35240 82660
rect 65656 82716 65720 82720
rect 65656 82660 65660 82716
rect 65660 82660 65716 82716
rect 65716 82660 65720 82716
rect 65656 82656 65720 82660
rect 65736 82716 65800 82720
rect 65736 82660 65740 82716
rect 65740 82660 65796 82716
rect 65796 82660 65800 82716
rect 65736 82656 65800 82660
rect 65816 82716 65880 82720
rect 65816 82660 65820 82716
rect 65820 82660 65876 82716
rect 65876 82660 65880 82716
rect 65816 82656 65880 82660
rect 65896 82716 65960 82720
rect 65896 82660 65900 82716
rect 65900 82660 65956 82716
rect 65956 82660 65960 82716
rect 65896 82656 65960 82660
rect 96376 82716 96440 82720
rect 96376 82660 96380 82716
rect 96380 82660 96436 82716
rect 96436 82660 96440 82716
rect 96376 82656 96440 82660
rect 96456 82716 96520 82720
rect 96456 82660 96460 82716
rect 96460 82660 96516 82716
rect 96516 82660 96520 82716
rect 96456 82656 96520 82660
rect 96536 82716 96600 82720
rect 96536 82660 96540 82716
rect 96540 82660 96596 82716
rect 96596 82660 96600 82716
rect 96536 82656 96600 82660
rect 96616 82716 96680 82720
rect 96616 82660 96620 82716
rect 96620 82660 96676 82716
rect 96676 82660 96680 82716
rect 96616 82656 96680 82660
rect 127096 82716 127160 82720
rect 127096 82660 127100 82716
rect 127100 82660 127156 82716
rect 127156 82660 127160 82716
rect 127096 82656 127160 82660
rect 127176 82716 127240 82720
rect 127176 82660 127180 82716
rect 127180 82660 127236 82716
rect 127236 82660 127240 82716
rect 127176 82656 127240 82660
rect 127256 82716 127320 82720
rect 127256 82660 127260 82716
rect 127260 82660 127316 82716
rect 127316 82660 127320 82716
rect 127256 82656 127320 82660
rect 127336 82716 127400 82720
rect 127336 82660 127340 82716
rect 127340 82660 127396 82716
rect 127396 82660 127400 82716
rect 127336 82656 127400 82660
rect 157816 82716 157880 82720
rect 157816 82660 157820 82716
rect 157820 82660 157876 82716
rect 157876 82660 157880 82716
rect 157816 82656 157880 82660
rect 157896 82716 157960 82720
rect 157896 82660 157900 82716
rect 157900 82660 157956 82716
rect 157956 82660 157960 82716
rect 157896 82656 157960 82660
rect 157976 82716 158040 82720
rect 157976 82660 157980 82716
rect 157980 82660 158036 82716
rect 158036 82660 158040 82716
rect 157976 82656 158040 82660
rect 158056 82716 158120 82720
rect 158056 82660 158060 82716
rect 158060 82660 158116 82716
rect 158116 82660 158120 82716
rect 158056 82656 158120 82660
rect 19576 82172 19640 82176
rect 19576 82116 19580 82172
rect 19580 82116 19636 82172
rect 19636 82116 19640 82172
rect 19576 82112 19640 82116
rect 19656 82172 19720 82176
rect 19656 82116 19660 82172
rect 19660 82116 19716 82172
rect 19716 82116 19720 82172
rect 19656 82112 19720 82116
rect 19736 82172 19800 82176
rect 19736 82116 19740 82172
rect 19740 82116 19796 82172
rect 19796 82116 19800 82172
rect 19736 82112 19800 82116
rect 19816 82172 19880 82176
rect 19816 82116 19820 82172
rect 19820 82116 19876 82172
rect 19876 82116 19880 82172
rect 19816 82112 19880 82116
rect 50296 82172 50360 82176
rect 50296 82116 50300 82172
rect 50300 82116 50356 82172
rect 50356 82116 50360 82172
rect 50296 82112 50360 82116
rect 50376 82172 50440 82176
rect 50376 82116 50380 82172
rect 50380 82116 50436 82172
rect 50436 82116 50440 82172
rect 50376 82112 50440 82116
rect 50456 82172 50520 82176
rect 50456 82116 50460 82172
rect 50460 82116 50516 82172
rect 50516 82116 50520 82172
rect 50456 82112 50520 82116
rect 50536 82172 50600 82176
rect 50536 82116 50540 82172
rect 50540 82116 50596 82172
rect 50596 82116 50600 82172
rect 50536 82112 50600 82116
rect 81016 82172 81080 82176
rect 81016 82116 81020 82172
rect 81020 82116 81076 82172
rect 81076 82116 81080 82172
rect 81016 82112 81080 82116
rect 81096 82172 81160 82176
rect 81096 82116 81100 82172
rect 81100 82116 81156 82172
rect 81156 82116 81160 82172
rect 81096 82112 81160 82116
rect 81176 82172 81240 82176
rect 81176 82116 81180 82172
rect 81180 82116 81236 82172
rect 81236 82116 81240 82172
rect 81176 82112 81240 82116
rect 81256 82172 81320 82176
rect 81256 82116 81260 82172
rect 81260 82116 81316 82172
rect 81316 82116 81320 82172
rect 81256 82112 81320 82116
rect 111736 82172 111800 82176
rect 111736 82116 111740 82172
rect 111740 82116 111796 82172
rect 111796 82116 111800 82172
rect 111736 82112 111800 82116
rect 111816 82172 111880 82176
rect 111816 82116 111820 82172
rect 111820 82116 111876 82172
rect 111876 82116 111880 82172
rect 111816 82112 111880 82116
rect 111896 82172 111960 82176
rect 111896 82116 111900 82172
rect 111900 82116 111956 82172
rect 111956 82116 111960 82172
rect 111896 82112 111960 82116
rect 111976 82172 112040 82176
rect 111976 82116 111980 82172
rect 111980 82116 112036 82172
rect 112036 82116 112040 82172
rect 111976 82112 112040 82116
rect 142456 82172 142520 82176
rect 142456 82116 142460 82172
rect 142460 82116 142516 82172
rect 142516 82116 142520 82172
rect 142456 82112 142520 82116
rect 142536 82172 142600 82176
rect 142536 82116 142540 82172
rect 142540 82116 142596 82172
rect 142596 82116 142600 82172
rect 142536 82112 142600 82116
rect 142616 82172 142680 82176
rect 142616 82116 142620 82172
rect 142620 82116 142676 82172
rect 142676 82116 142680 82172
rect 142616 82112 142680 82116
rect 142696 82172 142760 82176
rect 142696 82116 142700 82172
rect 142700 82116 142756 82172
rect 142756 82116 142760 82172
rect 142696 82112 142760 82116
rect 173176 82172 173240 82176
rect 173176 82116 173180 82172
rect 173180 82116 173236 82172
rect 173236 82116 173240 82172
rect 173176 82112 173240 82116
rect 173256 82172 173320 82176
rect 173256 82116 173260 82172
rect 173260 82116 173316 82172
rect 173316 82116 173320 82172
rect 173256 82112 173320 82116
rect 173336 82172 173400 82176
rect 173336 82116 173340 82172
rect 173340 82116 173396 82172
rect 173396 82116 173400 82172
rect 173336 82112 173400 82116
rect 173416 82172 173480 82176
rect 173416 82116 173420 82172
rect 173420 82116 173476 82172
rect 173476 82116 173480 82172
rect 173416 82112 173480 82116
rect 4216 81628 4280 81632
rect 4216 81572 4220 81628
rect 4220 81572 4276 81628
rect 4276 81572 4280 81628
rect 4216 81568 4280 81572
rect 4296 81628 4360 81632
rect 4296 81572 4300 81628
rect 4300 81572 4356 81628
rect 4356 81572 4360 81628
rect 4296 81568 4360 81572
rect 4376 81628 4440 81632
rect 4376 81572 4380 81628
rect 4380 81572 4436 81628
rect 4436 81572 4440 81628
rect 4376 81568 4440 81572
rect 4456 81628 4520 81632
rect 4456 81572 4460 81628
rect 4460 81572 4516 81628
rect 4516 81572 4520 81628
rect 4456 81568 4520 81572
rect 34936 81628 35000 81632
rect 34936 81572 34940 81628
rect 34940 81572 34996 81628
rect 34996 81572 35000 81628
rect 34936 81568 35000 81572
rect 35016 81628 35080 81632
rect 35016 81572 35020 81628
rect 35020 81572 35076 81628
rect 35076 81572 35080 81628
rect 35016 81568 35080 81572
rect 35096 81628 35160 81632
rect 35096 81572 35100 81628
rect 35100 81572 35156 81628
rect 35156 81572 35160 81628
rect 35096 81568 35160 81572
rect 35176 81628 35240 81632
rect 35176 81572 35180 81628
rect 35180 81572 35236 81628
rect 35236 81572 35240 81628
rect 35176 81568 35240 81572
rect 65656 81628 65720 81632
rect 65656 81572 65660 81628
rect 65660 81572 65716 81628
rect 65716 81572 65720 81628
rect 65656 81568 65720 81572
rect 65736 81628 65800 81632
rect 65736 81572 65740 81628
rect 65740 81572 65796 81628
rect 65796 81572 65800 81628
rect 65736 81568 65800 81572
rect 65816 81628 65880 81632
rect 65816 81572 65820 81628
rect 65820 81572 65876 81628
rect 65876 81572 65880 81628
rect 65816 81568 65880 81572
rect 65896 81628 65960 81632
rect 65896 81572 65900 81628
rect 65900 81572 65956 81628
rect 65956 81572 65960 81628
rect 65896 81568 65960 81572
rect 96376 81628 96440 81632
rect 96376 81572 96380 81628
rect 96380 81572 96436 81628
rect 96436 81572 96440 81628
rect 96376 81568 96440 81572
rect 96456 81628 96520 81632
rect 96456 81572 96460 81628
rect 96460 81572 96516 81628
rect 96516 81572 96520 81628
rect 96456 81568 96520 81572
rect 96536 81628 96600 81632
rect 96536 81572 96540 81628
rect 96540 81572 96596 81628
rect 96596 81572 96600 81628
rect 96536 81568 96600 81572
rect 96616 81628 96680 81632
rect 96616 81572 96620 81628
rect 96620 81572 96676 81628
rect 96676 81572 96680 81628
rect 96616 81568 96680 81572
rect 127096 81628 127160 81632
rect 127096 81572 127100 81628
rect 127100 81572 127156 81628
rect 127156 81572 127160 81628
rect 127096 81568 127160 81572
rect 127176 81628 127240 81632
rect 127176 81572 127180 81628
rect 127180 81572 127236 81628
rect 127236 81572 127240 81628
rect 127176 81568 127240 81572
rect 127256 81628 127320 81632
rect 127256 81572 127260 81628
rect 127260 81572 127316 81628
rect 127316 81572 127320 81628
rect 127256 81568 127320 81572
rect 127336 81628 127400 81632
rect 127336 81572 127340 81628
rect 127340 81572 127396 81628
rect 127396 81572 127400 81628
rect 127336 81568 127400 81572
rect 157816 81628 157880 81632
rect 157816 81572 157820 81628
rect 157820 81572 157876 81628
rect 157876 81572 157880 81628
rect 157816 81568 157880 81572
rect 157896 81628 157960 81632
rect 157896 81572 157900 81628
rect 157900 81572 157956 81628
rect 157956 81572 157960 81628
rect 157896 81568 157960 81572
rect 157976 81628 158040 81632
rect 157976 81572 157980 81628
rect 157980 81572 158036 81628
rect 158036 81572 158040 81628
rect 157976 81568 158040 81572
rect 158056 81628 158120 81632
rect 158056 81572 158060 81628
rect 158060 81572 158116 81628
rect 158116 81572 158120 81628
rect 158056 81568 158120 81572
rect 19576 81084 19640 81088
rect 19576 81028 19580 81084
rect 19580 81028 19636 81084
rect 19636 81028 19640 81084
rect 19576 81024 19640 81028
rect 19656 81084 19720 81088
rect 19656 81028 19660 81084
rect 19660 81028 19716 81084
rect 19716 81028 19720 81084
rect 19656 81024 19720 81028
rect 19736 81084 19800 81088
rect 19736 81028 19740 81084
rect 19740 81028 19796 81084
rect 19796 81028 19800 81084
rect 19736 81024 19800 81028
rect 19816 81084 19880 81088
rect 19816 81028 19820 81084
rect 19820 81028 19876 81084
rect 19876 81028 19880 81084
rect 19816 81024 19880 81028
rect 50296 81084 50360 81088
rect 50296 81028 50300 81084
rect 50300 81028 50356 81084
rect 50356 81028 50360 81084
rect 50296 81024 50360 81028
rect 50376 81084 50440 81088
rect 50376 81028 50380 81084
rect 50380 81028 50436 81084
rect 50436 81028 50440 81084
rect 50376 81024 50440 81028
rect 50456 81084 50520 81088
rect 50456 81028 50460 81084
rect 50460 81028 50516 81084
rect 50516 81028 50520 81084
rect 50456 81024 50520 81028
rect 50536 81084 50600 81088
rect 50536 81028 50540 81084
rect 50540 81028 50596 81084
rect 50596 81028 50600 81084
rect 50536 81024 50600 81028
rect 81016 81084 81080 81088
rect 81016 81028 81020 81084
rect 81020 81028 81076 81084
rect 81076 81028 81080 81084
rect 81016 81024 81080 81028
rect 81096 81084 81160 81088
rect 81096 81028 81100 81084
rect 81100 81028 81156 81084
rect 81156 81028 81160 81084
rect 81096 81024 81160 81028
rect 81176 81084 81240 81088
rect 81176 81028 81180 81084
rect 81180 81028 81236 81084
rect 81236 81028 81240 81084
rect 81176 81024 81240 81028
rect 81256 81084 81320 81088
rect 81256 81028 81260 81084
rect 81260 81028 81316 81084
rect 81316 81028 81320 81084
rect 81256 81024 81320 81028
rect 111736 81084 111800 81088
rect 111736 81028 111740 81084
rect 111740 81028 111796 81084
rect 111796 81028 111800 81084
rect 111736 81024 111800 81028
rect 111816 81084 111880 81088
rect 111816 81028 111820 81084
rect 111820 81028 111876 81084
rect 111876 81028 111880 81084
rect 111816 81024 111880 81028
rect 111896 81084 111960 81088
rect 111896 81028 111900 81084
rect 111900 81028 111956 81084
rect 111956 81028 111960 81084
rect 111896 81024 111960 81028
rect 111976 81084 112040 81088
rect 111976 81028 111980 81084
rect 111980 81028 112036 81084
rect 112036 81028 112040 81084
rect 111976 81024 112040 81028
rect 142456 81084 142520 81088
rect 142456 81028 142460 81084
rect 142460 81028 142516 81084
rect 142516 81028 142520 81084
rect 142456 81024 142520 81028
rect 142536 81084 142600 81088
rect 142536 81028 142540 81084
rect 142540 81028 142596 81084
rect 142596 81028 142600 81084
rect 142536 81024 142600 81028
rect 142616 81084 142680 81088
rect 142616 81028 142620 81084
rect 142620 81028 142676 81084
rect 142676 81028 142680 81084
rect 142616 81024 142680 81028
rect 142696 81084 142760 81088
rect 142696 81028 142700 81084
rect 142700 81028 142756 81084
rect 142756 81028 142760 81084
rect 142696 81024 142760 81028
rect 173176 81084 173240 81088
rect 173176 81028 173180 81084
rect 173180 81028 173236 81084
rect 173236 81028 173240 81084
rect 173176 81024 173240 81028
rect 173256 81084 173320 81088
rect 173256 81028 173260 81084
rect 173260 81028 173316 81084
rect 173316 81028 173320 81084
rect 173256 81024 173320 81028
rect 173336 81084 173400 81088
rect 173336 81028 173340 81084
rect 173340 81028 173396 81084
rect 173396 81028 173400 81084
rect 173336 81024 173400 81028
rect 173416 81084 173480 81088
rect 173416 81028 173420 81084
rect 173420 81028 173476 81084
rect 173476 81028 173480 81084
rect 173416 81024 173480 81028
rect 4216 80540 4280 80544
rect 4216 80484 4220 80540
rect 4220 80484 4276 80540
rect 4276 80484 4280 80540
rect 4216 80480 4280 80484
rect 4296 80540 4360 80544
rect 4296 80484 4300 80540
rect 4300 80484 4356 80540
rect 4356 80484 4360 80540
rect 4296 80480 4360 80484
rect 4376 80540 4440 80544
rect 4376 80484 4380 80540
rect 4380 80484 4436 80540
rect 4436 80484 4440 80540
rect 4376 80480 4440 80484
rect 4456 80540 4520 80544
rect 4456 80484 4460 80540
rect 4460 80484 4516 80540
rect 4516 80484 4520 80540
rect 4456 80480 4520 80484
rect 34936 80540 35000 80544
rect 34936 80484 34940 80540
rect 34940 80484 34996 80540
rect 34996 80484 35000 80540
rect 34936 80480 35000 80484
rect 35016 80540 35080 80544
rect 35016 80484 35020 80540
rect 35020 80484 35076 80540
rect 35076 80484 35080 80540
rect 35016 80480 35080 80484
rect 35096 80540 35160 80544
rect 35096 80484 35100 80540
rect 35100 80484 35156 80540
rect 35156 80484 35160 80540
rect 35096 80480 35160 80484
rect 35176 80540 35240 80544
rect 35176 80484 35180 80540
rect 35180 80484 35236 80540
rect 35236 80484 35240 80540
rect 35176 80480 35240 80484
rect 65656 80540 65720 80544
rect 65656 80484 65660 80540
rect 65660 80484 65716 80540
rect 65716 80484 65720 80540
rect 65656 80480 65720 80484
rect 65736 80540 65800 80544
rect 65736 80484 65740 80540
rect 65740 80484 65796 80540
rect 65796 80484 65800 80540
rect 65736 80480 65800 80484
rect 65816 80540 65880 80544
rect 65816 80484 65820 80540
rect 65820 80484 65876 80540
rect 65876 80484 65880 80540
rect 65816 80480 65880 80484
rect 65896 80540 65960 80544
rect 65896 80484 65900 80540
rect 65900 80484 65956 80540
rect 65956 80484 65960 80540
rect 65896 80480 65960 80484
rect 96376 80540 96440 80544
rect 96376 80484 96380 80540
rect 96380 80484 96436 80540
rect 96436 80484 96440 80540
rect 96376 80480 96440 80484
rect 96456 80540 96520 80544
rect 96456 80484 96460 80540
rect 96460 80484 96516 80540
rect 96516 80484 96520 80540
rect 96456 80480 96520 80484
rect 96536 80540 96600 80544
rect 96536 80484 96540 80540
rect 96540 80484 96596 80540
rect 96596 80484 96600 80540
rect 96536 80480 96600 80484
rect 96616 80540 96680 80544
rect 96616 80484 96620 80540
rect 96620 80484 96676 80540
rect 96676 80484 96680 80540
rect 96616 80480 96680 80484
rect 127096 80540 127160 80544
rect 127096 80484 127100 80540
rect 127100 80484 127156 80540
rect 127156 80484 127160 80540
rect 127096 80480 127160 80484
rect 127176 80540 127240 80544
rect 127176 80484 127180 80540
rect 127180 80484 127236 80540
rect 127236 80484 127240 80540
rect 127176 80480 127240 80484
rect 127256 80540 127320 80544
rect 127256 80484 127260 80540
rect 127260 80484 127316 80540
rect 127316 80484 127320 80540
rect 127256 80480 127320 80484
rect 127336 80540 127400 80544
rect 127336 80484 127340 80540
rect 127340 80484 127396 80540
rect 127396 80484 127400 80540
rect 127336 80480 127400 80484
rect 157816 80540 157880 80544
rect 157816 80484 157820 80540
rect 157820 80484 157876 80540
rect 157876 80484 157880 80540
rect 157816 80480 157880 80484
rect 157896 80540 157960 80544
rect 157896 80484 157900 80540
rect 157900 80484 157956 80540
rect 157956 80484 157960 80540
rect 157896 80480 157960 80484
rect 157976 80540 158040 80544
rect 157976 80484 157980 80540
rect 157980 80484 158036 80540
rect 158036 80484 158040 80540
rect 157976 80480 158040 80484
rect 158056 80540 158120 80544
rect 158056 80484 158060 80540
rect 158060 80484 158116 80540
rect 158116 80484 158120 80540
rect 158056 80480 158120 80484
rect 19576 79996 19640 80000
rect 19576 79940 19580 79996
rect 19580 79940 19636 79996
rect 19636 79940 19640 79996
rect 19576 79936 19640 79940
rect 19656 79996 19720 80000
rect 19656 79940 19660 79996
rect 19660 79940 19716 79996
rect 19716 79940 19720 79996
rect 19656 79936 19720 79940
rect 19736 79996 19800 80000
rect 19736 79940 19740 79996
rect 19740 79940 19796 79996
rect 19796 79940 19800 79996
rect 19736 79936 19800 79940
rect 19816 79996 19880 80000
rect 19816 79940 19820 79996
rect 19820 79940 19876 79996
rect 19876 79940 19880 79996
rect 19816 79936 19880 79940
rect 50296 79996 50360 80000
rect 50296 79940 50300 79996
rect 50300 79940 50356 79996
rect 50356 79940 50360 79996
rect 50296 79936 50360 79940
rect 50376 79996 50440 80000
rect 50376 79940 50380 79996
rect 50380 79940 50436 79996
rect 50436 79940 50440 79996
rect 50376 79936 50440 79940
rect 50456 79996 50520 80000
rect 50456 79940 50460 79996
rect 50460 79940 50516 79996
rect 50516 79940 50520 79996
rect 50456 79936 50520 79940
rect 50536 79996 50600 80000
rect 50536 79940 50540 79996
rect 50540 79940 50596 79996
rect 50596 79940 50600 79996
rect 50536 79936 50600 79940
rect 81016 79996 81080 80000
rect 81016 79940 81020 79996
rect 81020 79940 81076 79996
rect 81076 79940 81080 79996
rect 81016 79936 81080 79940
rect 81096 79996 81160 80000
rect 81096 79940 81100 79996
rect 81100 79940 81156 79996
rect 81156 79940 81160 79996
rect 81096 79936 81160 79940
rect 81176 79996 81240 80000
rect 81176 79940 81180 79996
rect 81180 79940 81236 79996
rect 81236 79940 81240 79996
rect 81176 79936 81240 79940
rect 81256 79996 81320 80000
rect 81256 79940 81260 79996
rect 81260 79940 81316 79996
rect 81316 79940 81320 79996
rect 81256 79936 81320 79940
rect 111736 79996 111800 80000
rect 111736 79940 111740 79996
rect 111740 79940 111796 79996
rect 111796 79940 111800 79996
rect 111736 79936 111800 79940
rect 111816 79996 111880 80000
rect 111816 79940 111820 79996
rect 111820 79940 111876 79996
rect 111876 79940 111880 79996
rect 111816 79936 111880 79940
rect 111896 79996 111960 80000
rect 111896 79940 111900 79996
rect 111900 79940 111956 79996
rect 111956 79940 111960 79996
rect 111896 79936 111960 79940
rect 111976 79996 112040 80000
rect 111976 79940 111980 79996
rect 111980 79940 112036 79996
rect 112036 79940 112040 79996
rect 111976 79936 112040 79940
rect 142456 79996 142520 80000
rect 142456 79940 142460 79996
rect 142460 79940 142516 79996
rect 142516 79940 142520 79996
rect 142456 79936 142520 79940
rect 142536 79996 142600 80000
rect 142536 79940 142540 79996
rect 142540 79940 142596 79996
rect 142596 79940 142600 79996
rect 142536 79936 142600 79940
rect 142616 79996 142680 80000
rect 142616 79940 142620 79996
rect 142620 79940 142676 79996
rect 142676 79940 142680 79996
rect 142616 79936 142680 79940
rect 142696 79996 142760 80000
rect 142696 79940 142700 79996
rect 142700 79940 142756 79996
rect 142756 79940 142760 79996
rect 142696 79936 142760 79940
rect 173176 79996 173240 80000
rect 173176 79940 173180 79996
rect 173180 79940 173236 79996
rect 173236 79940 173240 79996
rect 173176 79936 173240 79940
rect 173256 79996 173320 80000
rect 173256 79940 173260 79996
rect 173260 79940 173316 79996
rect 173316 79940 173320 79996
rect 173256 79936 173320 79940
rect 173336 79996 173400 80000
rect 173336 79940 173340 79996
rect 173340 79940 173396 79996
rect 173396 79940 173400 79996
rect 173336 79936 173400 79940
rect 173416 79996 173480 80000
rect 173416 79940 173420 79996
rect 173420 79940 173476 79996
rect 173476 79940 173480 79996
rect 173416 79936 173480 79940
rect 4216 79452 4280 79456
rect 4216 79396 4220 79452
rect 4220 79396 4276 79452
rect 4276 79396 4280 79452
rect 4216 79392 4280 79396
rect 4296 79452 4360 79456
rect 4296 79396 4300 79452
rect 4300 79396 4356 79452
rect 4356 79396 4360 79452
rect 4296 79392 4360 79396
rect 4376 79452 4440 79456
rect 4376 79396 4380 79452
rect 4380 79396 4436 79452
rect 4436 79396 4440 79452
rect 4376 79392 4440 79396
rect 4456 79452 4520 79456
rect 4456 79396 4460 79452
rect 4460 79396 4516 79452
rect 4516 79396 4520 79452
rect 4456 79392 4520 79396
rect 34936 79452 35000 79456
rect 34936 79396 34940 79452
rect 34940 79396 34996 79452
rect 34996 79396 35000 79452
rect 34936 79392 35000 79396
rect 35016 79452 35080 79456
rect 35016 79396 35020 79452
rect 35020 79396 35076 79452
rect 35076 79396 35080 79452
rect 35016 79392 35080 79396
rect 35096 79452 35160 79456
rect 35096 79396 35100 79452
rect 35100 79396 35156 79452
rect 35156 79396 35160 79452
rect 35096 79392 35160 79396
rect 35176 79452 35240 79456
rect 35176 79396 35180 79452
rect 35180 79396 35236 79452
rect 35236 79396 35240 79452
rect 35176 79392 35240 79396
rect 65656 79452 65720 79456
rect 65656 79396 65660 79452
rect 65660 79396 65716 79452
rect 65716 79396 65720 79452
rect 65656 79392 65720 79396
rect 65736 79452 65800 79456
rect 65736 79396 65740 79452
rect 65740 79396 65796 79452
rect 65796 79396 65800 79452
rect 65736 79392 65800 79396
rect 65816 79452 65880 79456
rect 65816 79396 65820 79452
rect 65820 79396 65876 79452
rect 65876 79396 65880 79452
rect 65816 79392 65880 79396
rect 65896 79452 65960 79456
rect 65896 79396 65900 79452
rect 65900 79396 65956 79452
rect 65956 79396 65960 79452
rect 65896 79392 65960 79396
rect 96376 79452 96440 79456
rect 96376 79396 96380 79452
rect 96380 79396 96436 79452
rect 96436 79396 96440 79452
rect 96376 79392 96440 79396
rect 96456 79452 96520 79456
rect 96456 79396 96460 79452
rect 96460 79396 96516 79452
rect 96516 79396 96520 79452
rect 96456 79392 96520 79396
rect 96536 79452 96600 79456
rect 96536 79396 96540 79452
rect 96540 79396 96596 79452
rect 96596 79396 96600 79452
rect 96536 79392 96600 79396
rect 96616 79452 96680 79456
rect 96616 79396 96620 79452
rect 96620 79396 96676 79452
rect 96676 79396 96680 79452
rect 96616 79392 96680 79396
rect 127096 79452 127160 79456
rect 127096 79396 127100 79452
rect 127100 79396 127156 79452
rect 127156 79396 127160 79452
rect 127096 79392 127160 79396
rect 127176 79452 127240 79456
rect 127176 79396 127180 79452
rect 127180 79396 127236 79452
rect 127236 79396 127240 79452
rect 127176 79392 127240 79396
rect 127256 79452 127320 79456
rect 127256 79396 127260 79452
rect 127260 79396 127316 79452
rect 127316 79396 127320 79452
rect 127256 79392 127320 79396
rect 127336 79452 127400 79456
rect 127336 79396 127340 79452
rect 127340 79396 127396 79452
rect 127396 79396 127400 79452
rect 127336 79392 127400 79396
rect 157816 79452 157880 79456
rect 157816 79396 157820 79452
rect 157820 79396 157876 79452
rect 157876 79396 157880 79452
rect 157816 79392 157880 79396
rect 157896 79452 157960 79456
rect 157896 79396 157900 79452
rect 157900 79396 157956 79452
rect 157956 79396 157960 79452
rect 157896 79392 157960 79396
rect 157976 79452 158040 79456
rect 157976 79396 157980 79452
rect 157980 79396 158036 79452
rect 158036 79396 158040 79452
rect 157976 79392 158040 79396
rect 158056 79452 158120 79456
rect 158056 79396 158060 79452
rect 158060 79396 158116 79452
rect 158116 79396 158120 79452
rect 158056 79392 158120 79396
rect 19576 78908 19640 78912
rect 19576 78852 19580 78908
rect 19580 78852 19636 78908
rect 19636 78852 19640 78908
rect 19576 78848 19640 78852
rect 19656 78908 19720 78912
rect 19656 78852 19660 78908
rect 19660 78852 19716 78908
rect 19716 78852 19720 78908
rect 19656 78848 19720 78852
rect 19736 78908 19800 78912
rect 19736 78852 19740 78908
rect 19740 78852 19796 78908
rect 19796 78852 19800 78908
rect 19736 78848 19800 78852
rect 19816 78908 19880 78912
rect 19816 78852 19820 78908
rect 19820 78852 19876 78908
rect 19876 78852 19880 78908
rect 19816 78848 19880 78852
rect 50296 78908 50360 78912
rect 50296 78852 50300 78908
rect 50300 78852 50356 78908
rect 50356 78852 50360 78908
rect 50296 78848 50360 78852
rect 50376 78908 50440 78912
rect 50376 78852 50380 78908
rect 50380 78852 50436 78908
rect 50436 78852 50440 78908
rect 50376 78848 50440 78852
rect 50456 78908 50520 78912
rect 50456 78852 50460 78908
rect 50460 78852 50516 78908
rect 50516 78852 50520 78908
rect 50456 78848 50520 78852
rect 50536 78908 50600 78912
rect 50536 78852 50540 78908
rect 50540 78852 50596 78908
rect 50596 78852 50600 78908
rect 50536 78848 50600 78852
rect 81016 78908 81080 78912
rect 81016 78852 81020 78908
rect 81020 78852 81076 78908
rect 81076 78852 81080 78908
rect 81016 78848 81080 78852
rect 81096 78908 81160 78912
rect 81096 78852 81100 78908
rect 81100 78852 81156 78908
rect 81156 78852 81160 78908
rect 81096 78848 81160 78852
rect 81176 78908 81240 78912
rect 81176 78852 81180 78908
rect 81180 78852 81236 78908
rect 81236 78852 81240 78908
rect 81176 78848 81240 78852
rect 81256 78908 81320 78912
rect 81256 78852 81260 78908
rect 81260 78852 81316 78908
rect 81316 78852 81320 78908
rect 81256 78848 81320 78852
rect 111736 78908 111800 78912
rect 111736 78852 111740 78908
rect 111740 78852 111796 78908
rect 111796 78852 111800 78908
rect 111736 78848 111800 78852
rect 111816 78908 111880 78912
rect 111816 78852 111820 78908
rect 111820 78852 111876 78908
rect 111876 78852 111880 78908
rect 111816 78848 111880 78852
rect 111896 78908 111960 78912
rect 111896 78852 111900 78908
rect 111900 78852 111956 78908
rect 111956 78852 111960 78908
rect 111896 78848 111960 78852
rect 111976 78908 112040 78912
rect 111976 78852 111980 78908
rect 111980 78852 112036 78908
rect 112036 78852 112040 78908
rect 111976 78848 112040 78852
rect 142456 78908 142520 78912
rect 142456 78852 142460 78908
rect 142460 78852 142516 78908
rect 142516 78852 142520 78908
rect 142456 78848 142520 78852
rect 142536 78908 142600 78912
rect 142536 78852 142540 78908
rect 142540 78852 142596 78908
rect 142596 78852 142600 78908
rect 142536 78848 142600 78852
rect 142616 78908 142680 78912
rect 142616 78852 142620 78908
rect 142620 78852 142676 78908
rect 142676 78852 142680 78908
rect 142616 78848 142680 78852
rect 142696 78908 142760 78912
rect 142696 78852 142700 78908
rect 142700 78852 142756 78908
rect 142756 78852 142760 78908
rect 142696 78848 142760 78852
rect 173176 78908 173240 78912
rect 173176 78852 173180 78908
rect 173180 78852 173236 78908
rect 173236 78852 173240 78908
rect 173176 78848 173240 78852
rect 173256 78908 173320 78912
rect 173256 78852 173260 78908
rect 173260 78852 173316 78908
rect 173316 78852 173320 78908
rect 173256 78848 173320 78852
rect 173336 78908 173400 78912
rect 173336 78852 173340 78908
rect 173340 78852 173396 78908
rect 173396 78852 173400 78908
rect 173336 78848 173400 78852
rect 173416 78908 173480 78912
rect 173416 78852 173420 78908
rect 173420 78852 173476 78908
rect 173476 78852 173480 78908
rect 173416 78848 173480 78852
rect 4216 78364 4280 78368
rect 4216 78308 4220 78364
rect 4220 78308 4276 78364
rect 4276 78308 4280 78364
rect 4216 78304 4280 78308
rect 4296 78364 4360 78368
rect 4296 78308 4300 78364
rect 4300 78308 4356 78364
rect 4356 78308 4360 78364
rect 4296 78304 4360 78308
rect 4376 78364 4440 78368
rect 4376 78308 4380 78364
rect 4380 78308 4436 78364
rect 4436 78308 4440 78364
rect 4376 78304 4440 78308
rect 4456 78364 4520 78368
rect 4456 78308 4460 78364
rect 4460 78308 4516 78364
rect 4516 78308 4520 78364
rect 4456 78304 4520 78308
rect 34936 78364 35000 78368
rect 34936 78308 34940 78364
rect 34940 78308 34996 78364
rect 34996 78308 35000 78364
rect 34936 78304 35000 78308
rect 35016 78364 35080 78368
rect 35016 78308 35020 78364
rect 35020 78308 35076 78364
rect 35076 78308 35080 78364
rect 35016 78304 35080 78308
rect 35096 78364 35160 78368
rect 35096 78308 35100 78364
rect 35100 78308 35156 78364
rect 35156 78308 35160 78364
rect 35096 78304 35160 78308
rect 35176 78364 35240 78368
rect 35176 78308 35180 78364
rect 35180 78308 35236 78364
rect 35236 78308 35240 78364
rect 35176 78304 35240 78308
rect 65656 78364 65720 78368
rect 65656 78308 65660 78364
rect 65660 78308 65716 78364
rect 65716 78308 65720 78364
rect 65656 78304 65720 78308
rect 65736 78364 65800 78368
rect 65736 78308 65740 78364
rect 65740 78308 65796 78364
rect 65796 78308 65800 78364
rect 65736 78304 65800 78308
rect 65816 78364 65880 78368
rect 65816 78308 65820 78364
rect 65820 78308 65876 78364
rect 65876 78308 65880 78364
rect 65816 78304 65880 78308
rect 65896 78364 65960 78368
rect 65896 78308 65900 78364
rect 65900 78308 65956 78364
rect 65956 78308 65960 78364
rect 65896 78304 65960 78308
rect 96376 78364 96440 78368
rect 96376 78308 96380 78364
rect 96380 78308 96436 78364
rect 96436 78308 96440 78364
rect 96376 78304 96440 78308
rect 96456 78364 96520 78368
rect 96456 78308 96460 78364
rect 96460 78308 96516 78364
rect 96516 78308 96520 78364
rect 96456 78304 96520 78308
rect 96536 78364 96600 78368
rect 96536 78308 96540 78364
rect 96540 78308 96596 78364
rect 96596 78308 96600 78364
rect 96536 78304 96600 78308
rect 96616 78364 96680 78368
rect 96616 78308 96620 78364
rect 96620 78308 96676 78364
rect 96676 78308 96680 78364
rect 96616 78304 96680 78308
rect 127096 78364 127160 78368
rect 127096 78308 127100 78364
rect 127100 78308 127156 78364
rect 127156 78308 127160 78364
rect 127096 78304 127160 78308
rect 127176 78364 127240 78368
rect 127176 78308 127180 78364
rect 127180 78308 127236 78364
rect 127236 78308 127240 78364
rect 127176 78304 127240 78308
rect 127256 78364 127320 78368
rect 127256 78308 127260 78364
rect 127260 78308 127316 78364
rect 127316 78308 127320 78364
rect 127256 78304 127320 78308
rect 127336 78364 127400 78368
rect 127336 78308 127340 78364
rect 127340 78308 127396 78364
rect 127396 78308 127400 78364
rect 127336 78304 127400 78308
rect 157816 78364 157880 78368
rect 157816 78308 157820 78364
rect 157820 78308 157876 78364
rect 157876 78308 157880 78364
rect 157816 78304 157880 78308
rect 157896 78364 157960 78368
rect 157896 78308 157900 78364
rect 157900 78308 157956 78364
rect 157956 78308 157960 78364
rect 157896 78304 157960 78308
rect 157976 78364 158040 78368
rect 157976 78308 157980 78364
rect 157980 78308 158036 78364
rect 158036 78308 158040 78364
rect 157976 78304 158040 78308
rect 158056 78364 158120 78368
rect 158056 78308 158060 78364
rect 158060 78308 158116 78364
rect 158116 78308 158120 78364
rect 158056 78304 158120 78308
rect 19576 77820 19640 77824
rect 19576 77764 19580 77820
rect 19580 77764 19636 77820
rect 19636 77764 19640 77820
rect 19576 77760 19640 77764
rect 19656 77820 19720 77824
rect 19656 77764 19660 77820
rect 19660 77764 19716 77820
rect 19716 77764 19720 77820
rect 19656 77760 19720 77764
rect 19736 77820 19800 77824
rect 19736 77764 19740 77820
rect 19740 77764 19796 77820
rect 19796 77764 19800 77820
rect 19736 77760 19800 77764
rect 19816 77820 19880 77824
rect 19816 77764 19820 77820
rect 19820 77764 19876 77820
rect 19876 77764 19880 77820
rect 19816 77760 19880 77764
rect 50296 77820 50360 77824
rect 50296 77764 50300 77820
rect 50300 77764 50356 77820
rect 50356 77764 50360 77820
rect 50296 77760 50360 77764
rect 50376 77820 50440 77824
rect 50376 77764 50380 77820
rect 50380 77764 50436 77820
rect 50436 77764 50440 77820
rect 50376 77760 50440 77764
rect 50456 77820 50520 77824
rect 50456 77764 50460 77820
rect 50460 77764 50516 77820
rect 50516 77764 50520 77820
rect 50456 77760 50520 77764
rect 50536 77820 50600 77824
rect 50536 77764 50540 77820
rect 50540 77764 50596 77820
rect 50596 77764 50600 77820
rect 50536 77760 50600 77764
rect 81016 77820 81080 77824
rect 81016 77764 81020 77820
rect 81020 77764 81076 77820
rect 81076 77764 81080 77820
rect 81016 77760 81080 77764
rect 81096 77820 81160 77824
rect 81096 77764 81100 77820
rect 81100 77764 81156 77820
rect 81156 77764 81160 77820
rect 81096 77760 81160 77764
rect 81176 77820 81240 77824
rect 81176 77764 81180 77820
rect 81180 77764 81236 77820
rect 81236 77764 81240 77820
rect 81176 77760 81240 77764
rect 81256 77820 81320 77824
rect 81256 77764 81260 77820
rect 81260 77764 81316 77820
rect 81316 77764 81320 77820
rect 81256 77760 81320 77764
rect 111736 77820 111800 77824
rect 111736 77764 111740 77820
rect 111740 77764 111796 77820
rect 111796 77764 111800 77820
rect 111736 77760 111800 77764
rect 111816 77820 111880 77824
rect 111816 77764 111820 77820
rect 111820 77764 111876 77820
rect 111876 77764 111880 77820
rect 111816 77760 111880 77764
rect 111896 77820 111960 77824
rect 111896 77764 111900 77820
rect 111900 77764 111956 77820
rect 111956 77764 111960 77820
rect 111896 77760 111960 77764
rect 111976 77820 112040 77824
rect 111976 77764 111980 77820
rect 111980 77764 112036 77820
rect 112036 77764 112040 77820
rect 111976 77760 112040 77764
rect 142456 77820 142520 77824
rect 142456 77764 142460 77820
rect 142460 77764 142516 77820
rect 142516 77764 142520 77820
rect 142456 77760 142520 77764
rect 142536 77820 142600 77824
rect 142536 77764 142540 77820
rect 142540 77764 142596 77820
rect 142596 77764 142600 77820
rect 142536 77760 142600 77764
rect 142616 77820 142680 77824
rect 142616 77764 142620 77820
rect 142620 77764 142676 77820
rect 142676 77764 142680 77820
rect 142616 77760 142680 77764
rect 142696 77820 142760 77824
rect 142696 77764 142700 77820
rect 142700 77764 142756 77820
rect 142756 77764 142760 77820
rect 142696 77760 142760 77764
rect 173176 77820 173240 77824
rect 173176 77764 173180 77820
rect 173180 77764 173236 77820
rect 173236 77764 173240 77820
rect 173176 77760 173240 77764
rect 173256 77820 173320 77824
rect 173256 77764 173260 77820
rect 173260 77764 173316 77820
rect 173316 77764 173320 77820
rect 173256 77760 173320 77764
rect 173336 77820 173400 77824
rect 173336 77764 173340 77820
rect 173340 77764 173396 77820
rect 173396 77764 173400 77820
rect 173336 77760 173400 77764
rect 173416 77820 173480 77824
rect 173416 77764 173420 77820
rect 173420 77764 173476 77820
rect 173476 77764 173480 77820
rect 173416 77760 173480 77764
rect 4216 77276 4280 77280
rect 4216 77220 4220 77276
rect 4220 77220 4276 77276
rect 4276 77220 4280 77276
rect 4216 77216 4280 77220
rect 4296 77276 4360 77280
rect 4296 77220 4300 77276
rect 4300 77220 4356 77276
rect 4356 77220 4360 77276
rect 4296 77216 4360 77220
rect 4376 77276 4440 77280
rect 4376 77220 4380 77276
rect 4380 77220 4436 77276
rect 4436 77220 4440 77276
rect 4376 77216 4440 77220
rect 4456 77276 4520 77280
rect 4456 77220 4460 77276
rect 4460 77220 4516 77276
rect 4516 77220 4520 77276
rect 4456 77216 4520 77220
rect 34936 77276 35000 77280
rect 34936 77220 34940 77276
rect 34940 77220 34996 77276
rect 34996 77220 35000 77276
rect 34936 77216 35000 77220
rect 35016 77276 35080 77280
rect 35016 77220 35020 77276
rect 35020 77220 35076 77276
rect 35076 77220 35080 77276
rect 35016 77216 35080 77220
rect 35096 77276 35160 77280
rect 35096 77220 35100 77276
rect 35100 77220 35156 77276
rect 35156 77220 35160 77276
rect 35096 77216 35160 77220
rect 35176 77276 35240 77280
rect 35176 77220 35180 77276
rect 35180 77220 35236 77276
rect 35236 77220 35240 77276
rect 35176 77216 35240 77220
rect 65656 77276 65720 77280
rect 65656 77220 65660 77276
rect 65660 77220 65716 77276
rect 65716 77220 65720 77276
rect 65656 77216 65720 77220
rect 65736 77276 65800 77280
rect 65736 77220 65740 77276
rect 65740 77220 65796 77276
rect 65796 77220 65800 77276
rect 65736 77216 65800 77220
rect 65816 77276 65880 77280
rect 65816 77220 65820 77276
rect 65820 77220 65876 77276
rect 65876 77220 65880 77276
rect 65816 77216 65880 77220
rect 65896 77276 65960 77280
rect 65896 77220 65900 77276
rect 65900 77220 65956 77276
rect 65956 77220 65960 77276
rect 65896 77216 65960 77220
rect 96376 77276 96440 77280
rect 96376 77220 96380 77276
rect 96380 77220 96436 77276
rect 96436 77220 96440 77276
rect 96376 77216 96440 77220
rect 96456 77276 96520 77280
rect 96456 77220 96460 77276
rect 96460 77220 96516 77276
rect 96516 77220 96520 77276
rect 96456 77216 96520 77220
rect 96536 77276 96600 77280
rect 96536 77220 96540 77276
rect 96540 77220 96596 77276
rect 96596 77220 96600 77276
rect 96536 77216 96600 77220
rect 96616 77276 96680 77280
rect 96616 77220 96620 77276
rect 96620 77220 96676 77276
rect 96676 77220 96680 77276
rect 96616 77216 96680 77220
rect 127096 77276 127160 77280
rect 127096 77220 127100 77276
rect 127100 77220 127156 77276
rect 127156 77220 127160 77276
rect 127096 77216 127160 77220
rect 127176 77276 127240 77280
rect 127176 77220 127180 77276
rect 127180 77220 127236 77276
rect 127236 77220 127240 77276
rect 127176 77216 127240 77220
rect 127256 77276 127320 77280
rect 127256 77220 127260 77276
rect 127260 77220 127316 77276
rect 127316 77220 127320 77276
rect 127256 77216 127320 77220
rect 127336 77276 127400 77280
rect 127336 77220 127340 77276
rect 127340 77220 127396 77276
rect 127396 77220 127400 77276
rect 127336 77216 127400 77220
rect 157816 77276 157880 77280
rect 157816 77220 157820 77276
rect 157820 77220 157876 77276
rect 157876 77220 157880 77276
rect 157816 77216 157880 77220
rect 157896 77276 157960 77280
rect 157896 77220 157900 77276
rect 157900 77220 157956 77276
rect 157956 77220 157960 77276
rect 157896 77216 157960 77220
rect 157976 77276 158040 77280
rect 157976 77220 157980 77276
rect 157980 77220 158036 77276
rect 158036 77220 158040 77276
rect 157976 77216 158040 77220
rect 158056 77276 158120 77280
rect 158056 77220 158060 77276
rect 158060 77220 158116 77276
rect 158116 77220 158120 77276
rect 158056 77216 158120 77220
rect 19576 76732 19640 76736
rect 19576 76676 19580 76732
rect 19580 76676 19636 76732
rect 19636 76676 19640 76732
rect 19576 76672 19640 76676
rect 19656 76732 19720 76736
rect 19656 76676 19660 76732
rect 19660 76676 19716 76732
rect 19716 76676 19720 76732
rect 19656 76672 19720 76676
rect 19736 76732 19800 76736
rect 19736 76676 19740 76732
rect 19740 76676 19796 76732
rect 19796 76676 19800 76732
rect 19736 76672 19800 76676
rect 19816 76732 19880 76736
rect 19816 76676 19820 76732
rect 19820 76676 19876 76732
rect 19876 76676 19880 76732
rect 19816 76672 19880 76676
rect 50296 76732 50360 76736
rect 50296 76676 50300 76732
rect 50300 76676 50356 76732
rect 50356 76676 50360 76732
rect 50296 76672 50360 76676
rect 50376 76732 50440 76736
rect 50376 76676 50380 76732
rect 50380 76676 50436 76732
rect 50436 76676 50440 76732
rect 50376 76672 50440 76676
rect 50456 76732 50520 76736
rect 50456 76676 50460 76732
rect 50460 76676 50516 76732
rect 50516 76676 50520 76732
rect 50456 76672 50520 76676
rect 50536 76732 50600 76736
rect 50536 76676 50540 76732
rect 50540 76676 50596 76732
rect 50596 76676 50600 76732
rect 50536 76672 50600 76676
rect 81016 76732 81080 76736
rect 81016 76676 81020 76732
rect 81020 76676 81076 76732
rect 81076 76676 81080 76732
rect 81016 76672 81080 76676
rect 81096 76732 81160 76736
rect 81096 76676 81100 76732
rect 81100 76676 81156 76732
rect 81156 76676 81160 76732
rect 81096 76672 81160 76676
rect 81176 76732 81240 76736
rect 81176 76676 81180 76732
rect 81180 76676 81236 76732
rect 81236 76676 81240 76732
rect 81176 76672 81240 76676
rect 81256 76732 81320 76736
rect 81256 76676 81260 76732
rect 81260 76676 81316 76732
rect 81316 76676 81320 76732
rect 81256 76672 81320 76676
rect 111736 76732 111800 76736
rect 111736 76676 111740 76732
rect 111740 76676 111796 76732
rect 111796 76676 111800 76732
rect 111736 76672 111800 76676
rect 111816 76732 111880 76736
rect 111816 76676 111820 76732
rect 111820 76676 111876 76732
rect 111876 76676 111880 76732
rect 111816 76672 111880 76676
rect 111896 76732 111960 76736
rect 111896 76676 111900 76732
rect 111900 76676 111956 76732
rect 111956 76676 111960 76732
rect 111896 76672 111960 76676
rect 111976 76732 112040 76736
rect 111976 76676 111980 76732
rect 111980 76676 112036 76732
rect 112036 76676 112040 76732
rect 111976 76672 112040 76676
rect 142456 76732 142520 76736
rect 142456 76676 142460 76732
rect 142460 76676 142516 76732
rect 142516 76676 142520 76732
rect 142456 76672 142520 76676
rect 142536 76732 142600 76736
rect 142536 76676 142540 76732
rect 142540 76676 142596 76732
rect 142596 76676 142600 76732
rect 142536 76672 142600 76676
rect 142616 76732 142680 76736
rect 142616 76676 142620 76732
rect 142620 76676 142676 76732
rect 142676 76676 142680 76732
rect 142616 76672 142680 76676
rect 142696 76732 142760 76736
rect 142696 76676 142700 76732
rect 142700 76676 142756 76732
rect 142756 76676 142760 76732
rect 142696 76672 142760 76676
rect 173176 76732 173240 76736
rect 173176 76676 173180 76732
rect 173180 76676 173236 76732
rect 173236 76676 173240 76732
rect 173176 76672 173240 76676
rect 173256 76732 173320 76736
rect 173256 76676 173260 76732
rect 173260 76676 173316 76732
rect 173316 76676 173320 76732
rect 173256 76672 173320 76676
rect 173336 76732 173400 76736
rect 173336 76676 173340 76732
rect 173340 76676 173396 76732
rect 173396 76676 173400 76732
rect 173336 76672 173400 76676
rect 173416 76732 173480 76736
rect 173416 76676 173420 76732
rect 173420 76676 173476 76732
rect 173476 76676 173480 76732
rect 173416 76672 173480 76676
rect 4216 76188 4280 76192
rect 4216 76132 4220 76188
rect 4220 76132 4276 76188
rect 4276 76132 4280 76188
rect 4216 76128 4280 76132
rect 4296 76188 4360 76192
rect 4296 76132 4300 76188
rect 4300 76132 4356 76188
rect 4356 76132 4360 76188
rect 4296 76128 4360 76132
rect 4376 76188 4440 76192
rect 4376 76132 4380 76188
rect 4380 76132 4436 76188
rect 4436 76132 4440 76188
rect 4376 76128 4440 76132
rect 4456 76188 4520 76192
rect 4456 76132 4460 76188
rect 4460 76132 4516 76188
rect 4516 76132 4520 76188
rect 4456 76128 4520 76132
rect 34936 76188 35000 76192
rect 34936 76132 34940 76188
rect 34940 76132 34996 76188
rect 34996 76132 35000 76188
rect 34936 76128 35000 76132
rect 35016 76188 35080 76192
rect 35016 76132 35020 76188
rect 35020 76132 35076 76188
rect 35076 76132 35080 76188
rect 35016 76128 35080 76132
rect 35096 76188 35160 76192
rect 35096 76132 35100 76188
rect 35100 76132 35156 76188
rect 35156 76132 35160 76188
rect 35096 76128 35160 76132
rect 35176 76188 35240 76192
rect 35176 76132 35180 76188
rect 35180 76132 35236 76188
rect 35236 76132 35240 76188
rect 35176 76128 35240 76132
rect 65656 76188 65720 76192
rect 65656 76132 65660 76188
rect 65660 76132 65716 76188
rect 65716 76132 65720 76188
rect 65656 76128 65720 76132
rect 65736 76188 65800 76192
rect 65736 76132 65740 76188
rect 65740 76132 65796 76188
rect 65796 76132 65800 76188
rect 65736 76128 65800 76132
rect 65816 76188 65880 76192
rect 65816 76132 65820 76188
rect 65820 76132 65876 76188
rect 65876 76132 65880 76188
rect 65816 76128 65880 76132
rect 65896 76188 65960 76192
rect 65896 76132 65900 76188
rect 65900 76132 65956 76188
rect 65956 76132 65960 76188
rect 65896 76128 65960 76132
rect 96376 76188 96440 76192
rect 96376 76132 96380 76188
rect 96380 76132 96436 76188
rect 96436 76132 96440 76188
rect 96376 76128 96440 76132
rect 96456 76188 96520 76192
rect 96456 76132 96460 76188
rect 96460 76132 96516 76188
rect 96516 76132 96520 76188
rect 96456 76128 96520 76132
rect 96536 76188 96600 76192
rect 96536 76132 96540 76188
rect 96540 76132 96596 76188
rect 96596 76132 96600 76188
rect 96536 76128 96600 76132
rect 96616 76188 96680 76192
rect 96616 76132 96620 76188
rect 96620 76132 96676 76188
rect 96676 76132 96680 76188
rect 96616 76128 96680 76132
rect 127096 76188 127160 76192
rect 127096 76132 127100 76188
rect 127100 76132 127156 76188
rect 127156 76132 127160 76188
rect 127096 76128 127160 76132
rect 127176 76188 127240 76192
rect 127176 76132 127180 76188
rect 127180 76132 127236 76188
rect 127236 76132 127240 76188
rect 127176 76128 127240 76132
rect 127256 76188 127320 76192
rect 127256 76132 127260 76188
rect 127260 76132 127316 76188
rect 127316 76132 127320 76188
rect 127256 76128 127320 76132
rect 127336 76188 127400 76192
rect 127336 76132 127340 76188
rect 127340 76132 127396 76188
rect 127396 76132 127400 76188
rect 127336 76128 127400 76132
rect 157816 76188 157880 76192
rect 157816 76132 157820 76188
rect 157820 76132 157876 76188
rect 157876 76132 157880 76188
rect 157816 76128 157880 76132
rect 157896 76188 157960 76192
rect 157896 76132 157900 76188
rect 157900 76132 157956 76188
rect 157956 76132 157960 76188
rect 157896 76128 157960 76132
rect 157976 76188 158040 76192
rect 157976 76132 157980 76188
rect 157980 76132 158036 76188
rect 158036 76132 158040 76188
rect 157976 76128 158040 76132
rect 158056 76188 158120 76192
rect 158056 76132 158060 76188
rect 158060 76132 158116 76188
rect 158116 76132 158120 76188
rect 158056 76128 158120 76132
rect 19576 75644 19640 75648
rect 19576 75588 19580 75644
rect 19580 75588 19636 75644
rect 19636 75588 19640 75644
rect 19576 75584 19640 75588
rect 19656 75644 19720 75648
rect 19656 75588 19660 75644
rect 19660 75588 19716 75644
rect 19716 75588 19720 75644
rect 19656 75584 19720 75588
rect 19736 75644 19800 75648
rect 19736 75588 19740 75644
rect 19740 75588 19796 75644
rect 19796 75588 19800 75644
rect 19736 75584 19800 75588
rect 19816 75644 19880 75648
rect 19816 75588 19820 75644
rect 19820 75588 19876 75644
rect 19876 75588 19880 75644
rect 19816 75584 19880 75588
rect 50296 75644 50360 75648
rect 50296 75588 50300 75644
rect 50300 75588 50356 75644
rect 50356 75588 50360 75644
rect 50296 75584 50360 75588
rect 50376 75644 50440 75648
rect 50376 75588 50380 75644
rect 50380 75588 50436 75644
rect 50436 75588 50440 75644
rect 50376 75584 50440 75588
rect 50456 75644 50520 75648
rect 50456 75588 50460 75644
rect 50460 75588 50516 75644
rect 50516 75588 50520 75644
rect 50456 75584 50520 75588
rect 50536 75644 50600 75648
rect 50536 75588 50540 75644
rect 50540 75588 50596 75644
rect 50596 75588 50600 75644
rect 50536 75584 50600 75588
rect 81016 75644 81080 75648
rect 81016 75588 81020 75644
rect 81020 75588 81076 75644
rect 81076 75588 81080 75644
rect 81016 75584 81080 75588
rect 81096 75644 81160 75648
rect 81096 75588 81100 75644
rect 81100 75588 81156 75644
rect 81156 75588 81160 75644
rect 81096 75584 81160 75588
rect 81176 75644 81240 75648
rect 81176 75588 81180 75644
rect 81180 75588 81236 75644
rect 81236 75588 81240 75644
rect 81176 75584 81240 75588
rect 81256 75644 81320 75648
rect 81256 75588 81260 75644
rect 81260 75588 81316 75644
rect 81316 75588 81320 75644
rect 81256 75584 81320 75588
rect 111736 75644 111800 75648
rect 111736 75588 111740 75644
rect 111740 75588 111796 75644
rect 111796 75588 111800 75644
rect 111736 75584 111800 75588
rect 111816 75644 111880 75648
rect 111816 75588 111820 75644
rect 111820 75588 111876 75644
rect 111876 75588 111880 75644
rect 111816 75584 111880 75588
rect 111896 75644 111960 75648
rect 111896 75588 111900 75644
rect 111900 75588 111956 75644
rect 111956 75588 111960 75644
rect 111896 75584 111960 75588
rect 111976 75644 112040 75648
rect 111976 75588 111980 75644
rect 111980 75588 112036 75644
rect 112036 75588 112040 75644
rect 111976 75584 112040 75588
rect 142456 75644 142520 75648
rect 142456 75588 142460 75644
rect 142460 75588 142516 75644
rect 142516 75588 142520 75644
rect 142456 75584 142520 75588
rect 142536 75644 142600 75648
rect 142536 75588 142540 75644
rect 142540 75588 142596 75644
rect 142596 75588 142600 75644
rect 142536 75584 142600 75588
rect 142616 75644 142680 75648
rect 142616 75588 142620 75644
rect 142620 75588 142676 75644
rect 142676 75588 142680 75644
rect 142616 75584 142680 75588
rect 142696 75644 142760 75648
rect 142696 75588 142700 75644
rect 142700 75588 142756 75644
rect 142756 75588 142760 75644
rect 142696 75584 142760 75588
rect 173176 75644 173240 75648
rect 173176 75588 173180 75644
rect 173180 75588 173236 75644
rect 173236 75588 173240 75644
rect 173176 75584 173240 75588
rect 173256 75644 173320 75648
rect 173256 75588 173260 75644
rect 173260 75588 173316 75644
rect 173316 75588 173320 75644
rect 173256 75584 173320 75588
rect 173336 75644 173400 75648
rect 173336 75588 173340 75644
rect 173340 75588 173396 75644
rect 173396 75588 173400 75644
rect 173336 75584 173400 75588
rect 173416 75644 173480 75648
rect 173416 75588 173420 75644
rect 173420 75588 173476 75644
rect 173476 75588 173480 75644
rect 173416 75584 173480 75588
rect 4216 75100 4280 75104
rect 4216 75044 4220 75100
rect 4220 75044 4276 75100
rect 4276 75044 4280 75100
rect 4216 75040 4280 75044
rect 4296 75100 4360 75104
rect 4296 75044 4300 75100
rect 4300 75044 4356 75100
rect 4356 75044 4360 75100
rect 4296 75040 4360 75044
rect 4376 75100 4440 75104
rect 4376 75044 4380 75100
rect 4380 75044 4436 75100
rect 4436 75044 4440 75100
rect 4376 75040 4440 75044
rect 4456 75100 4520 75104
rect 4456 75044 4460 75100
rect 4460 75044 4516 75100
rect 4516 75044 4520 75100
rect 4456 75040 4520 75044
rect 34936 75100 35000 75104
rect 34936 75044 34940 75100
rect 34940 75044 34996 75100
rect 34996 75044 35000 75100
rect 34936 75040 35000 75044
rect 35016 75100 35080 75104
rect 35016 75044 35020 75100
rect 35020 75044 35076 75100
rect 35076 75044 35080 75100
rect 35016 75040 35080 75044
rect 35096 75100 35160 75104
rect 35096 75044 35100 75100
rect 35100 75044 35156 75100
rect 35156 75044 35160 75100
rect 35096 75040 35160 75044
rect 35176 75100 35240 75104
rect 35176 75044 35180 75100
rect 35180 75044 35236 75100
rect 35236 75044 35240 75100
rect 35176 75040 35240 75044
rect 65656 75100 65720 75104
rect 65656 75044 65660 75100
rect 65660 75044 65716 75100
rect 65716 75044 65720 75100
rect 65656 75040 65720 75044
rect 65736 75100 65800 75104
rect 65736 75044 65740 75100
rect 65740 75044 65796 75100
rect 65796 75044 65800 75100
rect 65736 75040 65800 75044
rect 65816 75100 65880 75104
rect 65816 75044 65820 75100
rect 65820 75044 65876 75100
rect 65876 75044 65880 75100
rect 65816 75040 65880 75044
rect 65896 75100 65960 75104
rect 65896 75044 65900 75100
rect 65900 75044 65956 75100
rect 65956 75044 65960 75100
rect 65896 75040 65960 75044
rect 96376 75100 96440 75104
rect 96376 75044 96380 75100
rect 96380 75044 96436 75100
rect 96436 75044 96440 75100
rect 96376 75040 96440 75044
rect 96456 75100 96520 75104
rect 96456 75044 96460 75100
rect 96460 75044 96516 75100
rect 96516 75044 96520 75100
rect 96456 75040 96520 75044
rect 96536 75100 96600 75104
rect 96536 75044 96540 75100
rect 96540 75044 96596 75100
rect 96596 75044 96600 75100
rect 96536 75040 96600 75044
rect 96616 75100 96680 75104
rect 96616 75044 96620 75100
rect 96620 75044 96676 75100
rect 96676 75044 96680 75100
rect 96616 75040 96680 75044
rect 127096 75100 127160 75104
rect 127096 75044 127100 75100
rect 127100 75044 127156 75100
rect 127156 75044 127160 75100
rect 127096 75040 127160 75044
rect 127176 75100 127240 75104
rect 127176 75044 127180 75100
rect 127180 75044 127236 75100
rect 127236 75044 127240 75100
rect 127176 75040 127240 75044
rect 127256 75100 127320 75104
rect 127256 75044 127260 75100
rect 127260 75044 127316 75100
rect 127316 75044 127320 75100
rect 127256 75040 127320 75044
rect 127336 75100 127400 75104
rect 127336 75044 127340 75100
rect 127340 75044 127396 75100
rect 127396 75044 127400 75100
rect 127336 75040 127400 75044
rect 157816 75100 157880 75104
rect 157816 75044 157820 75100
rect 157820 75044 157876 75100
rect 157876 75044 157880 75100
rect 157816 75040 157880 75044
rect 157896 75100 157960 75104
rect 157896 75044 157900 75100
rect 157900 75044 157956 75100
rect 157956 75044 157960 75100
rect 157896 75040 157960 75044
rect 157976 75100 158040 75104
rect 157976 75044 157980 75100
rect 157980 75044 158036 75100
rect 158036 75044 158040 75100
rect 157976 75040 158040 75044
rect 158056 75100 158120 75104
rect 158056 75044 158060 75100
rect 158060 75044 158116 75100
rect 158116 75044 158120 75100
rect 158056 75040 158120 75044
rect 19576 74556 19640 74560
rect 19576 74500 19580 74556
rect 19580 74500 19636 74556
rect 19636 74500 19640 74556
rect 19576 74496 19640 74500
rect 19656 74556 19720 74560
rect 19656 74500 19660 74556
rect 19660 74500 19716 74556
rect 19716 74500 19720 74556
rect 19656 74496 19720 74500
rect 19736 74556 19800 74560
rect 19736 74500 19740 74556
rect 19740 74500 19796 74556
rect 19796 74500 19800 74556
rect 19736 74496 19800 74500
rect 19816 74556 19880 74560
rect 19816 74500 19820 74556
rect 19820 74500 19876 74556
rect 19876 74500 19880 74556
rect 19816 74496 19880 74500
rect 50296 74556 50360 74560
rect 50296 74500 50300 74556
rect 50300 74500 50356 74556
rect 50356 74500 50360 74556
rect 50296 74496 50360 74500
rect 50376 74556 50440 74560
rect 50376 74500 50380 74556
rect 50380 74500 50436 74556
rect 50436 74500 50440 74556
rect 50376 74496 50440 74500
rect 50456 74556 50520 74560
rect 50456 74500 50460 74556
rect 50460 74500 50516 74556
rect 50516 74500 50520 74556
rect 50456 74496 50520 74500
rect 50536 74556 50600 74560
rect 50536 74500 50540 74556
rect 50540 74500 50596 74556
rect 50596 74500 50600 74556
rect 50536 74496 50600 74500
rect 81016 74556 81080 74560
rect 81016 74500 81020 74556
rect 81020 74500 81076 74556
rect 81076 74500 81080 74556
rect 81016 74496 81080 74500
rect 81096 74556 81160 74560
rect 81096 74500 81100 74556
rect 81100 74500 81156 74556
rect 81156 74500 81160 74556
rect 81096 74496 81160 74500
rect 81176 74556 81240 74560
rect 81176 74500 81180 74556
rect 81180 74500 81236 74556
rect 81236 74500 81240 74556
rect 81176 74496 81240 74500
rect 81256 74556 81320 74560
rect 81256 74500 81260 74556
rect 81260 74500 81316 74556
rect 81316 74500 81320 74556
rect 81256 74496 81320 74500
rect 111736 74556 111800 74560
rect 111736 74500 111740 74556
rect 111740 74500 111796 74556
rect 111796 74500 111800 74556
rect 111736 74496 111800 74500
rect 111816 74556 111880 74560
rect 111816 74500 111820 74556
rect 111820 74500 111876 74556
rect 111876 74500 111880 74556
rect 111816 74496 111880 74500
rect 111896 74556 111960 74560
rect 111896 74500 111900 74556
rect 111900 74500 111956 74556
rect 111956 74500 111960 74556
rect 111896 74496 111960 74500
rect 111976 74556 112040 74560
rect 111976 74500 111980 74556
rect 111980 74500 112036 74556
rect 112036 74500 112040 74556
rect 111976 74496 112040 74500
rect 142456 74556 142520 74560
rect 142456 74500 142460 74556
rect 142460 74500 142516 74556
rect 142516 74500 142520 74556
rect 142456 74496 142520 74500
rect 142536 74556 142600 74560
rect 142536 74500 142540 74556
rect 142540 74500 142596 74556
rect 142596 74500 142600 74556
rect 142536 74496 142600 74500
rect 142616 74556 142680 74560
rect 142616 74500 142620 74556
rect 142620 74500 142676 74556
rect 142676 74500 142680 74556
rect 142616 74496 142680 74500
rect 142696 74556 142760 74560
rect 142696 74500 142700 74556
rect 142700 74500 142756 74556
rect 142756 74500 142760 74556
rect 142696 74496 142760 74500
rect 173176 74556 173240 74560
rect 173176 74500 173180 74556
rect 173180 74500 173236 74556
rect 173236 74500 173240 74556
rect 173176 74496 173240 74500
rect 173256 74556 173320 74560
rect 173256 74500 173260 74556
rect 173260 74500 173316 74556
rect 173316 74500 173320 74556
rect 173256 74496 173320 74500
rect 173336 74556 173400 74560
rect 173336 74500 173340 74556
rect 173340 74500 173396 74556
rect 173396 74500 173400 74556
rect 173336 74496 173400 74500
rect 173416 74556 173480 74560
rect 173416 74500 173420 74556
rect 173420 74500 173476 74556
rect 173476 74500 173480 74556
rect 173416 74496 173480 74500
rect 4216 74012 4280 74016
rect 4216 73956 4220 74012
rect 4220 73956 4276 74012
rect 4276 73956 4280 74012
rect 4216 73952 4280 73956
rect 4296 74012 4360 74016
rect 4296 73956 4300 74012
rect 4300 73956 4356 74012
rect 4356 73956 4360 74012
rect 4296 73952 4360 73956
rect 4376 74012 4440 74016
rect 4376 73956 4380 74012
rect 4380 73956 4436 74012
rect 4436 73956 4440 74012
rect 4376 73952 4440 73956
rect 4456 74012 4520 74016
rect 4456 73956 4460 74012
rect 4460 73956 4516 74012
rect 4516 73956 4520 74012
rect 4456 73952 4520 73956
rect 34936 74012 35000 74016
rect 34936 73956 34940 74012
rect 34940 73956 34996 74012
rect 34996 73956 35000 74012
rect 34936 73952 35000 73956
rect 35016 74012 35080 74016
rect 35016 73956 35020 74012
rect 35020 73956 35076 74012
rect 35076 73956 35080 74012
rect 35016 73952 35080 73956
rect 35096 74012 35160 74016
rect 35096 73956 35100 74012
rect 35100 73956 35156 74012
rect 35156 73956 35160 74012
rect 35096 73952 35160 73956
rect 35176 74012 35240 74016
rect 35176 73956 35180 74012
rect 35180 73956 35236 74012
rect 35236 73956 35240 74012
rect 35176 73952 35240 73956
rect 65656 74012 65720 74016
rect 65656 73956 65660 74012
rect 65660 73956 65716 74012
rect 65716 73956 65720 74012
rect 65656 73952 65720 73956
rect 65736 74012 65800 74016
rect 65736 73956 65740 74012
rect 65740 73956 65796 74012
rect 65796 73956 65800 74012
rect 65736 73952 65800 73956
rect 65816 74012 65880 74016
rect 65816 73956 65820 74012
rect 65820 73956 65876 74012
rect 65876 73956 65880 74012
rect 65816 73952 65880 73956
rect 65896 74012 65960 74016
rect 65896 73956 65900 74012
rect 65900 73956 65956 74012
rect 65956 73956 65960 74012
rect 65896 73952 65960 73956
rect 96376 74012 96440 74016
rect 96376 73956 96380 74012
rect 96380 73956 96436 74012
rect 96436 73956 96440 74012
rect 96376 73952 96440 73956
rect 96456 74012 96520 74016
rect 96456 73956 96460 74012
rect 96460 73956 96516 74012
rect 96516 73956 96520 74012
rect 96456 73952 96520 73956
rect 96536 74012 96600 74016
rect 96536 73956 96540 74012
rect 96540 73956 96596 74012
rect 96596 73956 96600 74012
rect 96536 73952 96600 73956
rect 96616 74012 96680 74016
rect 96616 73956 96620 74012
rect 96620 73956 96676 74012
rect 96676 73956 96680 74012
rect 96616 73952 96680 73956
rect 127096 74012 127160 74016
rect 127096 73956 127100 74012
rect 127100 73956 127156 74012
rect 127156 73956 127160 74012
rect 127096 73952 127160 73956
rect 127176 74012 127240 74016
rect 127176 73956 127180 74012
rect 127180 73956 127236 74012
rect 127236 73956 127240 74012
rect 127176 73952 127240 73956
rect 127256 74012 127320 74016
rect 127256 73956 127260 74012
rect 127260 73956 127316 74012
rect 127316 73956 127320 74012
rect 127256 73952 127320 73956
rect 127336 74012 127400 74016
rect 127336 73956 127340 74012
rect 127340 73956 127396 74012
rect 127396 73956 127400 74012
rect 127336 73952 127400 73956
rect 157816 74012 157880 74016
rect 157816 73956 157820 74012
rect 157820 73956 157876 74012
rect 157876 73956 157880 74012
rect 157816 73952 157880 73956
rect 157896 74012 157960 74016
rect 157896 73956 157900 74012
rect 157900 73956 157956 74012
rect 157956 73956 157960 74012
rect 157896 73952 157960 73956
rect 157976 74012 158040 74016
rect 157976 73956 157980 74012
rect 157980 73956 158036 74012
rect 158036 73956 158040 74012
rect 157976 73952 158040 73956
rect 158056 74012 158120 74016
rect 158056 73956 158060 74012
rect 158060 73956 158116 74012
rect 158116 73956 158120 74012
rect 158056 73952 158120 73956
rect 19576 73468 19640 73472
rect 19576 73412 19580 73468
rect 19580 73412 19636 73468
rect 19636 73412 19640 73468
rect 19576 73408 19640 73412
rect 19656 73468 19720 73472
rect 19656 73412 19660 73468
rect 19660 73412 19716 73468
rect 19716 73412 19720 73468
rect 19656 73408 19720 73412
rect 19736 73468 19800 73472
rect 19736 73412 19740 73468
rect 19740 73412 19796 73468
rect 19796 73412 19800 73468
rect 19736 73408 19800 73412
rect 19816 73468 19880 73472
rect 19816 73412 19820 73468
rect 19820 73412 19876 73468
rect 19876 73412 19880 73468
rect 19816 73408 19880 73412
rect 50296 73468 50360 73472
rect 50296 73412 50300 73468
rect 50300 73412 50356 73468
rect 50356 73412 50360 73468
rect 50296 73408 50360 73412
rect 50376 73468 50440 73472
rect 50376 73412 50380 73468
rect 50380 73412 50436 73468
rect 50436 73412 50440 73468
rect 50376 73408 50440 73412
rect 50456 73468 50520 73472
rect 50456 73412 50460 73468
rect 50460 73412 50516 73468
rect 50516 73412 50520 73468
rect 50456 73408 50520 73412
rect 50536 73468 50600 73472
rect 50536 73412 50540 73468
rect 50540 73412 50596 73468
rect 50596 73412 50600 73468
rect 50536 73408 50600 73412
rect 81016 73468 81080 73472
rect 81016 73412 81020 73468
rect 81020 73412 81076 73468
rect 81076 73412 81080 73468
rect 81016 73408 81080 73412
rect 81096 73468 81160 73472
rect 81096 73412 81100 73468
rect 81100 73412 81156 73468
rect 81156 73412 81160 73468
rect 81096 73408 81160 73412
rect 81176 73468 81240 73472
rect 81176 73412 81180 73468
rect 81180 73412 81236 73468
rect 81236 73412 81240 73468
rect 81176 73408 81240 73412
rect 81256 73468 81320 73472
rect 81256 73412 81260 73468
rect 81260 73412 81316 73468
rect 81316 73412 81320 73468
rect 81256 73408 81320 73412
rect 111736 73468 111800 73472
rect 111736 73412 111740 73468
rect 111740 73412 111796 73468
rect 111796 73412 111800 73468
rect 111736 73408 111800 73412
rect 111816 73468 111880 73472
rect 111816 73412 111820 73468
rect 111820 73412 111876 73468
rect 111876 73412 111880 73468
rect 111816 73408 111880 73412
rect 111896 73468 111960 73472
rect 111896 73412 111900 73468
rect 111900 73412 111956 73468
rect 111956 73412 111960 73468
rect 111896 73408 111960 73412
rect 111976 73468 112040 73472
rect 111976 73412 111980 73468
rect 111980 73412 112036 73468
rect 112036 73412 112040 73468
rect 111976 73408 112040 73412
rect 142456 73468 142520 73472
rect 142456 73412 142460 73468
rect 142460 73412 142516 73468
rect 142516 73412 142520 73468
rect 142456 73408 142520 73412
rect 142536 73468 142600 73472
rect 142536 73412 142540 73468
rect 142540 73412 142596 73468
rect 142596 73412 142600 73468
rect 142536 73408 142600 73412
rect 142616 73468 142680 73472
rect 142616 73412 142620 73468
rect 142620 73412 142676 73468
rect 142676 73412 142680 73468
rect 142616 73408 142680 73412
rect 142696 73468 142760 73472
rect 142696 73412 142700 73468
rect 142700 73412 142756 73468
rect 142756 73412 142760 73468
rect 142696 73408 142760 73412
rect 173176 73468 173240 73472
rect 173176 73412 173180 73468
rect 173180 73412 173236 73468
rect 173236 73412 173240 73468
rect 173176 73408 173240 73412
rect 173256 73468 173320 73472
rect 173256 73412 173260 73468
rect 173260 73412 173316 73468
rect 173316 73412 173320 73468
rect 173256 73408 173320 73412
rect 173336 73468 173400 73472
rect 173336 73412 173340 73468
rect 173340 73412 173396 73468
rect 173396 73412 173400 73468
rect 173336 73408 173400 73412
rect 173416 73468 173480 73472
rect 173416 73412 173420 73468
rect 173420 73412 173476 73468
rect 173476 73412 173480 73468
rect 173416 73408 173480 73412
rect 4216 72924 4280 72928
rect 4216 72868 4220 72924
rect 4220 72868 4276 72924
rect 4276 72868 4280 72924
rect 4216 72864 4280 72868
rect 4296 72924 4360 72928
rect 4296 72868 4300 72924
rect 4300 72868 4356 72924
rect 4356 72868 4360 72924
rect 4296 72864 4360 72868
rect 4376 72924 4440 72928
rect 4376 72868 4380 72924
rect 4380 72868 4436 72924
rect 4436 72868 4440 72924
rect 4376 72864 4440 72868
rect 4456 72924 4520 72928
rect 4456 72868 4460 72924
rect 4460 72868 4516 72924
rect 4516 72868 4520 72924
rect 4456 72864 4520 72868
rect 34936 72924 35000 72928
rect 34936 72868 34940 72924
rect 34940 72868 34996 72924
rect 34996 72868 35000 72924
rect 34936 72864 35000 72868
rect 35016 72924 35080 72928
rect 35016 72868 35020 72924
rect 35020 72868 35076 72924
rect 35076 72868 35080 72924
rect 35016 72864 35080 72868
rect 35096 72924 35160 72928
rect 35096 72868 35100 72924
rect 35100 72868 35156 72924
rect 35156 72868 35160 72924
rect 35096 72864 35160 72868
rect 35176 72924 35240 72928
rect 35176 72868 35180 72924
rect 35180 72868 35236 72924
rect 35236 72868 35240 72924
rect 35176 72864 35240 72868
rect 65656 72924 65720 72928
rect 65656 72868 65660 72924
rect 65660 72868 65716 72924
rect 65716 72868 65720 72924
rect 65656 72864 65720 72868
rect 65736 72924 65800 72928
rect 65736 72868 65740 72924
rect 65740 72868 65796 72924
rect 65796 72868 65800 72924
rect 65736 72864 65800 72868
rect 65816 72924 65880 72928
rect 65816 72868 65820 72924
rect 65820 72868 65876 72924
rect 65876 72868 65880 72924
rect 65816 72864 65880 72868
rect 65896 72924 65960 72928
rect 65896 72868 65900 72924
rect 65900 72868 65956 72924
rect 65956 72868 65960 72924
rect 65896 72864 65960 72868
rect 96376 72924 96440 72928
rect 96376 72868 96380 72924
rect 96380 72868 96436 72924
rect 96436 72868 96440 72924
rect 96376 72864 96440 72868
rect 96456 72924 96520 72928
rect 96456 72868 96460 72924
rect 96460 72868 96516 72924
rect 96516 72868 96520 72924
rect 96456 72864 96520 72868
rect 96536 72924 96600 72928
rect 96536 72868 96540 72924
rect 96540 72868 96596 72924
rect 96596 72868 96600 72924
rect 96536 72864 96600 72868
rect 96616 72924 96680 72928
rect 96616 72868 96620 72924
rect 96620 72868 96676 72924
rect 96676 72868 96680 72924
rect 96616 72864 96680 72868
rect 127096 72924 127160 72928
rect 127096 72868 127100 72924
rect 127100 72868 127156 72924
rect 127156 72868 127160 72924
rect 127096 72864 127160 72868
rect 127176 72924 127240 72928
rect 127176 72868 127180 72924
rect 127180 72868 127236 72924
rect 127236 72868 127240 72924
rect 127176 72864 127240 72868
rect 127256 72924 127320 72928
rect 127256 72868 127260 72924
rect 127260 72868 127316 72924
rect 127316 72868 127320 72924
rect 127256 72864 127320 72868
rect 127336 72924 127400 72928
rect 127336 72868 127340 72924
rect 127340 72868 127396 72924
rect 127396 72868 127400 72924
rect 127336 72864 127400 72868
rect 157816 72924 157880 72928
rect 157816 72868 157820 72924
rect 157820 72868 157876 72924
rect 157876 72868 157880 72924
rect 157816 72864 157880 72868
rect 157896 72924 157960 72928
rect 157896 72868 157900 72924
rect 157900 72868 157956 72924
rect 157956 72868 157960 72924
rect 157896 72864 157960 72868
rect 157976 72924 158040 72928
rect 157976 72868 157980 72924
rect 157980 72868 158036 72924
rect 158036 72868 158040 72924
rect 157976 72864 158040 72868
rect 158056 72924 158120 72928
rect 158056 72868 158060 72924
rect 158060 72868 158116 72924
rect 158116 72868 158120 72924
rect 158056 72864 158120 72868
rect 19576 72380 19640 72384
rect 19576 72324 19580 72380
rect 19580 72324 19636 72380
rect 19636 72324 19640 72380
rect 19576 72320 19640 72324
rect 19656 72380 19720 72384
rect 19656 72324 19660 72380
rect 19660 72324 19716 72380
rect 19716 72324 19720 72380
rect 19656 72320 19720 72324
rect 19736 72380 19800 72384
rect 19736 72324 19740 72380
rect 19740 72324 19796 72380
rect 19796 72324 19800 72380
rect 19736 72320 19800 72324
rect 19816 72380 19880 72384
rect 19816 72324 19820 72380
rect 19820 72324 19876 72380
rect 19876 72324 19880 72380
rect 19816 72320 19880 72324
rect 50296 72380 50360 72384
rect 50296 72324 50300 72380
rect 50300 72324 50356 72380
rect 50356 72324 50360 72380
rect 50296 72320 50360 72324
rect 50376 72380 50440 72384
rect 50376 72324 50380 72380
rect 50380 72324 50436 72380
rect 50436 72324 50440 72380
rect 50376 72320 50440 72324
rect 50456 72380 50520 72384
rect 50456 72324 50460 72380
rect 50460 72324 50516 72380
rect 50516 72324 50520 72380
rect 50456 72320 50520 72324
rect 50536 72380 50600 72384
rect 50536 72324 50540 72380
rect 50540 72324 50596 72380
rect 50596 72324 50600 72380
rect 50536 72320 50600 72324
rect 81016 72380 81080 72384
rect 81016 72324 81020 72380
rect 81020 72324 81076 72380
rect 81076 72324 81080 72380
rect 81016 72320 81080 72324
rect 81096 72380 81160 72384
rect 81096 72324 81100 72380
rect 81100 72324 81156 72380
rect 81156 72324 81160 72380
rect 81096 72320 81160 72324
rect 81176 72380 81240 72384
rect 81176 72324 81180 72380
rect 81180 72324 81236 72380
rect 81236 72324 81240 72380
rect 81176 72320 81240 72324
rect 81256 72380 81320 72384
rect 81256 72324 81260 72380
rect 81260 72324 81316 72380
rect 81316 72324 81320 72380
rect 81256 72320 81320 72324
rect 111736 72380 111800 72384
rect 111736 72324 111740 72380
rect 111740 72324 111796 72380
rect 111796 72324 111800 72380
rect 111736 72320 111800 72324
rect 111816 72380 111880 72384
rect 111816 72324 111820 72380
rect 111820 72324 111876 72380
rect 111876 72324 111880 72380
rect 111816 72320 111880 72324
rect 111896 72380 111960 72384
rect 111896 72324 111900 72380
rect 111900 72324 111956 72380
rect 111956 72324 111960 72380
rect 111896 72320 111960 72324
rect 111976 72380 112040 72384
rect 111976 72324 111980 72380
rect 111980 72324 112036 72380
rect 112036 72324 112040 72380
rect 111976 72320 112040 72324
rect 142456 72380 142520 72384
rect 142456 72324 142460 72380
rect 142460 72324 142516 72380
rect 142516 72324 142520 72380
rect 142456 72320 142520 72324
rect 142536 72380 142600 72384
rect 142536 72324 142540 72380
rect 142540 72324 142596 72380
rect 142596 72324 142600 72380
rect 142536 72320 142600 72324
rect 142616 72380 142680 72384
rect 142616 72324 142620 72380
rect 142620 72324 142676 72380
rect 142676 72324 142680 72380
rect 142616 72320 142680 72324
rect 142696 72380 142760 72384
rect 142696 72324 142700 72380
rect 142700 72324 142756 72380
rect 142756 72324 142760 72380
rect 142696 72320 142760 72324
rect 173176 72380 173240 72384
rect 173176 72324 173180 72380
rect 173180 72324 173236 72380
rect 173236 72324 173240 72380
rect 173176 72320 173240 72324
rect 173256 72380 173320 72384
rect 173256 72324 173260 72380
rect 173260 72324 173316 72380
rect 173316 72324 173320 72380
rect 173256 72320 173320 72324
rect 173336 72380 173400 72384
rect 173336 72324 173340 72380
rect 173340 72324 173396 72380
rect 173396 72324 173400 72380
rect 173336 72320 173400 72324
rect 173416 72380 173480 72384
rect 173416 72324 173420 72380
rect 173420 72324 173476 72380
rect 173476 72324 173480 72380
rect 173416 72320 173480 72324
rect 4216 71836 4280 71840
rect 4216 71780 4220 71836
rect 4220 71780 4276 71836
rect 4276 71780 4280 71836
rect 4216 71776 4280 71780
rect 4296 71836 4360 71840
rect 4296 71780 4300 71836
rect 4300 71780 4356 71836
rect 4356 71780 4360 71836
rect 4296 71776 4360 71780
rect 4376 71836 4440 71840
rect 4376 71780 4380 71836
rect 4380 71780 4436 71836
rect 4436 71780 4440 71836
rect 4376 71776 4440 71780
rect 4456 71836 4520 71840
rect 4456 71780 4460 71836
rect 4460 71780 4516 71836
rect 4516 71780 4520 71836
rect 4456 71776 4520 71780
rect 34936 71836 35000 71840
rect 34936 71780 34940 71836
rect 34940 71780 34996 71836
rect 34996 71780 35000 71836
rect 34936 71776 35000 71780
rect 35016 71836 35080 71840
rect 35016 71780 35020 71836
rect 35020 71780 35076 71836
rect 35076 71780 35080 71836
rect 35016 71776 35080 71780
rect 35096 71836 35160 71840
rect 35096 71780 35100 71836
rect 35100 71780 35156 71836
rect 35156 71780 35160 71836
rect 35096 71776 35160 71780
rect 35176 71836 35240 71840
rect 35176 71780 35180 71836
rect 35180 71780 35236 71836
rect 35236 71780 35240 71836
rect 35176 71776 35240 71780
rect 65656 71836 65720 71840
rect 65656 71780 65660 71836
rect 65660 71780 65716 71836
rect 65716 71780 65720 71836
rect 65656 71776 65720 71780
rect 65736 71836 65800 71840
rect 65736 71780 65740 71836
rect 65740 71780 65796 71836
rect 65796 71780 65800 71836
rect 65736 71776 65800 71780
rect 65816 71836 65880 71840
rect 65816 71780 65820 71836
rect 65820 71780 65876 71836
rect 65876 71780 65880 71836
rect 65816 71776 65880 71780
rect 65896 71836 65960 71840
rect 65896 71780 65900 71836
rect 65900 71780 65956 71836
rect 65956 71780 65960 71836
rect 65896 71776 65960 71780
rect 96376 71836 96440 71840
rect 96376 71780 96380 71836
rect 96380 71780 96436 71836
rect 96436 71780 96440 71836
rect 96376 71776 96440 71780
rect 96456 71836 96520 71840
rect 96456 71780 96460 71836
rect 96460 71780 96516 71836
rect 96516 71780 96520 71836
rect 96456 71776 96520 71780
rect 96536 71836 96600 71840
rect 96536 71780 96540 71836
rect 96540 71780 96596 71836
rect 96596 71780 96600 71836
rect 96536 71776 96600 71780
rect 96616 71836 96680 71840
rect 96616 71780 96620 71836
rect 96620 71780 96676 71836
rect 96676 71780 96680 71836
rect 96616 71776 96680 71780
rect 127096 71836 127160 71840
rect 127096 71780 127100 71836
rect 127100 71780 127156 71836
rect 127156 71780 127160 71836
rect 127096 71776 127160 71780
rect 127176 71836 127240 71840
rect 127176 71780 127180 71836
rect 127180 71780 127236 71836
rect 127236 71780 127240 71836
rect 127176 71776 127240 71780
rect 127256 71836 127320 71840
rect 127256 71780 127260 71836
rect 127260 71780 127316 71836
rect 127316 71780 127320 71836
rect 127256 71776 127320 71780
rect 127336 71836 127400 71840
rect 127336 71780 127340 71836
rect 127340 71780 127396 71836
rect 127396 71780 127400 71836
rect 127336 71776 127400 71780
rect 157816 71836 157880 71840
rect 157816 71780 157820 71836
rect 157820 71780 157876 71836
rect 157876 71780 157880 71836
rect 157816 71776 157880 71780
rect 157896 71836 157960 71840
rect 157896 71780 157900 71836
rect 157900 71780 157956 71836
rect 157956 71780 157960 71836
rect 157896 71776 157960 71780
rect 157976 71836 158040 71840
rect 157976 71780 157980 71836
rect 157980 71780 158036 71836
rect 158036 71780 158040 71836
rect 157976 71776 158040 71780
rect 158056 71836 158120 71840
rect 158056 71780 158060 71836
rect 158060 71780 158116 71836
rect 158116 71780 158120 71836
rect 158056 71776 158120 71780
rect 19576 71292 19640 71296
rect 19576 71236 19580 71292
rect 19580 71236 19636 71292
rect 19636 71236 19640 71292
rect 19576 71232 19640 71236
rect 19656 71292 19720 71296
rect 19656 71236 19660 71292
rect 19660 71236 19716 71292
rect 19716 71236 19720 71292
rect 19656 71232 19720 71236
rect 19736 71292 19800 71296
rect 19736 71236 19740 71292
rect 19740 71236 19796 71292
rect 19796 71236 19800 71292
rect 19736 71232 19800 71236
rect 19816 71292 19880 71296
rect 19816 71236 19820 71292
rect 19820 71236 19876 71292
rect 19876 71236 19880 71292
rect 19816 71232 19880 71236
rect 50296 71292 50360 71296
rect 50296 71236 50300 71292
rect 50300 71236 50356 71292
rect 50356 71236 50360 71292
rect 50296 71232 50360 71236
rect 50376 71292 50440 71296
rect 50376 71236 50380 71292
rect 50380 71236 50436 71292
rect 50436 71236 50440 71292
rect 50376 71232 50440 71236
rect 50456 71292 50520 71296
rect 50456 71236 50460 71292
rect 50460 71236 50516 71292
rect 50516 71236 50520 71292
rect 50456 71232 50520 71236
rect 50536 71292 50600 71296
rect 50536 71236 50540 71292
rect 50540 71236 50596 71292
rect 50596 71236 50600 71292
rect 50536 71232 50600 71236
rect 81016 71292 81080 71296
rect 81016 71236 81020 71292
rect 81020 71236 81076 71292
rect 81076 71236 81080 71292
rect 81016 71232 81080 71236
rect 81096 71292 81160 71296
rect 81096 71236 81100 71292
rect 81100 71236 81156 71292
rect 81156 71236 81160 71292
rect 81096 71232 81160 71236
rect 81176 71292 81240 71296
rect 81176 71236 81180 71292
rect 81180 71236 81236 71292
rect 81236 71236 81240 71292
rect 81176 71232 81240 71236
rect 81256 71292 81320 71296
rect 81256 71236 81260 71292
rect 81260 71236 81316 71292
rect 81316 71236 81320 71292
rect 81256 71232 81320 71236
rect 111736 71292 111800 71296
rect 111736 71236 111740 71292
rect 111740 71236 111796 71292
rect 111796 71236 111800 71292
rect 111736 71232 111800 71236
rect 111816 71292 111880 71296
rect 111816 71236 111820 71292
rect 111820 71236 111876 71292
rect 111876 71236 111880 71292
rect 111816 71232 111880 71236
rect 111896 71292 111960 71296
rect 111896 71236 111900 71292
rect 111900 71236 111956 71292
rect 111956 71236 111960 71292
rect 111896 71232 111960 71236
rect 111976 71292 112040 71296
rect 111976 71236 111980 71292
rect 111980 71236 112036 71292
rect 112036 71236 112040 71292
rect 111976 71232 112040 71236
rect 142456 71292 142520 71296
rect 142456 71236 142460 71292
rect 142460 71236 142516 71292
rect 142516 71236 142520 71292
rect 142456 71232 142520 71236
rect 142536 71292 142600 71296
rect 142536 71236 142540 71292
rect 142540 71236 142596 71292
rect 142596 71236 142600 71292
rect 142536 71232 142600 71236
rect 142616 71292 142680 71296
rect 142616 71236 142620 71292
rect 142620 71236 142676 71292
rect 142676 71236 142680 71292
rect 142616 71232 142680 71236
rect 142696 71292 142760 71296
rect 142696 71236 142700 71292
rect 142700 71236 142756 71292
rect 142756 71236 142760 71292
rect 142696 71232 142760 71236
rect 173176 71292 173240 71296
rect 173176 71236 173180 71292
rect 173180 71236 173236 71292
rect 173236 71236 173240 71292
rect 173176 71232 173240 71236
rect 173256 71292 173320 71296
rect 173256 71236 173260 71292
rect 173260 71236 173316 71292
rect 173316 71236 173320 71292
rect 173256 71232 173320 71236
rect 173336 71292 173400 71296
rect 173336 71236 173340 71292
rect 173340 71236 173396 71292
rect 173396 71236 173400 71292
rect 173336 71232 173400 71236
rect 173416 71292 173480 71296
rect 173416 71236 173420 71292
rect 173420 71236 173476 71292
rect 173476 71236 173480 71292
rect 173416 71232 173480 71236
rect 4216 70748 4280 70752
rect 4216 70692 4220 70748
rect 4220 70692 4276 70748
rect 4276 70692 4280 70748
rect 4216 70688 4280 70692
rect 4296 70748 4360 70752
rect 4296 70692 4300 70748
rect 4300 70692 4356 70748
rect 4356 70692 4360 70748
rect 4296 70688 4360 70692
rect 4376 70748 4440 70752
rect 4376 70692 4380 70748
rect 4380 70692 4436 70748
rect 4436 70692 4440 70748
rect 4376 70688 4440 70692
rect 4456 70748 4520 70752
rect 4456 70692 4460 70748
rect 4460 70692 4516 70748
rect 4516 70692 4520 70748
rect 4456 70688 4520 70692
rect 34936 70748 35000 70752
rect 34936 70692 34940 70748
rect 34940 70692 34996 70748
rect 34996 70692 35000 70748
rect 34936 70688 35000 70692
rect 35016 70748 35080 70752
rect 35016 70692 35020 70748
rect 35020 70692 35076 70748
rect 35076 70692 35080 70748
rect 35016 70688 35080 70692
rect 35096 70748 35160 70752
rect 35096 70692 35100 70748
rect 35100 70692 35156 70748
rect 35156 70692 35160 70748
rect 35096 70688 35160 70692
rect 35176 70748 35240 70752
rect 35176 70692 35180 70748
rect 35180 70692 35236 70748
rect 35236 70692 35240 70748
rect 35176 70688 35240 70692
rect 65656 70748 65720 70752
rect 65656 70692 65660 70748
rect 65660 70692 65716 70748
rect 65716 70692 65720 70748
rect 65656 70688 65720 70692
rect 65736 70748 65800 70752
rect 65736 70692 65740 70748
rect 65740 70692 65796 70748
rect 65796 70692 65800 70748
rect 65736 70688 65800 70692
rect 65816 70748 65880 70752
rect 65816 70692 65820 70748
rect 65820 70692 65876 70748
rect 65876 70692 65880 70748
rect 65816 70688 65880 70692
rect 65896 70748 65960 70752
rect 65896 70692 65900 70748
rect 65900 70692 65956 70748
rect 65956 70692 65960 70748
rect 65896 70688 65960 70692
rect 96376 70748 96440 70752
rect 96376 70692 96380 70748
rect 96380 70692 96436 70748
rect 96436 70692 96440 70748
rect 96376 70688 96440 70692
rect 96456 70748 96520 70752
rect 96456 70692 96460 70748
rect 96460 70692 96516 70748
rect 96516 70692 96520 70748
rect 96456 70688 96520 70692
rect 96536 70748 96600 70752
rect 96536 70692 96540 70748
rect 96540 70692 96596 70748
rect 96596 70692 96600 70748
rect 96536 70688 96600 70692
rect 96616 70748 96680 70752
rect 96616 70692 96620 70748
rect 96620 70692 96676 70748
rect 96676 70692 96680 70748
rect 96616 70688 96680 70692
rect 127096 70748 127160 70752
rect 127096 70692 127100 70748
rect 127100 70692 127156 70748
rect 127156 70692 127160 70748
rect 127096 70688 127160 70692
rect 127176 70748 127240 70752
rect 127176 70692 127180 70748
rect 127180 70692 127236 70748
rect 127236 70692 127240 70748
rect 127176 70688 127240 70692
rect 127256 70748 127320 70752
rect 127256 70692 127260 70748
rect 127260 70692 127316 70748
rect 127316 70692 127320 70748
rect 127256 70688 127320 70692
rect 127336 70748 127400 70752
rect 127336 70692 127340 70748
rect 127340 70692 127396 70748
rect 127396 70692 127400 70748
rect 127336 70688 127400 70692
rect 157816 70748 157880 70752
rect 157816 70692 157820 70748
rect 157820 70692 157876 70748
rect 157876 70692 157880 70748
rect 157816 70688 157880 70692
rect 157896 70748 157960 70752
rect 157896 70692 157900 70748
rect 157900 70692 157956 70748
rect 157956 70692 157960 70748
rect 157896 70688 157960 70692
rect 157976 70748 158040 70752
rect 157976 70692 157980 70748
rect 157980 70692 158036 70748
rect 158036 70692 158040 70748
rect 157976 70688 158040 70692
rect 158056 70748 158120 70752
rect 158056 70692 158060 70748
rect 158060 70692 158116 70748
rect 158116 70692 158120 70748
rect 158056 70688 158120 70692
rect 19576 70204 19640 70208
rect 19576 70148 19580 70204
rect 19580 70148 19636 70204
rect 19636 70148 19640 70204
rect 19576 70144 19640 70148
rect 19656 70204 19720 70208
rect 19656 70148 19660 70204
rect 19660 70148 19716 70204
rect 19716 70148 19720 70204
rect 19656 70144 19720 70148
rect 19736 70204 19800 70208
rect 19736 70148 19740 70204
rect 19740 70148 19796 70204
rect 19796 70148 19800 70204
rect 19736 70144 19800 70148
rect 19816 70204 19880 70208
rect 19816 70148 19820 70204
rect 19820 70148 19876 70204
rect 19876 70148 19880 70204
rect 19816 70144 19880 70148
rect 50296 70204 50360 70208
rect 50296 70148 50300 70204
rect 50300 70148 50356 70204
rect 50356 70148 50360 70204
rect 50296 70144 50360 70148
rect 50376 70204 50440 70208
rect 50376 70148 50380 70204
rect 50380 70148 50436 70204
rect 50436 70148 50440 70204
rect 50376 70144 50440 70148
rect 50456 70204 50520 70208
rect 50456 70148 50460 70204
rect 50460 70148 50516 70204
rect 50516 70148 50520 70204
rect 50456 70144 50520 70148
rect 50536 70204 50600 70208
rect 50536 70148 50540 70204
rect 50540 70148 50596 70204
rect 50596 70148 50600 70204
rect 50536 70144 50600 70148
rect 81016 70204 81080 70208
rect 81016 70148 81020 70204
rect 81020 70148 81076 70204
rect 81076 70148 81080 70204
rect 81016 70144 81080 70148
rect 81096 70204 81160 70208
rect 81096 70148 81100 70204
rect 81100 70148 81156 70204
rect 81156 70148 81160 70204
rect 81096 70144 81160 70148
rect 81176 70204 81240 70208
rect 81176 70148 81180 70204
rect 81180 70148 81236 70204
rect 81236 70148 81240 70204
rect 81176 70144 81240 70148
rect 81256 70204 81320 70208
rect 81256 70148 81260 70204
rect 81260 70148 81316 70204
rect 81316 70148 81320 70204
rect 81256 70144 81320 70148
rect 111736 70204 111800 70208
rect 111736 70148 111740 70204
rect 111740 70148 111796 70204
rect 111796 70148 111800 70204
rect 111736 70144 111800 70148
rect 111816 70204 111880 70208
rect 111816 70148 111820 70204
rect 111820 70148 111876 70204
rect 111876 70148 111880 70204
rect 111816 70144 111880 70148
rect 111896 70204 111960 70208
rect 111896 70148 111900 70204
rect 111900 70148 111956 70204
rect 111956 70148 111960 70204
rect 111896 70144 111960 70148
rect 111976 70204 112040 70208
rect 111976 70148 111980 70204
rect 111980 70148 112036 70204
rect 112036 70148 112040 70204
rect 111976 70144 112040 70148
rect 142456 70204 142520 70208
rect 142456 70148 142460 70204
rect 142460 70148 142516 70204
rect 142516 70148 142520 70204
rect 142456 70144 142520 70148
rect 142536 70204 142600 70208
rect 142536 70148 142540 70204
rect 142540 70148 142596 70204
rect 142596 70148 142600 70204
rect 142536 70144 142600 70148
rect 142616 70204 142680 70208
rect 142616 70148 142620 70204
rect 142620 70148 142676 70204
rect 142676 70148 142680 70204
rect 142616 70144 142680 70148
rect 142696 70204 142760 70208
rect 142696 70148 142700 70204
rect 142700 70148 142756 70204
rect 142756 70148 142760 70204
rect 142696 70144 142760 70148
rect 173176 70204 173240 70208
rect 173176 70148 173180 70204
rect 173180 70148 173236 70204
rect 173236 70148 173240 70204
rect 173176 70144 173240 70148
rect 173256 70204 173320 70208
rect 173256 70148 173260 70204
rect 173260 70148 173316 70204
rect 173316 70148 173320 70204
rect 173256 70144 173320 70148
rect 173336 70204 173400 70208
rect 173336 70148 173340 70204
rect 173340 70148 173396 70204
rect 173396 70148 173400 70204
rect 173336 70144 173400 70148
rect 173416 70204 173480 70208
rect 173416 70148 173420 70204
rect 173420 70148 173476 70204
rect 173476 70148 173480 70204
rect 173416 70144 173480 70148
rect 4216 69660 4280 69664
rect 4216 69604 4220 69660
rect 4220 69604 4276 69660
rect 4276 69604 4280 69660
rect 4216 69600 4280 69604
rect 4296 69660 4360 69664
rect 4296 69604 4300 69660
rect 4300 69604 4356 69660
rect 4356 69604 4360 69660
rect 4296 69600 4360 69604
rect 4376 69660 4440 69664
rect 4376 69604 4380 69660
rect 4380 69604 4436 69660
rect 4436 69604 4440 69660
rect 4376 69600 4440 69604
rect 4456 69660 4520 69664
rect 4456 69604 4460 69660
rect 4460 69604 4516 69660
rect 4516 69604 4520 69660
rect 4456 69600 4520 69604
rect 34936 69660 35000 69664
rect 34936 69604 34940 69660
rect 34940 69604 34996 69660
rect 34996 69604 35000 69660
rect 34936 69600 35000 69604
rect 35016 69660 35080 69664
rect 35016 69604 35020 69660
rect 35020 69604 35076 69660
rect 35076 69604 35080 69660
rect 35016 69600 35080 69604
rect 35096 69660 35160 69664
rect 35096 69604 35100 69660
rect 35100 69604 35156 69660
rect 35156 69604 35160 69660
rect 35096 69600 35160 69604
rect 35176 69660 35240 69664
rect 35176 69604 35180 69660
rect 35180 69604 35236 69660
rect 35236 69604 35240 69660
rect 35176 69600 35240 69604
rect 65656 69660 65720 69664
rect 65656 69604 65660 69660
rect 65660 69604 65716 69660
rect 65716 69604 65720 69660
rect 65656 69600 65720 69604
rect 65736 69660 65800 69664
rect 65736 69604 65740 69660
rect 65740 69604 65796 69660
rect 65796 69604 65800 69660
rect 65736 69600 65800 69604
rect 65816 69660 65880 69664
rect 65816 69604 65820 69660
rect 65820 69604 65876 69660
rect 65876 69604 65880 69660
rect 65816 69600 65880 69604
rect 65896 69660 65960 69664
rect 65896 69604 65900 69660
rect 65900 69604 65956 69660
rect 65956 69604 65960 69660
rect 65896 69600 65960 69604
rect 96376 69660 96440 69664
rect 96376 69604 96380 69660
rect 96380 69604 96436 69660
rect 96436 69604 96440 69660
rect 96376 69600 96440 69604
rect 96456 69660 96520 69664
rect 96456 69604 96460 69660
rect 96460 69604 96516 69660
rect 96516 69604 96520 69660
rect 96456 69600 96520 69604
rect 96536 69660 96600 69664
rect 96536 69604 96540 69660
rect 96540 69604 96596 69660
rect 96596 69604 96600 69660
rect 96536 69600 96600 69604
rect 96616 69660 96680 69664
rect 96616 69604 96620 69660
rect 96620 69604 96676 69660
rect 96676 69604 96680 69660
rect 96616 69600 96680 69604
rect 127096 69660 127160 69664
rect 127096 69604 127100 69660
rect 127100 69604 127156 69660
rect 127156 69604 127160 69660
rect 127096 69600 127160 69604
rect 127176 69660 127240 69664
rect 127176 69604 127180 69660
rect 127180 69604 127236 69660
rect 127236 69604 127240 69660
rect 127176 69600 127240 69604
rect 127256 69660 127320 69664
rect 127256 69604 127260 69660
rect 127260 69604 127316 69660
rect 127316 69604 127320 69660
rect 127256 69600 127320 69604
rect 127336 69660 127400 69664
rect 127336 69604 127340 69660
rect 127340 69604 127396 69660
rect 127396 69604 127400 69660
rect 127336 69600 127400 69604
rect 157816 69660 157880 69664
rect 157816 69604 157820 69660
rect 157820 69604 157876 69660
rect 157876 69604 157880 69660
rect 157816 69600 157880 69604
rect 157896 69660 157960 69664
rect 157896 69604 157900 69660
rect 157900 69604 157956 69660
rect 157956 69604 157960 69660
rect 157896 69600 157960 69604
rect 157976 69660 158040 69664
rect 157976 69604 157980 69660
rect 157980 69604 158036 69660
rect 158036 69604 158040 69660
rect 157976 69600 158040 69604
rect 158056 69660 158120 69664
rect 158056 69604 158060 69660
rect 158060 69604 158116 69660
rect 158116 69604 158120 69660
rect 158056 69600 158120 69604
rect 19576 69116 19640 69120
rect 19576 69060 19580 69116
rect 19580 69060 19636 69116
rect 19636 69060 19640 69116
rect 19576 69056 19640 69060
rect 19656 69116 19720 69120
rect 19656 69060 19660 69116
rect 19660 69060 19716 69116
rect 19716 69060 19720 69116
rect 19656 69056 19720 69060
rect 19736 69116 19800 69120
rect 19736 69060 19740 69116
rect 19740 69060 19796 69116
rect 19796 69060 19800 69116
rect 19736 69056 19800 69060
rect 19816 69116 19880 69120
rect 19816 69060 19820 69116
rect 19820 69060 19876 69116
rect 19876 69060 19880 69116
rect 19816 69056 19880 69060
rect 50296 69116 50360 69120
rect 50296 69060 50300 69116
rect 50300 69060 50356 69116
rect 50356 69060 50360 69116
rect 50296 69056 50360 69060
rect 50376 69116 50440 69120
rect 50376 69060 50380 69116
rect 50380 69060 50436 69116
rect 50436 69060 50440 69116
rect 50376 69056 50440 69060
rect 50456 69116 50520 69120
rect 50456 69060 50460 69116
rect 50460 69060 50516 69116
rect 50516 69060 50520 69116
rect 50456 69056 50520 69060
rect 50536 69116 50600 69120
rect 50536 69060 50540 69116
rect 50540 69060 50596 69116
rect 50596 69060 50600 69116
rect 50536 69056 50600 69060
rect 81016 69116 81080 69120
rect 81016 69060 81020 69116
rect 81020 69060 81076 69116
rect 81076 69060 81080 69116
rect 81016 69056 81080 69060
rect 81096 69116 81160 69120
rect 81096 69060 81100 69116
rect 81100 69060 81156 69116
rect 81156 69060 81160 69116
rect 81096 69056 81160 69060
rect 81176 69116 81240 69120
rect 81176 69060 81180 69116
rect 81180 69060 81236 69116
rect 81236 69060 81240 69116
rect 81176 69056 81240 69060
rect 81256 69116 81320 69120
rect 81256 69060 81260 69116
rect 81260 69060 81316 69116
rect 81316 69060 81320 69116
rect 81256 69056 81320 69060
rect 111736 69116 111800 69120
rect 111736 69060 111740 69116
rect 111740 69060 111796 69116
rect 111796 69060 111800 69116
rect 111736 69056 111800 69060
rect 111816 69116 111880 69120
rect 111816 69060 111820 69116
rect 111820 69060 111876 69116
rect 111876 69060 111880 69116
rect 111816 69056 111880 69060
rect 111896 69116 111960 69120
rect 111896 69060 111900 69116
rect 111900 69060 111956 69116
rect 111956 69060 111960 69116
rect 111896 69056 111960 69060
rect 111976 69116 112040 69120
rect 111976 69060 111980 69116
rect 111980 69060 112036 69116
rect 112036 69060 112040 69116
rect 111976 69056 112040 69060
rect 142456 69116 142520 69120
rect 142456 69060 142460 69116
rect 142460 69060 142516 69116
rect 142516 69060 142520 69116
rect 142456 69056 142520 69060
rect 142536 69116 142600 69120
rect 142536 69060 142540 69116
rect 142540 69060 142596 69116
rect 142596 69060 142600 69116
rect 142536 69056 142600 69060
rect 142616 69116 142680 69120
rect 142616 69060 142620 69116
rect 142620 69060 142676 69116
rect 142676 69060 142680 69116
rect 142616 69056 142680 69060
rect 142696 69116 142760 69120
rect 142696 69060 142700 69116
rect 142700 69060 142756 69116
rect 142756 69060 142760 69116
rect 142696 69056 142760 69060
rect 173176 69116 173240 69120
rect 173176 69060 173180 69116
rect 173180 69060 173236 69116
rect 173236 69060 173240 69116
rect 173176 69056 173240 69060
rect 173256 69116 173320 69120
rect 173256 69060 173260 69116
rect 173260 69060 173316 69116
rect 173316 69060 173320 69116
rect 173256 69056 173320 69060
rect 173336 69116 173400 69120
rect 173336 69060 173340 69116
rect 173340 69060 173396 69116
rect 173396 69060 173400 69116
rect 173336 69056 173400 69060
rect 173416 69116 173480 69120
rect 173416 69060 173420 69116
rect 173420 69060 173476 69116
rect 173476 69060 173480 69116
rect 173416 69056 173480 69060
rect 4216 68572 4280 68576
rect 4216 68516 4220 68572
rect 4220 68516 4276 68572
rect 4276 68516 4280 68572
rect 4216 68512 4280 68516
rect 4296 68572 4360 68576
rect 4296 68516 4300 68572
rect 4300 68516 4356 68572
rect 4356 68516 4360 68572
rect 4296 68512 4360 68516
rect 4376 68572 4440 68576
rect 4376 68516 4380 68572
rect 4380 68516 4436 68572
rect 4436 68516 4440 68572
rect 4376 68512 4440 68516
rect 4456 68572 4520 68576
rect 4456 68516 4460 68572
rect 4460 68516 4516 68572
rect 4516 68516 4520 68572
rect 4456 68512 4520 68516
rect 34936 68572 35000 68576
rect 34936 68516 34940 68572
rect 34940 68516 34996 68572
rect 34996 68516 35000 68572
rect 34936 68512 35000 68516
rect 35016 68572 35080 68576
rect 35016 68516 35020 68572
rect 35020 68516 35076 68572
rect 35076 68516 35080 68572
rect 35016 68512 35080 68516
rect 35096 68572 35160 68576
rect 35096 68516 35100 68572
rect 35100 68516 35156 68572
rect 35156 68516 35160 68572
rect 35096 68512 35160 68516
rect 35176 68572 35240 68576
rect 35176 68516 35180 68572
rect 35180 68516 35236 68572
rect 35236 68516 35240 68572
rect 35176 68512 35240 68516
rect 65656 68572 65720 68576
rect 65656 68516 65660 68572
rect 65660 68516 65716 68572
rect 65716 68516 65720 68572
rect 65656 68512 65720 68516
rect 65736 68572 65800 68576
rect 65736 68516 65740 68572
rect 65740 68516 65796 68572
rect 65796 68516 65800 68572
rect 65736 68512 65800 68516
rect 65816 68572 65880 68576
rect 65816 68516 65820 68572
rect 65820 68516 65876 68572
rect 65876 68516 65880 68572
rect 65816 68512 65880 68516
rect 65896 68572 65960 68576
rect 65896 68516 65900 68572
rect 65900 68516 65956 68572
rect 65956 68516 65960 68572
rect 65896 68512 65960 68516
rect 96376 68572 96440 68576
rect 96376 68516 96380 68572
rect 96380 68516 96436 68572
rect 96436 68516 96440 68572
rect 96376 68512 96440 68516
rect 96456 68572 96520 68576
rect 96456 68516 96460 68572
rect 96460 68516 96516 68572
rect 96516 68516 96520 68572
rect 96456 68512 96520 68516
rect 96536 68572 96600 68576
rect 96536 68516 96540 68572
rect 96540 68516 96596 68572
rect 96596 68516 96600 68572
rect 96536 68512 96600 68516
rect 96616 68572 96680 68576
rect 96616 68516 96620 68572
rect 96620 68516 96676 68572
rect 96676 68516 96680 68572
rect 96616 68512 96680 68516
rect 127096 68572 127160 68576
rect 127096 68516 127100 68572
rect 127100 68516 127156 68572
rect 127156 68516 127160 68572
rect 127096 68512 127160 68516
rect 127176 68572 127240 68576
rect 127176 68516 127180 68572
rect 127180 68516 127236 68572
rect 127236 68516 127240 68572
rect 127176 68512 127240 68516
rect 127256 68572 127320 68576
rect 127256 68516 127260 68572
rect 127260 68516 127316 68572
rect 127316 68516 127320 68572
rect 127256 68512 127320 68516
rect 127336 68572 127400 68576
rect 127336 68516 127340 68572
rect 127340 68516 127396 68572
rect 127396 68516 127400 68572
rect 127336 68512 127400 68516
rect 157816 68572 157880 68576
rect 157816 68516 157820 68572
rect 157820 68516 157876 68572
rect 157876 68516 157880 68572
rect 157816 68512 157880 68516
rect 157896 68572 157960 68576
rect 157896 68516 157900 68572
rect 157900 68516 157956 68572
rect 157956 68516 157960 68572
rect 157896 68512 157960 68516
rect 157976 68572 158040 68576
rect 157976 68516 157980 68572
rect 157980 68516 158036 68572
rect 158036 68516 158040 68572
rect 157976 68512 158040 68516
rect 158056 68572 158120 68576
rect 158056 68516 158060 68572
rect 158060 68516 158116 68572
rect 158116 68516 158120 68572
rect 158056 68512 158120 68516
rect 19576 68028 19640 68032
rect 19576 67972 19580 68028
rect 19580 67972 19636 68028
rect 19636 67972 19640 68028
rect 19576 67968 19640 67972
rect 19656 68028 19720 68032
rect 19656 67972 19660 68028
rect 19660 67972 19716 68028
rect 19716 67972 19720 68028
rect 19656 67968 19720 67972
rect 19736 68028 19800 68032
rect 19736 67972 19740 68028
rect 19740 67972 19796 68028
rect 19796 67972 19800 68028
rect 19736 67968 19800 67972
rect 19816 68028 19880 68032
rect 19816 67972 19820 68028
rect 19820 67972 19876 68028
rect 19876 67972 19880 68028
rect 19816 67968 19880 67972
rect 50296 68028 50360 68032
rect 50296 67972 50300 68028
rect 50300 67972 50356 68028
rect 50356 67972 50360 68028
rect 50296 67968 50360 67972
rect 50376 68028 50440 68032
rect 50376 67972 50380 68028
rect 50380 67972 50436 68028
rect 50436 67972 50440 68028
rect 50376 67968 50440 67972
rect 50456 68028 50520 68032
rect 50456 67972 50460 68028
rect 50460 67972 50516 68028
rect 50516 67972 50520 68028
rect 50456 67968 50520 67972
rect 50536 68028 50600 68032
rect 50536 67972 50540 68028
rect 50540 67972 50596 68028
rect 50596 67972 50600 68028
rect 50536 67968 50600 67972
rect 81016 68028 81080 68032
rect 81016 67972 81020 68028
rect 81020 67972 81076 68028
rect 81076 67972 81080 68028
rect 81016 67968 81080 67972
rect 81096 68028 81160 68032
rect 81096 67972 81100 68028
rect 81100 67972 81156 68028
rect 81156 67972 81160 68028
rect 81096 67968 81160 67972
rect 81176 68028 81240 68032
rect 81176 67972 81180 68028
rect 81180 67972 81236 68028
rect 81236 67972 81240 68028
rect 81176 67968 81240 67972
rect 81256 68028 81320 68032
rect 81256 67972 81260 68028
rect 81260 67972 81316 68028
rect 81316 67972 81320 68028
rect 81256 67968 81320 67972
rect 111736 68028 111800 68032
rect 111736 67972 111740 68028
rect 111740 67972 111796 68028
rect 111796 67972 111800 68028
rect 111736 67968 111800 67972
rect 111816 68028 111880 68032
rect 111816 67972 111820 68028
rect 111820 67972 111876 68028
rect 111876 67972 111880 68028
rect 111816 67968 111880 67972
rect 111896 68028 111960 68032
rect 111896 67972 111900 68028
rect 111900 67972 111956 68028
rect 111956 67972 111960 68028
rect 111896 67968 111960 67972
rect 111976 68028 112040 68032
rect 111976 67972 111980 68028
rect 111980 67972 112036 68028
rect 112036 67972 112040 68028
rect 111976 67968 112040 67972
rect 142456 68028 142520 68032
rect 142456 67972 142460 68028
rect 142460 67972 142516 68028
rect 142516 67972 142520 68028
rect 142456 67968 142520 67972
rect 142536 68028 142600 68032
rect 142536 67972 142540 68028
rect 142540 67972 142596 68028
rect 142596 67972 142600 68028
rect 142536 67968 142600 67972
rect 142616 68028 142680 68032
rect 142616 67972 142620 68028
rect 142620 67972 142676 68028
rect 142676 67972 142680 68028
rect 142616 67968 142680 67972
rect 142696 68028 142760 68032
rect 142696 67972 142700 68028
rect 142700 67972 142756 68028
rect 142756 67972 142760 68028
rect 142696 67968 142760 67972
rect 173176 68028 173240 68032
rect 173176 67972 173180 68028
rect 173180 67972 173236 68028
rect 173236 67972 173240 68028
rect 173176 67968 173240 67972
rect 173256 68028 173320 68032
rect 173256 67972 173260 68028
rect 173260 67972 173316 68028
rect 173316 67972 173320 68028
rect 173256 67968 173320 67972
rect 173336 68028 173400 68032
rect 173336 67972 173340 68028
rect 173340 67972 173396 68028
rect 173396 67972 173400 68028
rect 173336 67968 173400 67972
rect 173416 68028 173480 68032
rect 173416 67972 173420 68028
rect 173420 67972 173476 68028
rect 173476 67972 173480 68028
rect 173416 67968 173480 67972
rect 4216 67484 4280 67488
rect 4216 67428 4220 67484
rect 4220 67428 4276 67484
rect 4276 67428 4280 67484
rect 4216 67424 4280 67428
rect 4296 67484 4360 67488
rect 4296 67428 4300 67484
rect 4300 67428 4356 67484
rect 4356 67428 4360 67484
rect 4296 67424 4360 67428
rect 4376 67484 4440 67488
rect 4376 67428 4380 67484
rect 4380 67428 4436 67484
rect 4436 67428 4440 67484
rect 4376 67424 4440 67428
rect 4456 67484 4520 67488
rect 4456 67428 4460 67484
rect 4460 67428 4516 67484
rect 4516 67428 4520 67484
rect 4456 67424 4520 67428
rect 34936 67484 35000 67488
rect 34936 67428 34940 67484
rect 34940 67428 34996 67484
rect 34996 67428 35000 67484
rect 34936 67424 35000 67428
rect 35016 67484 35080 67488
rect 35016 67428 35020 67484
rect 35020 67428 35076 67484
rect 35076 67428 35080 67484
rect 35016 67424 35080 67428
rect 35096 67484 35160 67488
rect 35096 67428 35100 67484
rect 35100 67428 35156 67484
rect 35156 67428 35160 67484
rect 35096 67424 35160 67428
rect 35176 67484 35240 67488
rect 35176 67428 35180 67484
rect 35180 67428 35236 67484
rect 35236 67428 35240 67484
rect 35176 67424 35240 67428
rect 65656 67484 65720 67488
rect 65656 67428 65660 67484
rect 65660 67428 65716 67484
rect 65716 67428 65720 67484
rect 65656 67424 65720 67428
rect 65736 67484 65800 67488
rect 65736 67428 65740 67484
rect 65740 67428 65796 67484
rect 65796 67428 65800 67484
rect 65736 67424 65800 67428
rect 65816 67484 65880 67488
rect 65816 67428 65820 67484
rect 65820 67428 65876 67484
rect 65876 67428 65880 67484
rect 65816 67424 65880 67428
rect 65896 67484 65960 67488
rect 65896 67428 65900 67484
rect 65900 67428 65956 67484
rect 65956 67428 65960 67484
rect 65896 67424 65960 67428
rect 96376 67484 96440 67488
rect 96376 67428 96380 67484
rect 96380 67428 96436 67484
rect 96436 67428 96440 67484
rect 96376 67424 96440 67428
rect 96456 67484 96520 67488
rect 96456 67428 96460 67484
rect 96460 67428 96516 67484
rect 96516 67428 96520 67484
rect 96456 67424 96520 67428
rect 96536 67484 96600 67488
rect 96536 67428 96540 67484
rect 96540 67428 96596 67484
rect 96596 67428 96600 67484
rect 96536 67424 96600 67428
rect 96616 67484 96680 67488
rect 96616 67428 96620 67484
rect 96620 67428 96676 67484
rect 96676 67428 96680 67484
rect 96616 67424 96680 67428
rect 127096 67484 127160 67488
rect 127096 67428 127100 67484
rect 127100 67428 127156 67484
rect 127156 67428 127160 67484
rect 127096 67424 127160 67428
rect 127176 67484 127240 67488
rect 127176 67428 127180 67484
rect 127180 67428 127236 67484
rect 127236 67428 127240 67484
rect 127176 67424 127240 67428
rect 127256 67484 127320 67488
rect 127256 67428 127260 67484
rect 127260 67428 127316 67484
rect 127316 67428 127320 67484
rect 127256 67424 127320 67428
rect 127336 67484 127400 67488
rect 127336 67428 127340 67484
rect 127340 67428 127396 67484
rect 127396 67428 127400 67484
rect 127336 67424 127400 67428
rect 157816 67484 157880 67488
rect 157816 67428 157820 67484
rect 157820 67428 157876 67484
rect 157876 67428 157880 67484
rect 157816 67424 157880 67428
rect 157896 67484 157960 67488
rect 157896 67428 157900 67484
rect 157900 67428 157956 67484
rect 157956 67428 157960 67484
rect 157896 67424 157960 67428
rect 157976 67484 158040 67488
rect 157976 67428 157980 67484
rect 157980 67428 158036 67484
rect 158036 67428 158040 67484
rect 157976 67424 158040 67428
rect 158056 67484 158120 67488
rect 158056 67428 158060 67484
rect 158060 67428 158116 67484
rect 158116 67428 158120 67484
rect 158056 67424 158120 67428
rect 19576 66940 19640 66944
rect 19576 66884 19580 66940
rect 19580 66884 19636 66940
rect 19636 66884 19640 66940
rect 19576 66880 19640 66884
rect 19656 66940 19720 66944
rect 19656 66884 19660 66940
rect 19660 66884 19716 66940
rect 19716 66884 19720 66940
rect 19656 66880 19720 66884
rect 19736 66940 19800 66944
rect 19736 66884 19740 66940
rect 19740 66884 19796 66940
rect 19796 66884 19800 66940
rect 19736 66880 19800 66884
rect 19816 66940 19880 66944
rect 19816 66884 19820 66940
rect 19820 66884 19876 66940
rect 19876 66884 19880 66940
rect 19816 66880 19880 66884
rect 50296 66940 50360 66944
rect 50296 66884 50300 66940
rect 50300 66884 50356 66940
rect 50356 66884 50360 66940
rect 50296 66880 50360 66884
rect 50376 66940 50440 66944
rect 50376 66884 50380 66940
rect 50380 66884 50436 66940
rect 50436 66884 50440 66940
rect 50376 66880 50440 66884
rect 50456 66940 50520 66944
rect 50456 66884 50460 66940
rect 50460 66884 50516 66940
rect 50516 66884 50520 66940
rect 50456 66880 50520 66884
rect 50536 66940 50600 66944
rect 50536 66884 50540 66940
rect 50540 66884 50596 66940
rect 50596 66884 50600 66940
rect 50536 66880 50600 66884
rect 81016 66940 81080 66944
rect 81016 66884 81020 66940
rect 81020 66884 81076 66940
rect 81076 66884 81080 66940
rect 81016 66880 81080 66884
rect 81096 66940 81160 66944
rect 81096 66884 81100 66940
rect 81100 66884 81156 66940
rect 81156 66884 81160 66940
rect 81096 66880 81160 66884
rect 81176 66940 81240 66944
rect 81176 66884 81180 66940
rect 81180 66884 81236 66940
rect 81236 66884 81240 66940
rect 81176 66880 81240 66884
rect 81256 66940 81320 66944
rect 81256 66884 81260 66940
rect 81260 66884 81316 66940
rect 81316 66884 81320 66940
rect 81256 66880 81320 66884
rect 111736 66940 111800 66944
rect 111736 66884 111740 66940
rect 111740 66884 111796 66940
rect 111796 66884 111800 66940
rect 111736 66880 111800 66884
rect 111816 66940 111880 66944
rect 111816 66884 111820 66940
rect 111820 66884 111876 66940
rect 111876 66884 111880 66940
rect 111816 66880 111880 66884
rect 111896 66940 111960 66944
rect 111896 66884 111900 66940
rect 111900 66884 111956 66940
rect 111956 66884 111960 66940
rect 111896 66880 111960 66884
rect 111976 66940 112040 66944
rect 111976 66884 111980 66940
rect 111980 66884 112036 66940
rect 112036 66884 112040 66940
rect 111976 66880 112040 66884
rect 142456 66940 142520 66944
rect 142456 66884 142460 66940
rect 142460 66884 142516 66940
rect 142516 66884 142520 66940
rect 142456 66880 142520 66884
rect 142536 66940 142600 66944
rect 142536 66884 142540 66940
rect 142540 66884 142596 66940
rect 142596 66884 142600 66940
rect 142536 66880 142600 66884
rect 142616 66940 142680 66944
rect 142616 66884 142620 66940
rect 142620 66884 142676 66940
rect 142676 66884 142680 66940
rect 142616 66880 142680 66884
rect 142696 66940 142760 66944
rect 142696 66884 142700 66940
rect 142700 66884 142756 66940
rect 142756 66884 142760 66940
rect 142696 66880 142760 66884
rect 173176 66940 173240 66944
rect 173176 66884 173180 66940
rect 173180 66884 173236 66940
rect 173236 66884 173240 66940
rect 173176 66880 173240 66884
rect 173256 66940 173320 66944
rect 173256 66884 173260 66940
rect 173260 66884 173316 66940
rect 173316 66884 173320 66940
rect 173256 66880 173320 66884
rect 173336 66940 173400 66944
rect 173336 66884 173340 66940
rect 173340 66884 173396 66940
rect 173396 66884 173400 66940
rect 173336 66880 173400 66884
rect 173416 66940 173480 66944
rect 173416 66884 173420 66940
rect 173420 66884 173476 66940
rect 173476 66884 173480 66940
rect 173416 66880 173480 66884
rect 4216 66396 4280 66400
rect 4216 66340 4220 66396
rect 4220 66340 4276 66396
rect 4276 66340 4280 66396
rect 4216 66336 4280 66340
rect 4296 66396 4360 66400
rect 4296 66340 4300 66396
rect 4300 66340 4356 66396
rect 4356 66340 4360 66396
rect 4296 66336 4360 66340
rect 4376 66396 4440 66400
rect 4376 66340 4380 66396
rect 4380 66340 4436 66396
rect 4436 66340 4440 66396
rect 4376 66336 4440 66340
rect 4456 66396 4520 66400
rect 4456 66340 4460 66396
rect 4460 66340 4516 66396
rect 4516 66340 4520 66396
rect 4456 66336 4520 66340
rect 34936 66396 35000 66400
rect 34936 66340 34940 66396
rect 34940 66340 34996 66396
rect 34996 66340 35000 66396
rect 34936 66336 35000 66340
rect 35016 66396 35080 66400
rect 35016 66340 35020 66396
rect 35020 66340 35076 66396
rect 35076 66340 35080 66396
rect 35016 66336 35080 66340
rect 35096 66396 35160 66400
rect 35096 66340 35100 66396
rect 35100 66340 35156 66396
rect 35156 66340 35160 66396
rect 35096 66336 35160 66340
rect 35176 66396 35240 66400
rect 35176 66340 35180 66396
rect 35180 66340 35236 66396
rect 35236 66340 35240 66396
rect 35176 66336 35240 66340
rect 65656 66396 65720 66400
rect 65656 66340 65660 66396
rect 65660 66340 65716 66396
rect 65716 66340 65720 66396
rect 65656 66336 65720 66340
rect 65736 66396 65800 66400
rect 65736 66340 65740 66396
rect 65740 66340 65796 66396
rect 65796 66340 65800 66396
rect 65736 66336 65800 66340
rect 65816 66396 65880 66400
rect 65816 66340 65820 66396
rect 65820 66340 65876 66396
rect 65876 66340 65880 66396
rect 65816 66336 65880 66340
rect 65896 66396 65960 66400
rect 65896 66340 65900 66396
rect 65900 66340 65956 66396
rect 65956 66340 65960 66396
rect 65896 66336 65960 66340
rect 96376 66396 96440 66400
rect 96376 66340 96380 66396
rect 96380 66340 96436 66396
rect 96436 66340 96440 66396
rect 96376 66336 96440 66340
rect 96456 66396 96520 66400
rect 96456 66340 96460 66396
rect 96460 66340 96516 66396
rect 96516 66340 96520 66396
rect 96456 66336 96520 66340
rect 96536 66396 96600 66400
rect 96536 66340 96540 66396
rect 96540 66340 96596 66396
rect 96596 66340 96600 66396
rect 96536 66336 96600 66340
rect 96616 66396 96680 66400
rect 96616 66340 96620 66396
rect 96620 66340 96676 66396
rect 96676 66340 96680 66396
rect 96616 66336 96680 66340
rect 127096 66396 127160 66400
rect 127096 66340 127100 66396
rect 127100 66340 127156 66396
rect 127156 66340 127160 66396
rect 127096 66336 127160 66340
rect 127176 66396 127240 66400
rect 127176 66340 127180 66396
rect 127180 66340 127236 66396
rect 127236 66340 127240 66396
rect 127176 66336 127240 66340
rect 127256 66396 127320 66400
rect 127256 66340 127260 66396
rect 127260 66340 127316 66396
rect 127316 66340 127320 66396
rect 127256 66336 127320 66340
rect 127336 66396 127400 66400
rect 127336 66340 127340 66396
rect 127340 66340 127396 66396
rect 127396 66340 127400 66396
rect 127336 66336 127400 66340
rect 157816 66396 157880 66400
rect 157816 66340 157820 66396
rect 157820 66340 157876 66396
rect 157876 66340 157880 66396
rect 157816 66336 157880 66340
rect 157896 66396 157960 66400
rect 157896 66340 157900 66396
rect 157900 66340 157956 66396
rect 157956 66340 157960 66396
rect 157896 66336 157960 66340
rect 157976 66396 158040 66400
rect 157976 66340 157980 66396
rect 157980 66340 158036 66396
rect 158036 66340 158040 66396
rect 157976 66336 158040 66340
rect 158056 66396 158120 66400
rect 158056 66340 158060 66396
rect 158060 66340 158116 66396
rect 158116 66340 158120 66396
rect 158056 66336 158120 66340
rect 19576 65852 19640 65856
rect 19576 65796 19580 65852
rect 19580 65796 19636 65852
rect 19636 65796 19640 65852
rect 19576 65792 19640 65796
rect 19656 65852 19720 65856
rect 19656 65796 19660 65852
rect 19660 65796 19716 65852
rect 19716 65796 19720 65852
rect 19656 65792 19720 65796
rect 19736 65852 19800 65856
rect 19736 65796 19740 65852
rect 19740 65796 19796 65852
rect 19796 65796 19800 65852
rect 19736 65792 19800 65796
rect 19816 65852 19880 65856
rect 19816 65796 19820 65852
rect 19820 65796 19876 65852
rect 19876 65796 19880 65852
rect 19816 65792 19880 65796
rect 50296 65852 50360 65856
rect 50296 65796 50300 65852
rect 50300 65796 50356 65852
rect 50356 65796 50360 65852
rect 50296 65792 50360 65796
rect 50376 65852 50440 65856
rect 50376 65796 50380 65852
rect 50380 65796 50436 65852
rect 50436 65796 50440 65852
rect 50376 65792 50440 65796
rect 50456 65852 50520 65856
rect 50456 65796 50460 65852
rect 50460 65796 50516 65852
rect 50516 65796 50520 65852
rect 50456 65792 50520 65796
rect 50536 65852 50600 65856
rect 50536 65796 50540 65852
rect 50540 65796 50596 65852
rect 50596 65796 50600 65852
rect 50536 65792 50600 65796
rect 81016 65852 81080 65856
rect 81016 65796 81020 65852
rect 81020 65796 81076 65852
rect 81076 65796 81080 65852
rect 81016 65792 81080 65796
rect 81096 65852 81160 65856
rect 81096 65796 81100 65852
rect 81100 65796 81156 65852
rect 81156 65796 81160 65852
rect 81096 65792 81160 65796
rect 81176 65852 81240 65856
rect 81176 65796 81180 65852
rect 81180 65796 81236 65852
rect 81236 65796 81240 65852
rect 81176 65792 81240 65796
rect 81256 65852 81320 65856
rect 81256 65796 81260 65852
rect 81260 65796 81316 65852
rect 81316 65796 81320 65852
rect 81256 65792 81320 65796
rect 111736 65852 111800 65856
rect 111736 65796 111740 65852
rect 111740 65796 111796 65852
rect 111796 65796 111800 65852
rect 111736 65792 111800 65796
rect 111816 65852 111880 65856
rect 111816 65796 111820 65852
rect 111820 65796 111876 65852
rect 111876 65796 111880 65852
rect 111816 65792 111880 65796
rect 111896 65852 111960 65856
rect 111896 65796 111900 65852
rect 111900 65796 111956 65852
rect 111956 65796 111960 65852
rect 111896 65792 111960 65796
rect 111976 65852 112040 65856
rect 111976 65796 111980 65852
rect 111980 65796 112036 65852
rect 112036 65796 112040 65852
rect 111976 65792 112040 65796
rect 142456 65852 142520 65856
rect 142456 65796 142460 65852
rect 142460 65796 142516 65852
rect 142516 65796 142520 65852
rect 142456 65792 142520 65796
rect 142536 65852 142600 65856
rect 142536 65796 142540 65852
rect 142540 65796 142596 65852
rect 142596 65796 142600 65852
rect 142536 65792 142600 65796
rect 142616 65852 142680 65856
rect 142616 65796 142620 65852
rect 142620 65796 142676 65852
rect 142676 65796 142680 65852
rect 142616 65792 142680 65796
rect 142696 65852 142760 65856
rect 142696 65796 142700 65852
rect 142700 65796 142756 65852
rect 142756 65796 142760 65852
rect 142696 65792 142760 65796
rect 173176 65852 173240 65856
rect 173176 65796 173180 65852
rect 173180 65796 173236 65852
rect 173236 65796 173240 65852
rect 173176 65792 173240 65796
rect 173256 65852 173320 65856
rect 173256 65796 173260 65852
rect 173260 65796 173316 65852
rect 173316 65796 173320 65852
rect 173256 65792 173320 65796
rect 173336 65852 173400 65856
rect 173336 65796 173340 65852
rect 173340 65796 173396 65852
rect 173396 65796 173400 65852
rect 173336 65792 173400 65796
rect 173416 65852 173480 65856
rect 173416 65796 173420 65852
rect 173420 65796 173476 65852
rect 173476 65796 173480 65852
rect 173416 65792 173480 65796
rect 4216 65308 4280 65312
rect 4216 65252 4220 65308
rect 4220 65252 4276 65308
rect 4276 65252 4280 65308
rect 4216 65248 4280 65252
rect 4296 65308 4360 65312
rect 4296 65252 4300 65308
rect 4300 65252 4356 65308
rect 4356 65252 4360 65308
rect 4296 65248 4360 65252
rect 4376 65308 4440 65312
rect 4376 65252 4380 65308
rect 4380 65252 4436 65308
rect 4436 65252 4440 65308
rect 4376 65248 4440 65252
rect 4456 65308 4520 65312
rect 4456 65252 4460 65308
rect 4460 65252 4516 65308
rect 4516 65252 4520 65308
rect 4456 65248 4520 65252
rect 34936 65308 35000 65312
rect 34936 65252 34940 65308
rect 34940 65252 34996 65308
rect 34996 65252 35000 65308
rect 34936 65248 35000 65252
rect 35016 65308 35080 65312
rect 35016 65252 35020 65308
rect 35020 65252 35076 65308
rect 35076 65252 35080 65308
rect 35016 65248 35080 65252
rect 35096 65308 35160 65312
rect 35096 65252 35100 65308
rect 35100 65252 35156 65308
rect 35156 65252 35160 65308
rect 35096 65248 35160 65252
rect 35176 65308 35240 65312
rect 35176 65252 35180 65308
rect 35180 65252 35236 65308
rect 35236 65252 35240 65308
rect 35176 65248 35240 65252
rect 65656 65308 65720 65312
rect 65656 65252 65660 65308
rect 65660 65252 65716 65308
rect 65716 65252 65720 65308
rect 65656 65248 65720 65252
rect 65736 65308 65800 65312
rect 65736 65252 65740 65308
rect 65740 65252 65796 65308
rect 65796 65252 65800 65308
rect 65736 65248 65800 65252
rect 65816 65308 65880 65312
rect 65816 65252 65820 65308
rect 65820 65252 65876 65308
rect 65876 65252 65880 65308
rect 65816 65248 65880 65252
rect 65896 65308 65960 65312
rect 65896 65252 65900 65308
rect 65900 65252 65956 65308
rect 65956 65252 65960 65308
rect 65896 65248 65960 65252
rect 96376 65308 96440 65312
rect 96376 65252 96380 65308
rect 96380 65252 96436 65308
rect 96436 65252 96440 65308
rect 96376 65248 96440 65252
rect 96456 65308 96520 65312
rect 96456 65252 96460 65308
rect 96460 65252 96516 65308
rect 96516 65252 96520 65308
rect 96456 65248 96520 65252
rect 96536 65308 96600 65312
rect 96536 65252 96540 65308
rect 96540 65252 96596 65308
rect 96596 65252 96600 65308
rect 96536 65248 96600 65252
rect 96616 65308 96680 65312
rect 96616 65252 96620 65308
rect 96620 65252 96676 65308
rect 96676 65252 96680 65308
rect 96616 65248 96680 65252
rect 127096 65308 127160 65312
rect 127096 65252 127100 65308
rect 127100 65252 127156 65308
rect 127156 65252 127160 65308
rect 127096 65248 127160 65252
rect 127176 65308 127240 65312
rect 127176 65252 127180 65308
rect 127180 65252 127236 65308
rect 127236 65252 127240 65308
rect 127176 65248 127240 65252
rect 127256 65308 127320 65312
rect 127256 65252 127260 65308
rect 127260 65252 127316 65308
rect 127316 65252 127320 65308
rect 127256 65248 127320 65252
rect 127336 65308 127400 65312
rect 127336 65252 127340 65308
rect 127340 65252 127396 65308
rect 127396 65252 127400 65308
rect 127336 65248 127400 65252
rect 157816 65308 157880 65312
rect 157816 65252 157820 65308
rect 157820 65252 157876 65308
rect 157876 65252 157880 65308
rect 157816 65248 157880 65252
rect 157896 65308 157960 65312
rect 157896 65252 157900 65308
rect 157900 65252 157956 65308
rect 157956 65252 157960 65308
rect 157896 65248 157960 65252
rect 157976 65308 158040 65312
rect 157976 65252 157980 65308
rect 157980 65252 158036 65308
rect 158036 65252 158040 65308
rect 157976 65248 158040 65252
rect 158056 65308 158120 65312
rect 158056 65252 158060 65308
rect 158060 65252 158116 65308
rect 158116 65252 158120 65308
rect 158056 65248 158120 65252
rect 19576 64764 19640 64768
rect 19576 64708 19580 64764
rect 19580 64708 19636 64764
rect 19636 64708 19640 64764
rect 19576 64704 19640 64708
rect 19656 64764 19720 64768
rect 19656 64708 19660 64764
rect 19660 64708 19716 64764
rect 19716 64708 19720 64764
rect 19656 64704 19720 64708
rect 19736 64764 19800 64768
rect 19736 64708 19740 64764
rect 19740 64708 19796 64764
rect 19796 64708 19800 64764
rect 19736 64704 19800 64708
rect 19816 64764 19880 64768
rect 19816 64708 19820 64764
rect 19820 64708 19876 64764
rect 19876 64708 19880 64764
rect 19816 64704 19880 64708
rect 50296 64764 50360 64768
rect 50296 64708 50300 64764
rect 50300 64708 50356 64764
rect 50356 64708 50360 64764
rect 50296 64704 50360 64708
rect 50376 64764 50440 64768
rect 50376 64708 50380 64764
rect 50380 64708 50436 64764
rect 50436 64708 50440 64764
rect 50376 64704 50440 64708
rect 50456 64764 50520 64768
rect 50456 64708 50460 64764
rect 50460 64708 50516 64764
rect 50516 64708 50520 64764
rect 50456 64704 50520 64708
rect 50536 64764 50600 64768
rect 50536 64708 50540 64764
rect 50540 64708 50596 64764
rect 50596 64708 50600 64764
rect 50536 64704 50600 64708
rect 81016 64764 81080 64768
rect 81016 64708 81020 64764
rect 81020 64708 81076 64764
rect 81076 64708 81080 64764
rect 81016 64704 81080 64708
rect 81096 64764 81160 64768
rect 81096 64708 81100 64764
rect 81100 64708 81156 64764
rect 81156 64708 81160 64764
rect 81096 64704 81160 64708
rect 81176 64764 81240 64768
rect 81176 64708 81180 64764
rect 81180 64708 81236 64764
rect 81236 64708 81240 64764
rect 81176 64704 81240 64708
rect 81256 64764 81320 64768
rect 81256 64708 81260 64764
rect 81260 64708 81316 64764
rect 81316 64708 81320 64764
rect 81256 64704 81320 64708
rect 111736 64764 111800 64768
rect 111736 64708 111740 64764
rect 111740 64708 111796 64764
rect 111796 64708 111800 64764
rect 111736 64704 111800 64708
rect 111816 64764 111880 64768
rect 111816 64708 111820 64764
rect 111820 64708 111876 64764
rect 111876 64708 111880 64764
rect 111816 64704 111880 64708
rect 111896 64764 111960 64768
rect 111896 64708 111900 64764
rect 111900 64708 111956 64764
rect 111956 64708 111960 64764
rect 111896 64704 111960 64708
rect 111976 64764 112040 64768
rect 111976 64708 111980 64764
rect 111980 64708 112036 64764
rect 112036 64708 112040 64764
rect 111976 64704 112040 64708
rect 142456 64764 142520 64768
rect 142456 64708 142460 64764
rect 142460 64708 142516 64764
rect 142516 64708 142520 64764
rect 142456 64704 142520 64708
rect 142536 64764 142600 64768
rect 142536 64708 142540 64764
rect 142540 64708 142596 64764
rect 142596 64708 142600 64764
rect 142536 64704 142600 64708
rect 142616 64764 142680 64768
rect 142616 64708 142620 64764
rect 142620 64708 142676 64764
rect 142676 64708 142680 64764
rect 142616 64704 142680 64708
rect 142696 64764 142760 64768
rect 142696 64708 142700 64764
rect 142700 64708 142756 64764
rect 142756 64708 142760 64764
rect 142696 64704 142760 64708
rect 173176 64764 173240 64768
rect 173176 64708 173180 64764
rect 173180 64708 173236 64764
rect 173236 64708 173240 64764
rect 173176 64704 173240 64708
rect 173256 64764 173320 64768
rect 173256 64708 173260 64764
rect 173260 64708 173316 64764
rect 173316 64708 173320 64764
rect 173256 64704 173320 64708
rect 173336 64764 173400 64768
rect 173336 64708 173340 64764
rect 173340 64708 173396 64764
rect 173396 64708 173400 64764
rect 173336 64704 173400 64708
rect 173416 64764 173480 64768
rect 173416 64708 173420 64764
rect 173420 64708 173476 64764
rect 173476 64708 173480 64764
rect 173416 64704 173480 64708
rect 4216 64220 4280 64224
rect 4216 64164 4220 64220
rect 4220 64164 4276 64220
rect 4276 64164 4280 64220
rect 4216 64160 4280 64164
rect 4296 64220 4360 64224
rect 4296 64164 4300 64220
rect 4300 64164 4356 64220
rect 4356 64164 4360 64220
rect 4296 64160 4360 64164
rect 4376 64220 4440 64224
rect 4376 64164 4380 64220
rect 4380 64164 4436 64220
rect 4436 64164 4440 64220
rect 4376 64160 4440 64164
rect 4456 64220 4520 64224
rect 4456 64164 4460 64220
rect 4460 64164 4516 64220
rect 4516 64164 4520 64220
rect 4456 64160 4520 64164
rect 34936 64220 35000 64224
rect 34936 64164 34940 64220
rect 34940 64164 34996 64220
rect 34996 64164 35000 64220
rect 34936 64160 35000 64164
rect 35016 64220 35080 64224
rect 35016 64164 35020 64220
rect 35020 64164 35076 64220
rect 35076 64164 35080 64220
rect 35016 64160 35080 64164
rect 35096 64220 35160 64224
rect 35096 64164 35100 64220
rect 35100 64164 35156 64220
rect 35156 64164 35160 64220
rect 35096 64160 35160 64164
rect 35176 64220 35240 64224
rect 35176 64164 35180 64220
rect 35180 64164 35236 64220
rect 35236 64164 35240 64220
rect 35176 64160 35240 64164
rect 65656 64220 65720 64224
rect 65656 64164 65660 64220
rect 65660 64164 65716 64220
rect 65716 64164 65720 64220
rect 65656 64160 65720 64164
rect 65736 64220 65800 64224
rect 65736 64164 65740 64220
rect 65740 64164 65796 64220
rect 65796 64164 65800 64220
rect 65736 64160 65800 64164
rect 65816 64220 65880 64224
rect 65816 64164 65820 64220
rect 65820 64164 65876 64220
rect 65876 64164 65880 64220
rect 65816 64160 65880 64164
rect 65896 64220 65960 64224
rect 65896 64164 65900 64220
rect 65900 64164 65956 64220
rect 65956 64164 65960 64220
rect 65896 64160 65960 64164
rect 96376 64220 96440 64224
rect 96376 64164 96380 64220
rect 96380 64164 96436 64220
rect 96436 64164 96440 64220
rect 96376 64160 96440 64164
rect 96456 64220 96520 64224
rect 96456 64164 96460 64220
rect 96460 64164 96516 64220
rect 96516 64164 96520 64220
rect 96456 64160 96520 64164
rect 96536 64220 96600 64224
rect 96536 64164 96540 64220
rect 96540 64164 96596 64220
rect 96596 64164 96600 64220
rect 96536 64160 96600 64164
rect 96616 64220 96680 64224
rect 96616 64164 96620 64220
rect 96620 64164 96676 64220
rect 96676 64164 96680 64220
rect 96616 64160 96680 64164
rect 127096 64220 127160 64224
rect 127096 64164 127100 64220
rect 127100 64164 127156 64220
rect 127156 64164 127160 64220
rect 127096 64160 127160 64164
rect 127176 64220 127240 64224
rect 127176 64164 127180 64220
rect 127180 64164 127236 64220
rect 127236 64164 127240 64220
rect 127176 64160 127240 64164
rect 127256 64220 127320 64224
rect 127256 64164 127260 64220
rect 127260 64164 127316 64220
rect 127316 64164 127320 64220
rect 127256 64160 127320 64164
rect 127336 64220 127400 64224
rect 127336 64164 127340 64220
rect 127340 64164 127396 64220
rect 127396 64164 127400 64220
rect 127336 64160 127400 64164
rect 157816 64220 157880 64224
rect 157816 64164 157820 64220
rect 157820 64164 157876 64220
rect 157876 64164 157880 64220
rect 157816 64160 157880 64164
rect 157896 64220 157960 64224
rect 157896 64164 157900 64220
rect 157900 64164 157956 64220
rect 157956 64164 157960 64220
rect 157896 64160 157960 64164
rect 157976 64220 158040 64224
rect 157976 64164 157980 64220
rect 157980 64164 158036 64220
rect 158036 64164 158040 64220
rect 157976 64160 158040 64164
rect 158056 64220 158120 64224
rect 158056 64164 158060 64220
rect 158060 64164 158116 64220
rect 158116 64164 158120 64220
rect 158056 64160 158120 64164
rect 19576 63676 19640 63680
rect 19576 63620 19580 63676
rect 19580 63620 19636 63676
rect 19636 63620 19640 63676
rect 19576 63616 19640 63620
rect 19656 63676 19720 63680
rect 19656 63620 19660 63676
rect 19660 63620 19716 63676
rect 19716 63620 19720 63676
rect 19656 63616 19720 63620
rect 19736 63676 19800 63680
rect 19736 63620 19740 63676
rect 19740 63620 19796 63676
rect 19796 63620 19800 63676
rect 19736 63616 19800 63620
rect 19816 63676 19880 63680
rect 19816 63620 19820 63676
rect 19820 63620 19876 63676
rect 19876 63620 19880 63676
rect 19816 63616 19880 63620
rect 50296 63676 50360 63680
rect 50296 63620 50300 63676
rect 50300 63620 50356 63676
rect 50356 63620 50360 63676
rect 50296 63616 50360 63620
rect 50376 63676 50440 63680
rect 50376 63620 50380 63676
rect 50380 63620 50436 63676
rect 50436 63620 50440 63676
rect 50376 63616 50440 63620
rect 50456 63676 50520 63680
rect 50456 63620 50460 63676
rect 50460 63620 50516 63676
rect 50516 63620 50520 63676
rect 50456 63616 50520 63620
rect 50536 63676 50600 63680
rect 50536 63620 50540 63676
rect 50540 63620 50596 63676
rect 50596 63620 50600 63676
rect 50536 63616 50600 63620
rect 81016 63676 81080 63680
rect 81016 63620 81020 63676
rect 81020 63620 81076 63676
rect 81076 63620 81080 63676
rect 81016 63616 81080 63620
rect 81096 63676 81160 63680
rect 81096 63620 81100 63676
rect 81100 63620 81156 63676
rect 81156 63620 81160 63676
rect 81096 63616 81160 63620
rect 81176 63676 81240 63680
rect 81176 63620 81180 63676
rect 81180 63620 81236 63676
rect 81236 63620 81240 63676
rect 81176 63616 81240 63620
rect 81256 63676 81320 63680
rect 81256 63620 81260 63676
rect 81260 63620 81316 63676
rect 81316 63620 81320 63676
rect 81256 63616 81320 63620
rect 111736 63676 111800 63680
rect 111736 63620 111740 63676
rect 111740 63620 111796 63676
rect 111796 63620 111800 63676
rect 111736 63616 111800 63620
rect 111816 63676 111880 63680
rect 111816 63620 111820 63676
rect 111820 63620 111876 63676
rect 111876 63620 111880 63676
rect 111816 63616 111880 63620
rect 111896 63676 111960 63680
rect 111896 63620 111900 63676
rect 111900 63620 111956 63676
rect 111956 63620 111960 63676
rect 111896 63616 111960 63620
rect 111976 63676 112040 63680
rect 111976 63620 111980 63676
rect 111980 63620 112036 63676
rect 112036 63620 112040 63676
rect 111976 63616 112040 63620
rect 142456 63676 142520 63680
rect 142456 63620 142460 63676
rect 142460 63620 142516 63676
rect 142516 63620 142520 63676
rect 142456 63616 142520 63620
rect 142536 63676 142600 63680
rect 142536 63620 142540 63676
rect 142540 63620 142596 63676
rect 142596 63620 142600 63676
rect 142536 63616 142600 63620
rect 142616 63676 142680 63680
rect 142616 63620 142620 63676
rect 142620 63620 142676 63676
rect 142676 63620 142680 63676
rect 142616 63616 142680 63620
rect 142696 63676 142760 63680
rect 142696 63620 142700 63676
rect 142700 63620 142756 63676
rect 142756 63620 142760 63676
rect 142696 63616 142760 63620
rect 173176 63676 173240 63680
rect 173176 63620 173180 63676
rect 173180 63620 173236 63676
rect 173236 63620 173240 63676
rect 173176 63616 173240 63620
rect 173256 63676 173320 63680
rect 173256 63620 173260 63676
rect 173260 63620 173316 63676
rect 173316 63620 173320 63676
rect 173256 63616 173320 63620
rect 173336 63676 173400 63680
rect 173336 63620 173340 63676
rect 173340 63620 173396 63676
rect 173396 63620 173400 63676
rect 173336 63616 173400 63620
rect 173416 63676 173480 63680
rect 173416 63620 173420 63676
rect 173420 63620 173476 63676
rect 173476 63620 173480 63676
rect 173416 63616 173480 63620
rect 4216 63132 4280 63136
rect 4216 63076 4220 63132
rect 4220 63076 4276 63132
rect 4276 63076 4280 63132
rect 4216 63072 4280 63076
rect 4296 63132 4360 63136
rect 4296 63076 4300 63132
rect 4300 63076 4356 63132
rect 4356 63076 4360 63132
rect 4296 63072 4360 63076
rect 4376 63132 4440 63136
rect 4376 63076 4380 63132
rect 4380 63076 4436 63132
rect 4436 63076 4440 63132
rect 4376 63072 4440 63076
rect 4456 63132 4520 63136
rect 4456 63076 4460 63132
rect 4460 63076 4516 63132
rect 4516 63076 4520 63132
rect 4456 63072 4520 63076
rect 34936 63132 35000 63136
rect 34936 63076 34940 63132
rect 34940 63076 34996 63132
rect 34996 63076 35000 63132
rect 34936 63072 35000 63076
rect 35016 63132 35080 63136
rect 35016 63076 35020 63132
rect 35020 63076 35076 63132
rect 35076 63076 35080 63132
rect 35016 63072 35080 63076
rect 35096 63132 35160 63136
rect 35096 63076 35100 63132
rect 35100 63076 35156 63132
rect 35156 63076 35160 63132
rect 35096 63072 35160 63076
rect 35176 63132 35240 63136
rect 35176 63076 35180 63132
rect 35180 63076 35236 63132
rect 35236 63076 35240 63132
rect 35176 63072 35240 63076
rect 65656 63132 65720 63136
rect 65656 63076 65660 63132
rect 65660 63076 65716 63132
rect 65716 63076 65720 63132
rect 65656 63072 65720 63076
rect 65736 63132 65800 63136
rect 65736 63076 65740 63132
rect 65740 63076 65796 63132
rect 65796 63076 65800 63132
rect 65736 63072 65800 63076
rect 65816 63132 65880 63136
rect 65816 63076 65820 63132
rect 65820 63076 65876 63132
rect 65876 63076 65880 63132
rect 65816 63072 65880 63076
rect 65896 63132 65960 63136
rect 65896 63076 65900 63132
rect 65900 63076 65956 63132
rect 65956 63076 65960 63132
rect 65896 63072 65960 63076
rect 96376 63132 96440 63136
rect 96376 63076 96380 63132
rect 96380 63076 96436 63132
rect 96436 63076 96440 63132
rect 96376 63072 96440 63076
rect 96456 63132 96520 63136
rect 96456 63076 96460 63132
rect 96460 63076 96516 63132
rect 96516 63076 96520 63132
rect 96456 63072 96520 63076
rect 96536 63132 96600 63136
rect 96536 63076 96540 63132
rect 96540 63076 96596 63132
rect 96596 63076 96600 63132
rect 96536 63072 96600 63076
rect 96616 63132 96680 63136
rect 96616 63076 96620 63132
rect 96620 63076 96676 63132
rect 96676 63076 96680 63132
rect 96616 63072 96680 63076
rect 127096 63132 127160 63136
rect 127096 63076 127100 63132
rect 127100 63076 127156 63132
rect 127156 63076 127160 63132
rect 127096 63072 127160 63076
rect 127176 63132 127240 63136
rect 127176 63076 127180 63132
rect 127180 63076 127236 63132
rect 127236 63076 127240 63132
rect 127176 63072 127240 63076
rect 127256 63132 127320 63136
rect 127256 63076 127260 63132
rect 127260 63076 127316 63132
rect 127316 63076 127320 63132
rect 127256 63072 127320 63076
rect 127336 63132 127400 63136
rect 127336 63076 127340 63132
rect 127340 63076 127396 63132
rect 127396 63076 127400 63132
rect 127336 63072 127400 63076
rect 157816 63132 157880 63136
rect 157816 63076 157820 63132
rect 157820 63076 157876 63132
rect 157876 63076 157880 63132
rect 157816 63072 157880 63076
rect 157896 63132 157960 63136
rect 157896 63076 157900 63132
rect 157900 63076 157956 63132
rect 157956 63076 157960 63132
rect 157896 63072 157960 63076
rect 157976 63132 158040 63136
rect 157976 63076 157980 63132
rect 157980 63076 158036 63132
rect 158036 63076 158040 63132
rect 157976 63072 158040 63076
rect 158056 63132 158120 63136
rect 158056 63076 158060 63132
rect 158060 63076 158116 63132
rect 158116 63076 158120 63132
rect 158056 63072 158120 63076
rect 19576 62588 19640 62592
rect 19576 62532 19580 62588
rect 19580 62532 19636 62588
rect 19636 62532 19640 62588
rect 19576 62528 19640 62532
rect 19656 62588 19720 62592
rect 19656 62532 19660 62588
rect 19660 62532 19716 62588
rect 19716 62532 19720 62588
rect 19656 62528 19720 62532
rect 19736 62588 19800 62592
rect 19736 62532 19740 62588
rect 19740 62532 19796 62588
rect 19796 62532 19800 62588
rect 19736 62528 19800 62532
rect 19816 62588 19880 62592
rect 19816 62532 19820 62588
rect 19820 62532 19876 62588
rect 19876 62532 19880 62588
rect 19816 62528 19880 62532
rect 50296 62588 50360 62592
rect 50296 62532 50300 62588
rect 50300 62532 50356 62588
rect 50356 62532 50360 62588
rect 50296 62528 50360 62532
rect 50376 62588 50440 62592
rect 50376 62532 50380 62588
rect 50380 62532 50436 62588
rect 50436 62532 50440 62588
rect 50376 62528 50440 62532
rect 50456 62588 50520 62592
rect 50456 62532 50460 62588
rect 50460 62532 50516 62588
rect 50516 62532 50520 62588
rect 50456 62528 50520 62532
rect 50536 62588 50600 62592
rect 50536 62532 50540 62588
rect 50540 62532 50596 62588
rect 50596 62532 50600 62588
rect 50536 62528 50600 62532
rect 81016 62588 81080 62592
rect 81016 62532 81020 62588
rect 81020 62532 81076 62588
rect 81076 62532 81080 62588
rect 81016 62528 81080 62532
rect 81096 62588 81160 62592
rect 81096 62532 81100 62588
rect 81100 62532 81156 62588
rect 81156 62532 81160 62588
rect 81096 62528 81160 62532
rect 81176 62588 81240 62592
rect 81176 62532 81180 62588
rect 81180 62532 81236 62588
rect 81236 62532 81240 62588
rect 81176 62528 81240 62532
rect 81256 62588 81320 62592
rect 81256 62532 81260 62588
rect 81260 62532 81316 62588
rect 81316 62532 81320 62588
rect 81256 62528 81320 62532
rect 111736 62588 111800 62592
rect 111736 62532 111740 62588
rect 111740 62532 111796 62588
rect 111796 62532 111800 62588
rect 111736 62528 111800 62532
rect 111816 62588 111880 62592
rect 111816 62532 111820 62588
rect 111820 62532 111876 62588
rect 111876 62532 111880 62588
rect 111816 62528 111880 62532
rect 111896 62588 111960 62592
rect 111896 62532 111900 62588
rect 111900 62532 111956 62588
rect 111956 62532 111960 62588
rect 111896 62528 111960 62532
rect 111976 62588 112040 62592
rect 111976 62532 111980 62588
rect 111980 62532 112036 62588
rect 112036 62532 112040 62588
rect 111976 62528 112040 62532
rect 142456 62588 142520 62592
rect 142456 62532 142460 62588
rect 142460 62532 142516 62588
rect 142516 62532 142520 62588
rect 142456 62528 142520 62532
rect 142536 62588 142600 62592
rect 142536 62532 142540 62588
rect 142540 62532 142596 62588
rect 142596 62532 142600 62588
rect 142536 62528 142600 62532
rect 142616 62588 142680 62592
rect 142616 62532 142620 62588
rect 142620 62532 142676 62588
rect 142676 62532 142680 62588
rect 142616 62528 142680 62532
rect 142696 62588 142760 62592
rect 142696 62532 142700 62588
rect 142700 62532 142756 62588
rect 142756 62532 142760 62588
rect 142696 62528 142760 62532
rect 173176 62588 173240 62592
rect 173176 62532 173180 62588
rect 173180 62532 173236 62588
rect 173236 62532 173240 62588
rect 173176 62528 173240 62532
rect 173256 62588 173320 62592
rect 173256 62532 173260 62588
rect 173260 62532 173316 62588
rect 173316 62532 173320 62588
rect 173256 62528 173320 62532
rect 173336 62588 173400 62592
rect 173336 62532 173340 62588
rect 173340 62532 173396 62588
rect 173396 62532 173400 62588
rect 173336 62528 173400 62532
rect 173416 62588 173480 62592
rect 173416 62532 173420 62588
rect 173420 62532 173476 62588
rect 173476 62532 173480 62588
rect 173416 62528 173480 62532
rect 4216 62044 4280 62048
rect 4216 61988 4220 62044
rect 4220 61988 4276 62044
rect 4276 61988 4280 62044
rect 4216 61984 4280 61988
rect 4296 62044 4360 62048
rect 4296 61988 4300 62044
rect 4300 61988 4356 62044
rect 4356 61988 4360 62044
rect 4296 61984 4360 61988
rect 4376 62044 4440 62048
rect 4376 61988 4380 62044
rect 4380 61988 4436 62044
rect 4436 61988 4440 62044
rect 4376 61984 4440 61988
rect 4456 62044 4520 62048
rect 4456 61988 4460 62044
rect 4460 61988 4516 62044
rect 4516 61988 4520 62044
rect 4456 61984 4520 61988
rect 34936 62044 35000 62048
rect 34936 61988 34940 62044
rect 34940 61988 34996 62044
rect 34996 61988 35000 62044
rect 34936 61984 35000 61988
rect 35016 62044 35080 62048
rect 35016 61988 35020 62044
rect 35020 61988 35076 62044
rect 35076 61988 35080 62044
rect 35016 61984 35080 61988
rect 35096 62044 35160 62048
rect 35096 61988 35100 62044
rect 35100 61988 35156 62044
rect 35156 61988 35160 62044
rect 35096 61984 35160 61988
rect 35176 62044 35240 62048
rect 35176 61988 35180 62044
rect 35180 61988 35236 62044
rect 35236 61988 35240 62044
rect 35176 61984 35240 61988
rect 65656 62044 65720 62048
rect 65656 61988 65660 62044
rect 65660 61988 65716 62044
rect 65716 61988 65720 62044
rect 65656 61984 65720 61988
rect 65736 62044 65800 62048
rect 65736 61988 65740 62044
rect 65740 61988 65796 62044
rect 65796 61988 65800 62044
rect 65736 61984 65800 61988
rect 65816 62044 65880 62048
rect 65816 61988 65820 62044
rect 65820 61988 65876 62044
rect 65876 61988 65880 62044
rect 65816 61984 65880 61988
rect 65896 62044 65960 62048
rect 65896 61988 65900 62044
rect 65900 61988 65956 62044
rect 65956 61988 65960 62044
rect 65896 61984 65960 61988
rect 96376 62044 96440 62048
rect 96376 61988 96380 62044
rect 96380 61988 96436 62044
rect 96436 61988 96440 62044
rect 96376 61984 96440 61988
rect 96456 62044 96520 62048
rect 96456 61988 96460 62044
rect 96460 61988 96516 62044
rect 96516 61988 96520 62044
rect 96456 61984 96520 61988
rect 96536 62044 96600 62048
rect 96536 61988 96540 62044
rect 96540 61988 96596 62044
rect 96596 61988 96600 62044
rect 96536 61984 96600 61988
rect 96616 62044 96680 62048
rect 96616 61988 96620 62044
rect 96620 61988 96676 62044
rect 96676 61988 96680 62044
rect 96616 61984 96680 61988
rect 127096 62044 127160 62048
rect 127096 61988 127100 62044
rect 127100 61988 127156 62044
rect 127156 61988 127160 62044
rect 127096 61984 127160 61988
rect 127176 62044 127240 62048
rect 127176 61988 127180 62044
rect 127180 61988 127236 62044
rect 127236 61988 127240 62044
rect 127176 61984 127240 61988
rect 127256 62044 127320 62048
rect 127256 61988 127260 62044
rect 127260 61988 127316 62044
rect 127316 61988 127320 62044
rect 127256 61984 127320 61988
rect 127336 62044 127400 62048
rect 127336 61988 127340 62044
rect 127340 61988 127396 62044
rect 127396 61988 127400 62044
rect 127336 61984 127400 61988
rect 157816 62044 157880 62048
rect 157816 61988 157820 62044
rect 157820 61988 157876 62044
rect 157876 61988 157880 62044
rect 157816 61984 157880 61988
rect 157896 62044 157960 62048
rect 157896 61988 157900 62044
rect 157900 61988 157956 62044
rect 157956 61988 157960 62044
rect 157896 61984 157960 61988
rect 157976 62044 158040 62048
rect 157976 61988 157980 62044
rect 157980 61988 158036 62044
rect 158036 61988 158040 62044
rect 157976 61984 158040 61988
rect 158056 62044 158120 62048
rect 158056 61988 158060 62044
rect 158060 61988 158116 62044
rect 158116 61988 158120 62044
rect 158056 61984 158120 61988
rect 19576 61500 19640 61504
rect 19576 61444 19580 61500
rect 19580 61444 19636 61500
rect 19636 61444 19640 61500
rect 19576 61440 19640 61444
rect 19656 61500 19720 61504
rect 19656 61444 19660 61500
rect 19660 61444 19716 61500
rect 19716 61444 19720 61500
rect 19656 61440 19720 61444
rect 19736 61500 19800 61504
rect 19736 61444 19740 61500
rect 19740 61444 19796 61500
rect 19796 61444 19800 61500
rect 19736 61440 19800 61444
rect 19816 61500 19880 61504
rect 19816 61444 19820 61500
rect 19820 61444 19876 61500
rect 19876 61444 19880 61500
rect 19816 61440 19880 61444
rect 50296 61500 50360 61504
rect 50296 61444 50300 61500
rect 50300 61444 50356 61500
rect 50356 61444 50360 61500
rect 50296 61440 50360 61444
rect 50376 61500 50440 61504
rect 50376 61444 50380 61500
rect 50380 61444 50436 61500
rect 50436 61444 50440 61500
rect 50376 61440 50440 61444
rect 50456 61500 50520 61504
rect 50456 61444 50460 61500
rect 50460 61444 50516 61500
rect 50516 61444 50520 61500
rect 50456 61440 50520 61444
rect 50536 61500 50600 61504
rect 50536 61444 50540 61500
rect 50540 61444 50596 61500
rect 50596 61444 50600 61500
rect 50536 61440 50600 61444
rect 81016 61500 81080 61504
rect 81016 61444 81020 61500
rect 81020 61444 81076 61500
rect 81076 61444 81080 61500
rect 81016 61440 81080 61444
rect 81096 61500 81160 61504
rect 81096 61444 81100 61500
rect 81100 61444 81156 61500
rect 81156 61444 81160 61500
rect 81096 61440 81160 61444
rect 81176 61500 81240 61504
rect 81176 61444 81180 61500
rect 81180 61444 81236 61500
rect 81236 61444 81240 61500
rect 81176 61440 81240 61444
rect 81256 61500 81320 61504
rect 81256 61444 81260 61500
rect 81260 61444 81316 61500
rect 81316 61444 81320 61500
rect 81256 61440 81320 61444
rect 111736 61500 111800 61504
rect 111736 61444 111740 61500
rect 111740 61444 111796 61500
rect 111796 61444 111800 61500
rect 111736 61440 111800 61444
rect 111816 61500 111880 61504
rect 111816 61444 111820 61500
rect 111820 61444 111876 61500
rect 111876 61444 111880 61500
rect 111816 61440 111880 61444
rect 111896 61500 111960 61504
rect 111896 61444 111900 61500
rect 111900 61444 111956 61500
rect 111956 61444 111960 61500
rect 111896 61440 111960 61444
rect 111976 61500 112040 61504
rect 111976 61444 111980 61500
rect 111980 61444 112036 61500
rect 112036 61444 112040 61500
rect 111976 61440 112040 61444
rect 142456 61500 142520 61504
rect 142456 61444 142460 61500
rect 142460 61444 142516 61500
rect 142516 61444 142520 61500
rect 142456 61440 142520 61444
rect 142536 61500 142600 61504
rect 142536 61444 142540 61500
rect 142540 61444 142596 61500
rect 142596 61444 142600 61500
rect 142536 61440 142600 61444
rect 142616 61500 142680 61504
rect 142616 61444 142620 61500
rect 142620 61444 142676 61500
rect 142676 61444 142680 61500
rect 142616 61440 142680 61444
rect 142696 61500 142760 61504
rect 142696 61444 142700 61500
rect 142700 61444 142756 61500
rect 142756 61444 142760 61500
rect 142696 61440 142760 61444
rect 173176 61500 173240 61504
rect 173176 61444 173180 61500
rect 173180 61444 173236 61500
rect 173236 61444 173240 61500
rect 173176 61440 173240 61444
rect 173256 61500 173320 61504
rect 173256 61444 173260 61500
rect 173260 61444 173316 61500
rect 173316 61444 173320 61500
rect 173256 61440 173320 61444
rect 173336 61500 173400 61504
rect 173336 61444 173340 61500
rect 173340 61444 173396 61500
rect 173396 61444 173400 61500
rect 173336 61440 173400 61444
rect 173416 61500 173480 61504
rect 173416 61444 173420 61500
rect 173420 61444 173476 61500
rect 173476 61444 173480 61500
rect 173416 61440 173480 61444
rect 4216 60956 4280 60960
rect 4216 60900 4220 60956
rect 4220 60900 4276 60956
rect 4276 60900 4280 60956
rect 4216 60896 4280 60900
rect 4296 60956 4360 60960
rect 4296 60900 4300 60956
rect 4300 60900 4356 60956
rect 4356 60900 4360 60956
rect 4296 60896 4360 60900
rect 4376 60956 4440 60960
rect 4376 60900 4380 60956
rect 4380 60900 4436 60956
rect 4436 60900 4440 60956
rect 4376 60896 4440 60900
rect 4456 60956 4520 60960
rect 4456 60900 4460 60956
rect 4460 60900 4516 60956
rect 4516 60900 4520 60956
rect 4456 60896 4520 60900
rect 34936 60956 35000 60960
rect 34936 60900 34940 60956
rect 34940 60900 34996 60956
rect 34996 60900 35000 60956
rect 34936 60896 35000 60900
rect 35016 60956 35080 60960
rect 35016 60900 35020 60956
rect 35020 60900 35076 60956
rect 35076 60900 35080 60956
rect 35016 60896 35080 60900
rect 35096 60956 35160 60960
rect 35096 60900 35100 60956
rect 35100 60900 35156 60956
rect 35156 60900 35160 60956
rect 35096 60896 35160 60900
rect 35176 60956 35240 60960
rect 35176 60900 35180 60956
rect 35180 60900 35236 60956
rect 35236 60900 35240 60956
rect 35176 60896 35240 60900
rect 65656 60956 65720 60960
rect 65656 60900 65660 60956
rect 65660 60900 65716 60956
rect 65716 60900 65720 60956
rect 65656 60896 65720 60900
rect 65736 60956 65800 60960
rect 65736 60900 65740 60956
rect 65740 60900 65796 60956
rect 65796 60900 65800 60956
rect 65736 60896 65800 60900
rect 65816 60956 65880 60960
rect 65816 60900 65820 60956
rect 65820 60900 65876 60956
rect 65876 60900 65880 60956
rect 65816 60896 65880 60900
rect 65896 60956 65960 60960
rect 65896 60900 65900 60956
rect 65900 60900 65956 60956
rect 65956 60900 65960 60956
rect 65896 60896 65960 60900
rect 96376 60956 96440 60960
rect 96376 60900 96380 60956
rect 96380 60900 96436 60956
rect 96436 60900 96440 60956
rect 96376 60896 96440 60900
rect 96456 60956 96520 60960
rect 96456 60900 96460 60956
rect 96460 60900 96516 60956
rect 96516 60900 96520 60956
rect 96456 60896 96520 60900
rect 96536 60956 96600 60960
rect 96536 60900 96540 60956
rect 96540 60900 96596 60956
rect 96596 60900 96600 60956
rect 96536 60896 96600 60900
rect 96616 60956 96680 60960
rect 96616 60900 96620 60956
rect 96620 60900 96676 60956
rect 96676 60900 96680 60956
rect 96616 60896 96680 60900
rect 127096 60956 127160 60960
rect 127096 60900 127100 60956
rect 127100 60900 127156 60956
rect 127156 60900 127160 60956
rect 127096 60896 127160 60900
rect 127176 60956 127240 60960
rect 127176 60900 127180 60956
rect 127180 60900 127236 60956
rect 127236 60900 127240 60956
rect 127176 60896 127240 60900
rect 127256 60956 127320 60960
rect 127256 60900 127260 60956
rect 127260 60900 127316 60956
rect 127316 60900 127320 60956
rect 127256 60896 127320 60900
rect 127336 60956 127400 60960
rect 127336 60900 127340 60956
rect 127340 60900 127396 60956
rect 127396 60900 127400 60956
rect 127336 60896 127400 60900
rect 157816 60956 157880 60960
rect 157816 60900 157820 60956
rect 157820 60900 157876 60956
rect 157876 60900 157880 60956
rect 157816 60896 157880 60900
rect 157896 60956 157960 60960
rect 157896 60900 157900 60956
rect 157900 60900 157956 60956
rect 157956 60900 157960 60956
rect 157896 60896 157960 60900
rect 157976 60956 158040 60960
rect 157976 60900 157980 60956
rect 157980 60900 158036 60956
rect 158036 60900 158040 60956
rect 157976 60896 158040 60900
rect 158056 60956 158120 60960
rect 158056 60900 158060 60956
rect 158060 60900 158116 60956
rect 158116 60900 158120 60956
rect 158056 60896 158120 60900
rect 19576 60412 19640 60416
rect 19576 60356 19580 60412
rect 19580 60356 19636 60412
rect 19636 60356 19640 60412
rect 19576 60352 19640 60356
rect 19656 60412 19720 60416
rect 19656 60356 19660 60412
rect 19660 60356 19716 60412
rect 19716 60356 19720 60412
rect 19656 60352 19720 60356
rect 19736 60412 19800 60416
rect 19736 60356 19740 60412
rect 19740 60356 19796 60412
rect 19796 60356 19800 60412
rect 19736 60352 19800 60356
rect 19816 60412 19880 60416
rect 19816 60356 19820 60412
rect 19820 60356 19876 60412
rect 19876 60356 19880 60412
rect 19816 60352 19880 60356
rect 50296 60412 50360 60416
rect 50296 60356 50300 60412
rect 50300 60356 50356 60412
rect 50356 60356 50360 60412
rect 50296 60352 50360 60356
rect 50376 60412 50440 60416
rect 50376 60356 50380 60412
rect 50380 60356 50436 60412
rect 50436 60356 50440 60412
rect 50376 60352 50440 60356
rect 50456 60412 50520 60416
rect 50456 60356 50460 60412
rect 50460 60356 50516 60412
rect 50516 60356 50520 60412
rect 50456 60352 50520 60356
rect 50536 60412 50600 60416
rect 50536 60356 50540 60412
rect 50540 60356 50596 60412
rect 50596 60356 50600 60412
rect 50536 60352 50600 60356
rect 81016 60412 81080 60416
rect 81016 60356 81020 60412
rect 81020 60356 81076 60412
rect 81076 60356 81080 60412
rect 81016 60352 81080 60356
rect 81096 60412 81160 60416
rect 81096 60356 81100 60412
rect 81100 60356 81156 60412
rect 81156 60356 81160 60412
rect 81096 60352 81160 60356
rect 81176 60412 81240 60416
rect 81176 60356 81180 60412
rect 81180 60356 81236 60412
rect 81236 60356 81240 60412
rect 81176 60352 81240 60356
rect 81256 60412 81320 60416
rect 81256 60356 81260 60412
rect 81260 60356 81316 60412
rect 81316 60356 81320 60412
rect 81256 60352 81320 60356
rect 111736 60412 111800 60416
rect 111736 60356 111740 60412
rect 111740 60356 111796 60412
rect 111796 60356 111800 60412
rect 111736 60352 111800 60356
rect 111816 60412 111880 60416
rect 111816 60356 111820 60412
rect 111820 60356 111876 60412
rect 111876 60356 111880 60412
rect 111816 60352 111880 60356
rect 111896 60412 111960 60416
rect 111896 60356 111900 60412
rect 111900 60356 111956 60412
rect 111956 60356 111960 60412
rect 111896 60352 111960 60356
rect 111976 60412 112040 60416
rect 111976 60356 111980 60412
rect 111980 60356 112036 60412
rect 112036 60356 112040 60412
rect 111976 60352 112040 60356
rect 142456 60412 142520 60416
rect 142456 60356 142460 60412
rect 142460 60356 142516 60412
rect 142516 60356 142520 60412
rect 142456 60352 142520 60356
rect 142536 60412 142600 60416
rect 142536 60356 142540 60412
rect 142540 60356 142596 60412
rect 142596 60356 142600 60412
rect 142536 60352 142600 60356
rect 142616 60412 142680 60416
rect 142616 60356 142620 60412
rect 142620 60356 142676 60412
rect 142676 60356 142680 60412
rect 142616 60352 142680 60356
rect 142696 60412 142760 60416
rect 142696 60356 142700 60412
rect 142700 60356 142756 60412
rect 142756 60356 142760 60412
rect 142696 60352 142760 60356
rect 173176 60412 173240 60416
rect 173176 60356 173180 60412
rect 173180 60356 173236 60412
rect 173236 60356 173240 60412
rect 173176 60352 173240 60356
rect 173256 60412 173320 60416
rect 173256 60356 173260 60412
rect 173260 60356 173316 60412
rect 173316 60356 173320 60412
rect 173256 60352 173320 60356
rect 173336 60412 173400 60416
rect 173336 60356 173340 60412
rect 173340 60356 173396 60412
rect 173396 60356 173400 60412
rect 173336 60352 173400 60356
rect 173416 60412 173480 60416
rect 173416 60356 173420 60412
rect 173420 60356 173476 60412
rect 173476 60356 173480 60412
rect 173416 60352 173480 60356
rect 4216 59868 4280 59872
rect 4216 59812 4220 59868
rect 4220 59812 4276 59868
rect 4276 59812 4280 59868
rect 4216 59808 4280 59812
rect 4296 59868 4360 59872
rect 4296 59812 4300 59868
rect 4300 59812 4356 59868
rect 4356 59812 4360 59868
rect 4296 59808 4360 59812
rect 4376 59868 4440 59872
rect 4376 59812 4380 59868
rect 4380 59812 4436 59868
rect 4436 59812 4440 59868
rect 4376 59808 4440 59812
rect 4456 59868 4520 59872
rect 4456 59812 4460 59868
rect 4460 59812 4516 59868
rect 4516 59812 4520 59868
rect 4456 59808 4520 59812
rect 34936 59868 35000 59872
rect 34936 59812 34940 59868
rect 34940 59812 34996 59868
rect 34996 59812 35000 59868
rect 34936 59808 35000 59812
rect 35016 59868 35080 59872
rect 35016 59812 35020 59868
rect 35020 59812 35076 59868
rect 35076 59812 35080 59868
rect 35016 59808 35080 59812
rect 35096 59868 35160 59872
rect 35096 59812 35100 59868
rect 35100 59812 35156 59868
rect 35156 59812 35160 59868
rect 35096 59808 35160 59812
rect 35176 59868 35240 59872
rect 35176 59812 35180 59868
rect 35180 59812 35236 59868
rect 35236 59812 35240 59868
rect 35176 59808 35240 59812
rect 65656 59868 65720 59872
rect 65656 59812 65660 59868
rect 65660 59812 65716 59868
rect 65716 59812 65720 59868
rect 65656 59808 65720 59812
rect 65736 59868 65800 59872
rect 65736 59812 65740 59868
rect 65740 59812 65796 59868
rect 65796 59812 65800 59868
rect 65736 59808 65800 59812
rect 65816 59868 65880 59872
rect 65816 59812 65820 59868
rect 65820 59812 65876 59868
rect 65876 59812 65880 59868
rect 65816 59808 65880 59812
rect 65896 59868 65960 59872
rect 65896 59812 65900 59868
rect 65900 59812 65956 59868
rect 65956 59812 65960 59868
rect 65896 59808 65960 59812
rect 96376 59868 96440 59872
rect 96376 59812 96380 59868
rect 96380 59812 96436 59868
rect 96436 59812 96440 59868
rect 96376 59808 96440 59812
rect 96456 59868 96520 59872
rect 96456 59812 96460 59868
rect 96460 59812 96516 59868
rect 96516 59812 96520 59868
rect 96456 59808 96520 59812
rect 96536 59868 96600 59872
rect 96536 59812 96540 59868
rect 96540 59812 96596 59868
rect 96596 59812 96600 59868
rect 96536 59808 96600 59812
rect 96616 59868 96680 59872
rect 96616 59812 96620 59868
rect 96620 59812 96676 59868
rect 96676 59812 96680 59868
rect 96616 59808 96680 59812
rect 127096 59868 127160 59872
rect 127096 59812 127100 59868
rect 127100 59812 127156 59868
rect 127156 59812 127160 59868
rect 127096 59808 127160 59812
rect 127176 59868 127240 59872
rect 127176 59812 127180 59868
rect 127180 59812 127236 59868
rect 127236 59812 127240 59868
rect 127176 59808 127240 59812
rect 127256 59868 127320 59872
rect 127256 59812 127260 59868
rect 127260 59812 127316 59868
rect 127316 59812 127320 59868
rect 127256 59808 127320 59812
rect 127336 59868 127400 59872
rect 127336 59812 127340 59868
rect 127340 59812 127396 59868
rect 127396 59812 127400 59868
rect 127336 59808 127400 59812
rect 157816 59868 157880 59872
rect 157816 59812 157820 59868
rect 157820 59812 157876 59868
rect 157876 59812 157880 59868
rect 157816 59808 157880 59812
rect 157896 59868 157960 59872
rect 157896 59812 157900 59868
rect 157900 59812 157956 59868
rect 157956 59812 157960 59868
rect 157896 59808 157960 59812
rect 157976 59868 158040 59872
rect 157976 59812 157980 59868
rect 157980 59812 158036 59868
rect 158036 59812 158040 59868
rect 157976 59808 158040 59812
rect 158056 59868 158120 59872
rect 158056 59812 158060 59868
rect 158060 59812 158116 59868
rect 158116 59812 158120 59868
rect 158056 59808 158120 59812
rect 19576 59324 19640 59328
rect 19576 59268 19580 59324
rect 19580 59268 19636 59324
rect 19636 59268 19640 59324
rect 19576 59264 19640 59268
rect 19656 59324 19720 59328
rect 19656 59268 19660 59324
rect 19660 59268 19716 59324
rect 19716 59268 19720 59324
rect 19656 59264 19720 59268
rect 19736 59324 19800 59328
rect 19736 59268 19740 59324
rect 19740 59268 19796 59324
rect 19796 59268 19800 59324
rect 19736 59264 19800 59268
rect 19816 59324 19880 59328
rect 19816 59268 19820 59324
rect 19820 59268 19876 59324
rect 19876 59268 19880 59324
rect 19816 59264 19880 59268
rect 50296 59324 50360 59328
rect 50296 59268 50300 59324
rect 50300 59268 50356 59324
rect 50356 59268 50360 59324
rect 50296 59264 50360 59268
rect 50376 59324 50440 59328
rect 50376 59268 50380 59324
rect 50380 59268 50436 59324
rect 50436 59268 50440 59324
rect 50376 59264 50440 59268
rect 50456 59324 50520 59328
rect 50456 59268 50460 59324
rect 50460 59268 50516 59324
rect 50516 59268 50520 59324
rect 50456 59264 50520 59268
rect 50536 59324 50600 59328
rect 50536 59268 50540 59324
rect 50540 59268 50596 59324
rect 50596 59268 50600 59324
rect 50536 59264 50600 59268
rect 81016 59324 81080 59328
rect 81016 59268 81020 59324
rect 81020 59268 81076 59324
rect 81076 59268 81080 59324
rect 81016 59264 81080 59268
rect 81096 59324 81160 59328
rect 81096 59268 81100 59324
rect 81100 59268 81156 59324
rect 81156 59268 81160 59324
rect 81096 59264 81160 59268
rect 81176 59324 81240 59328
rect 81176 59268 81180 59324
rect 81180 59268 81236 59324
rect 81236 59268 81240 59324
rect 81176 59264 81240 59268
rect 81256 59324 81320 59328
rect 81256 59268 81260 59324
rect 81260 59268 81316 59324
rect 81316 59268 81320 59324
rect 81256 59264 81320 59268
rect 111736 59324 111800 59328
rect 111736 59268 111740 59324
rect 111740 59268 111796 59324
rect 111796 59268 111800 59324
rect 111736 59264 111800 59268
rect 111816 59324 111880 59328
rect 111816 59268 111820 59324
rect 111820 59268 111876 59324
rect 111876 59268 111880 59324
rect 111816 59264 111880 59268
rect 111896 59324 111960 59328
rect 111896 59268 111900 59324
rect 111900 59268 111956 59324
rect 111956 59268 111960 59324
rect 111896 59264 111960 59268
rect 111976 59324 112040 59328
rect 111976 59268 111980 59324
rect 111980 59268 112036 59324
rect 112036 59268 112040 59324
rect 111976 59264 112040 59268
rect 142456 59324 142520 59328
rect 142456 59268 142460 59324
rect 142460 59268 142516 59324
rect 142516 59268 142520 59324
rect 142456 59264 142520 59268
rect 142536 59324 142600 59328
rect 142536 59268 142540 59324
rect 142540 59268 142596 59324
rect 142596 59268 142600 59324
rect 142536 59264 142600 59268
rect 142616 59324 142680 59328
rect 142616 59268 142620 59324
rect 142620 59268 142676 59324
rect 142676 59268 142680 59324
rect 142616 59264 142680 59268
rect 142696 59324 142760 59328
rect 142696 59268 142700 59324
rect 142700 59268 142756 59324
rect 142756 59268 142760 59324
rect 142696 59264 142760 59268
rect 173176 59324 173240 59328
rect 173176 59268 173180 59324
rect 173180 59268 173236 59324
rect 173236 59268 173240 59324
rect 173176 59264 173240 59268
rect 173256 59324 173320 59328
rect 173256 59268 173260 59324
rect 173260 59268 173316 59324
rect 173316 59268 173320 59324
rect 173256 59264 173320 59268
rect 173336 59324 173400 59328
rect 173336 59268 173340 59324
rect 173340 59268 173396 59324
rect 173396 59268 173400 59324
rect 173336 59264 173400 59268
rect 173416 59324 173480 59328
rect 173416 59268 173420 59324
rect 173420 59268 173476 59324
rect 173476 59268 173480 59324
rect 173416 59264 173480 59268
rect 4216 58780 4280 58784
rect 4216 58724 4220 58780
rect 4220 58724 4276 58780
rect 4276 58724 4280 58780
rect 4216 58720 4280 58724
rect 4296 58780 4360 58784
rect 4296 58724 4300 58780
rect 4300 58724 4356 58780
rect 4356 58724 4360 58780
rect 4296 58720 4360 58724
rect 4376 58780 4440 58784
rect 4376 58724 4380 58780
rect 4380 58724 4436 58780
rect 4436 58724 4440 58780
rect 4376 58720 4440 58724
rect 4456 58780 4520 58784
rect 4456 58724 4460 58780
rect 4460 58724 4516 58780
rect 4516 58724 4520 58780
rect 4456 58720 4520 58724
rect 34936 58780 35000 58784
rect 34936 58724 34940 58780
rect 34940 58724 34996 58780
rect 34996 58724 35000 58780
rect 34936 58720 35000 58724
rect 35016 58780 35080 58784
rect 35016 58724 35020 58780
rect 35020 58724 35076 58780
rect 35076 58724 35080 58780
rect 35016 58720 35080 58724
rect 35096 58780 35160 58784
rect 35096 58724 35100 58780
rect 35100 58724 35156 58780
rect 35156 58724 35160 58780
rect 35096 58720 35160 58724
rect 35176 58780 35240 58784
rect 35176 58724 35180 58780
rect 35180 58724 35236 58780
rect 35236 58724 35240 58780
rect 35176 58720 35240 58724
rect 65656 58780 65720 58784
rect 65656 58724 65660 58780
rect 65660 58724 65716 58780
rect 65716 58724 65720 58780
rect 65656 58720 65720 58724
rect 65736 58780 65800 58784
rect 65736 58724 65740 58780
rect 65740 58724 65796 58780
rect 65796 58724 65800 58780
rect 65736 58720 65800 58724
rect 65816 58780 65880 58784
rect 65816 58724 65820 58780
rect 65820 58724 65876 58780
rect 65876 58724 65880 58780
rect 65816 58720 65880 58724
rect 65896 58780 65960 58784
rect 65896 58724 65900 58780
rect 65900 58724 65956 58780
rect 65956 58724 65960 58780
rect 65896 58720 65960 58724
rect 96376 58780 96440 58784
rect 96376 58724 96380 58780
rect 96380 58724 96436 58780
rect 96436 58724 96440 58780
rect 96376 58720 96440 58724
rect 96456 58780 96520 58784
rect 96456 58724 96460 58780
rect 96460 58724 96516 58780
rect 96516 58724 96520 58780
rect 96456 58720 96520 58724
rect 96536 58780 96600 58784
rect 96536 58724 96540 58780
rect 96540 58724 96596 58780
rect 96596 58724 96600 58780
rect 96536 58720 96600 58724
rect 96616 58780 96680 58784
rect 96616 58724 96620 58780
rect 96620 58724 96676 58780
rect 96676 58724 96680 58780
rect 96616 58720 96680 58724
rect 127096 58780 127160 58784
rect 127096 58724 127100 58780
rect 127100 58724 127156 58780
rect 127156 58724 127160 58780
rect 127096 58720 127160 58724
rect 127176 58780 127240 58784
rect 127176 58724 127180 58780
rect 127180 58724 127236 58780
rect 127236 58724 127240 58780
rect 127176 58720 127240 58724
rect 127256 58780 127320 58784
rect 127256 58724 127260 58780
rect 127260 58724 127316 58780
rect 127316 58724 127320 58780
rect 127256 58720 127320 58724
rect 127336 58780 127400 58784
rect 127336 58724 127340 58780
rect 127340 58724 127396 58780
rect 127396 58724 127400 58780
rect 127336 58720 127400 58724
rect 157816 58780 157880 58784
rect 157816 58724 157820 58780
rect 157820 58724 157876 58780
rect 157876 58724 157880 58780
rect 157816 58720 157880 58724
rect 157896 58780 157960 58784
rect 157896 58724 157900 58780
rect 157900 58724 157956 58780
rect 157956 58724 157960 58780
rect 157896 58720 157960 58724
rect 157976 58780 158040 58784
rect 157976 58724 157980 58780
rect 157980 58724 158036 58780
rect 158036 58724 158040 58780
rect 157976 58720 158040 58724
rect 158056 58780 158120 58784
rect 158056 58724 158060 58780
rect 158060 58724 158116 58780
rect 158116 58724 158120 58780
rect 158056 58720 158120 58724
rect 19576 58236 19640 58240
rect 19576 58180 19580 58236
rect 19580 58180 19636 58236
rect 19636 58180 19640 58236
rect 19576 58176 19640 58180
rect 19656 58236 19720 58240
rect 19656 58180 19660 58236
rect 19660 58180 19716 58236
rect 19716 58180 19720 58236
rect 19656 58176 19720 58180
rect 19736 58236 19800 58240
rect 19736 58180 19740 58236
rect 19740 58180 19796 58236
rect 19796 58180 19800 58236
rect 19736 58176 19800 58180
rect 19816 58236 19880 58240
rect 19816 58180 19820 58236
rect 19820 58180 19876 58236
rect 19876 58180 19880 58236
rect 19816 58176 19880 58180
rect 50296 58236 50360 58240
rect 50296 58180 50300 58236
rect 50300 58180 50356 58236
rect 50356 58180 50360 58236
rect 50296 58176 50360 58180
rect 50376 58236 50440 58240
rect 50376 58180 50380 58236
rect 50380 58180 50436 58236
rect 50436 58180 50440 58236
rect 50376 58176 50440 58180
rect 50456 58236 50520 58240
rect 50456 58180 50460 58236
rect 50460 58180 50516 58236
rect 50516 58180 50520 58236
rect 50456 58176 50520 58180
rect 50536 58236 50600 58240
rect 50536 58180 50540 58236
rect 50540 58180 50596 58236
rect 50596 58180 50600 58236
rect 50536 58176 50600 58180
rect 81016 58236 81080 58240
rect 81016 58180 81020 58236
rect 81020 58180 81076 58236
rect 81076 58180 81080 58236
rect 81016 58176 81080 58180
rect 81096 58236 81160 58240
rect 81096 58180 81100 58236
rect 81100 58180 81156 58236
rect 81156 58180 81160 58236
rect 81096 58176 81160 58180
rect 81176 58236 81240 58240
rect 81176 58180 81180 58236
rect 81180 58180 81236 58236
rect 81236 58180 81240 58236
rect 81176 58176 81240 58180
rect 81256 58236 81320 58240
rect 81256 58180 81260 58236
rect 81260 58180 81316 58236
rect 81316 58180 81320 58236
rect 81256 58176 81320 58180
rect 111736 58236 111800 58240
rect 111736 58180 111740 58236
rect 111740 58180 111796 58236
rect 111796 58180 111800 58236
rect 111736 58176 111800 58180
rect 111816 58236 111880 58240
rect 111816 58180 111820 58236
rect 111820 58180 111876 58236
rect 111876 58180 111880 58236
rect 111816 58176 111880 58180
rect 111896 58236 111960 58240
rect 111896 58180 111900 58236
rect 111900 58180 111956 58236
rect 111956 58180 111960 58236
rect 111896 58176 111960 58180
rect 111976 58236 112040 58240
rect 111976 58180 111980 58236
rect 111980 58180 112036 58236
rect 112036 58180 112040 58236
rect 111976 58176 112040 58180
rect 142456 58236 142520 58240
rect 142456 58180 142460 58236
rect 142460 58180 142516 58236
rect 142516 58180 142520 58236
rect 142456 58176 142520 58180
rect 142536 58236 142600 58240
rect 142536 58180 142540 58236
rect 142540 58180 142596 58236
rect 142596 58180 142600 58236
rect 142536 58176 142600 58180
rect 142616 58236 142680 58240
rect 142616 58180 142620 58236
rect 142620 58180 142676 58236
rect 142676 58180 142680 58236
rect 142616 58176 142680 58180
rect 142696 58236 142760 58240
rect 142696 58180 142700 58236
rect 142700 58180 142756 58236
rect 142756 58180 142760 58236
rect 142696 58176 142760 58180
rect 173176 58236 173240 58240
rect 173176 58180 173180 58236
rect 173180 58180 173236 58236
rect 173236 58180 173240 58236
rect 173176 58176 173240 58180
rect 173256 58236 173320 58240
rect 173256 58180 173260 58236
rect 173260 58180 173316 58236
rect 173316 58180 173320 58236
rect 173256 58176 173320 58180
rect 173336 58236 173400 58240
rect 173336 58180 173340 58236
rect 173340 58180 173396 58236
rect 173396 58180 173400 58236
rect 173336 58176 173400 58180
rect 173416 58236 173480 58240
rect 173416 58180 173420 58236
rect 173420 58180 173476 58236
rect 173476 58180 173480 58236
rect 173416 58176 173480 58180
rect 4216 57692 4280 57696
rect 4216 57636 4220 57692
rect 4220 57636 4276 57692
rect 4276 57636 4280 57692
rect 4216 57632 4280 57636
rect 4296 57692 4360 57696
rect 4296 57636 4300 57692
rect 4300 57636 4356 57692
rect 4356 57636 4360 57692
rect 4296 57632 4360 57636
rect 4376 57692 4440 57696
rect 4376 57636 4380 57692
rect 4380 57636 4436 57692
rect 4436 57636 4440 57692
rect 4376 57632 4440 57636
rect 4456 57692 4520 57696
rect 4456 57636 4460 57692
rect 4460 57636 4516 57692
rect 4516 57636 4520 57692
rect 4456 57632 4520 57636
rect 34936 57692 35000 57696
rect 34936 57636 34940 57692
rect 34940 57636 34996 57692
rect 34996 57636 35000 57692
rect 34936 57632 35000 57636
rect 35016 57692 35080 57696
rect 35016 57636 35020 57692
rect 35020 57636 35076 57692
rect 35076 57636 35080 57692
rect 35016 57632 35080 57636
rect 35096 57692 35160 57696
rect 35096 57636 35100 57692
rect 35100 57636 35156 57692
rect 35156 57636 35160 57692
rect 35096 57632 35160 57636
rect 35176 57692 35240 57696
rect 35176 57636 35180 57692
rect 35180 57636 35236 57692
rect 35236 57636 35240 57692
rect 35176 57632 35240 57636
rect 65656 57692 65720 57696
rect 65656 57636 65660 57692
rect 65660 57636 65716 57692
rect 65716 57636 65720 57692
rect 65656 57632 65720 57636
rect 65736 57692 65800 57696
rect 65736 57636 65740 57692
rect 65740 57636 65796 57692
rect 65796 57636 65800 57692
rect 65736 57632 65800 57636
rect 65816 57692 65880 57696
rect 65816 57636 65820 57692
rect 65820 57636 65876 57692
rect 65876 57636 65880 57692
rect 65816 57632 65880 57636
rect 65896 57692 65960 57696
rect 65896 57636 65900 57692
rect 65900 57636 65956 57692
rect 65956 57636 65960 57692
rect 65896 57632 65960 57636
rect 96376 57692 96440 57696
rect 96376 57636 96380 57692
rect 96380 57636 96436 57692
rect 96436 57636 96440 57692
rect 96376 57632 96440 57636
rect 96456 57692 96520 57696
rect 96456 57636 96460 57692
rect 96460 57636 96516 57692
rect 96516 57636 96520 57692
rect 96456 57632 96520 57636
rect 96536 57692 96600 57696
rect 96536 57636 96540 57692
rect 96540 57636 96596 57692
rect 96596 57636 96600 57692
rect 96536 57632 96600 57636
rect 96616 57692 96680 57696
rect 96616 57636 96620 57692
rect 96620 57636 96676 57692
rect 96676 57636 96680 57692
rect 96616 57632 96680 57636
rect 127096 57692 127160 57696
rect 127096 57636 127100 57692
rect 127100 57636 127156 57692
rect 127156 57636 127160 57692
rect 127096 57632 127160 57636
rect 127176 57692 127240 57696
rect 127176 57636 127180 57692
rect 127180 57636 127236 57692
rect 127236 57636 127240 57692
rect 127176 57632 127240 57636
rect 127256 57692 127320 57696
rect 127256 57636 127260 57692
rect 127260 57636 127316 57692
rect 127316 57636 127320 57692
rect 127256 57632 127320 57636
rect 127336 57692 127400 57696
rect 127336 57636 127340 57692
rect 127340 57636 127396 57692
rect 127396 57636 127400 57692
rect 127336 57632 127400 57636
rect 157816 57692 157880 57696
rect 157816 57636 157820 57692
rect 157820 57636 157876 57692
rect 157876 57636 157880 57692
rect 157816 57632 157880 57636
rect 157896 57692 157960 57696
rect 157896 57636 157900 57692
rect 157900 57636 157956 57692
rect 157956 57636 157960 57692
rect 157896 57632 157960 57636
rect 157976 57692 158040 57696
rect 157976 57636 157980 57692
rect 157980 57636 158036 57692
rect 158036 57636 158040 57692
rect 157976 57632 158040 57636
rect 158056 57692 158120 57696
rect 158056 57636 158060 57692
rect 158060 57636 158116 57692
rect 158116 57636 158120 57692
rect 158056 57632 158120 57636
rect 19576 57148 19640 57152
rect 19576 57092 19580 57148
rect 19580 57092 19636 57148
rect 19636 57092 19640 57148
rect 19576 57088 19640 57092
rect 19656 57148 19720 57152
rect 19656 57092 19660 57148
rect 19660 57092 19716 57148
rect 19716 57092 19720 57148
rect 19656 57088 19720 57092
rect 19736 57148 19800 57152
rect 19736 57092 19740 57148
rect 19740 57092 19796 57148
rect 19796 57092 19800 57148
rect 19736 57088 19800 57092
rect 19816 57148 19880 57152
rect 19816 57092 19820 57148
rect 19820 57092 19876 57148
rect 19876 57092 19880 57148
rect 19816 57088 19880 57092
rect 50296 57148 50360 57152
rect 50296 57092 50300 57148
rect 50300 57092 50356 57148
rect 50356 57092 50360 57148
rect 50296 57088 50360 57092
rect 50376 57148 50440 57152
rect 50376 57092 50380 57148
rect 50380 57092 50436 57148
rect 50436 57092 50440 57148
rect 50376 57088 50440 57092
rect 50456 57148 50520 57152
rect 50456 57092 50460 57148
rect 50460 57092 50516 57148
rect 50516 57092 50520 57148
rect 50456 57088 50520 57092
rect 50536 57148 50600 57152
rect 50536 57092 50540 57148
rect 50540 57092 50596 57148
rect 50596 57092 50600 57148
rect 50536 57088 50600 57092
rect 81016 57148 81080 57152
rect 81016 57092 81020 57148
rect 81020 57092 81076 57148
rect 81076 57092 81080 57148
rect 81016 57088 81080 57092
rect 81096 57148 81160 57152
rect 81096 57092 81100 57148
rect 81100 57092 81156 57148
rect 81156 57092 81160 57148
rect 81096 57088 81160 57092
rect 81176 57148 81240 57152
rect 81176 57092 81180 57148
rect 81180 57092 81236 57148
rect 81236 57092 81240 57148
rect 81176 57088 81240 57092
rect 81256 57148 81320 57152
rect 81256 57092 81260 57148
rect 81260 57092 81316 57148
rect 81316 57092 81320 57148
rect 81256 57088 81320 57092
rect 111736 57148 111800 57152
rect 111736 57092 111740 57148
rect 111740 57092 111796 57148
rect 111796 57092 111800 57148
rect 111736 57088 111800 57092
rect 111816 57148 111880 57152
rect 111816 57092 111820 57148
rect 111820 57092 111876 57148
rect 111876 57092 111880 57148
rect 111816 57088 111880 57092
rect 111896 57148 111960 57152
rect 111896 57092 111900 57148
rect 111900 57092 111956 57148
rect 111956 57092 111960 57148
rect 111896 57088 111960 57092
rect 111976 57148 112040 57152
rect 111976 57092 111980 57148
rect 111980 57092 112036 57148
rect 112036 57092 112040 57148
rect 111976 57088 112040 57092
rect 142456 57148 142520 57152
rect 142456 57092 142460 57148
rect 142460 57092 142516 57148
rect 142516 57092 142520 57148
rect 142456 57088 142520 57092
rect 142536 57148 142600 57152
rect 142536 57092 142540 57148
rect 142540 57092 142596 57148
rect 142596 57092 142600 57148
rect 142536 57088 142600 57092
rect 142616 57148 142680 57152
rect 142616 57092 142620 57148
rect 142620 57092 142676 57148
rect 142676 57092 142680 57148
rect 142616 57088 142680 57092
rect 142696 57148 142760 57152
rect 142696 57092 142700 57148
rect 142700 57092 142756 57148
rect 142756 57092 142760 57148
rect 142696 57088 142760 57092
rect 173176 57148 173240 57152
rect 173176 57092 173180 57148
rect 173180 57092 173236 57148
rect 173236 57092 173240 57148
rect 173176 57088 173240 57092
rect 173256 57148 173320 57152
rect 173256 57092 173260 57148
rect 173260 57092 173316 57148
rect 173316 57092 173320 57148
rect 173256 57088 173320 57092
rect 173336 57148 173400 57152
rect 173336 57092 173340 57148
rect 173340 57092 173396 57148
rect 173396 57092 173400 57148
rect 173336 57088 173400 57092
rect 173416 57148 173480 57152
rect 173416 57092 173420 57148
rect 173420 57092 173476 57148
rect 173476 57092 173480 57148
rect 173416 57088 173480 57092
rect 4216 56604 4280 56608
rect 4216 56548 4220 56604
rect 4220 56548 4276 56604
rect 4276 56548 4280 56604
rect 4216 56544 4280 56548
rect 4296 56604 4360 56608
rect 4296 56548 4300 56604
rect 4300 56548 4356 56604
rect 4356 56548 4360 56604
rect 4296 56544 4360 56548
rect 4376 56604 4440 56608
rect 4376 56548 4380 56604
rect 4380 56548 4436 56604
rect 4436 56548 4440 56604
rect 4376 56544 4440 56548
rect 4456 56604 4520 56608
rect 4456 56548 4460 56604
rect 4460 56548 4516 56604
rect 4516 56548 4520 56604
rect 4456 56544 4520 56548
rect 34936 56604 35000 56608
rect 34936 56548 34940 56604
rect 34940 56548 34996 56604
rect 34996 56548 35000 56604
rect 34936 56544 35000 56548
rect 35016 56604 35080 56608
rect 35016 56548 35020 56604
rect 35020 56548 35076 56604
rect 35076 56548 35080 56604
rect 35016 56544 35080 56548
rect 35096 56604 35160 56608
rect 35096 56548 35100 56604
rect 35100 56548 35156 56604
rect 35156 56548 35160 56604
rect 35096 56544 35160 56548
rect 35176 56604 35240 56608
rect 35176 56548 35180 56604
rect 35180 56548 35236 56604
rect 35236 56548 35240 56604
rect 35176 56544 35240 56548
rect 65656 56604 65720 56608
rect 65656 56548 65660 56604
rect 65660 56548 65716 56604
rect 65716 56548 65720 56604
rect 65656 56544 65720 56548
rect 65736 56604 65800 56608
rect 65736 56548 65740 56604
rect 65740 56548 65796 56604
rect 65796 56548 65800 56604
rect 65736 56544 65800 56548
rect 65816 56604 65880 56608
rect 65816 56548 65820 56604
rect 65820 56548 65876 56604
rect 65876 56548 65880 56604
rect 65816 56544 65880 56548
rect 65896 56604 65960 56608
rect 65896 56548 65900 56604
rect 65900 56548 65956 56604
rect 65956 56548 65960 56604
rect 65896 56544 65960 56548
rect 96376 56604 96440 56608
rect 96376 56548 96380 56604
rect 96380 56548 96436 56604
rect 96436 56548 96440 56604
rect 96376 56544 96440 56548
rect 96456 56604 96520 56608
rect 96456 56548 96460 56604
rect 96460 56548 96516 56604
rect 96516 56548 96520 56604
rect 96456 56544 96520 56548
rect 96536 56604 96600 56608
rect 96536 56548 96540 56604
rect 96540 56548 96596 56604
rect 96596 56548 96600 56604
rect 96536 56544 96600 56548
rect 96616 56604 96680 56608
rect 96616 56548 96620 56604
rect 96620 56548 96676 56604
rect 96676 56548 96680 56604
rect 96616 56544 96680 56548
rect 127096 56604 127160 56608
rect 127096 56548 127100 56604
rect 127100 56548 127156 56604
rect 127156 56548 127160 56604
rect 127096 56544 127160 56548
rect 127176 56604 127240 56608
rect 127176 56548 127180 56604
rect 127180 56548 127236 56604
rect 127236 56548 127240 56604
rect 127176 56544 127240 56548
rect 127256 56604 127320 56608
rect 127256 56548 127260 56604
rect 127260 56548 127316 56604
rect 127316 56548 127320 56604
rect 127256 56544 127320 56548
rect 127336 56604 127400 56608
rect 127336 56548 127340 56604
rect 127340 56548 127396 56604
rect 127396 56548 127400 56604
rect 127336 56544 127400 56548
rect 157816 56604 157880 56608
rect 157816 56548 157820 56604
rect 157820 56548 157876 56604
rect 157876 56548 157880 56604
rect 157816 56544 157880 56548
rect 157896 56604 157960 56608
rect 157896 56548 157900 56604
rect 157900 56548 157956 56604
rect 157956 56548 157960 56604
rect 157896 56544 157960 56548
rect 157976 56604 158040 56608
rect 157976 56548 157980 56604
rect 157980 56548 158036 56604
rect 158036 56548 158040 56604
rect 157976 56544 158040 56548
rect 158056 56604 158120 56608
rect 158056 56548 158060 56604
rect 158060 56548 158116 56604
rect 158116 56548 158120 56604
rect 158056 56544 158120 56548
rect 19576 56060 19640 56064
rect 19576 56004 19580 56060
rect 19580 56004 19636 56060
rect 19636 56004 19640 56060
rect 19576 56000 19640 56004
rect 19656 56060 19720 56064
rect 19656 56004 19660 56060
rect 19660 56004 19716 56060
rect 19716 56004 19720 56060
rect 19656 56000 19720 56004
rect 19736 56060 19800 56064
rect 19736 56004 19740 56060
rect 19740 56004 19796 56060
rect 19796 56004 19800 56060
rect 19736 56000 19800 56004
rect 19816 56060 19880 56064
rect 19816 56004 19820 56060
rect 19820 56004 19876 56060
rect 19876 56004 19880 56060
rect 19816 56000 19880 56004
rect 50296 56060 50360 56064
rect 50296 56004 50300 56060
rect 50300 56004 50356 56060
rect 50356 56004 50360 56060
rect 50296 56000 50360 56004
rect 50376 56060 50440 56064
rect 50376 56004 50380 56060
rect 50380 56004 50436 56060
rect 50436 56004 50440 56060
rect 50376 56000 50440 56004
rect 50456 56060 50520 56064
rect 50456 56004 50460 56060
rect 50460 56004 50516 56060
rect 50516 56004 50520 56060
rect 50456 56000 50520 56004
rect 50536 56060 50600 56064
rect 50536 56004 50540 56060
rect 50540 56004 50596 56060
rect 50596 56004 50600 56060
rect 50536 56000 50600 56004
rect 81016 56060 81080 56064
rect 81016 56004 81020 56060
rect 81020 56004 81076 56060
rect 81076 56004 81080 56060
rect 81016 56000 81080 56004
rect 81096 56060 81160 56064
rect 81096 56004 81100 56060
rect 81100 56004 81156 56060
rect 81156 56004 81160 56060
rect 81096 56000 81160 56004
rect 81176 56060 81240 56064
rect 81176 56004 81180 56060
rect 81180 56004 81236 56060
rect 81236 56004 81240 56060
rect 81176 56000 81240 56004
rect 81256 56060 81320 56064
rect 81256 56004 81260 56060
rect 81260 56004 81316 56060
rect 81316 56004 81320 56060
rect 81256 56000 81320 56004
rect 111736 56060 111800 56064
rect 111736 56004 111740 56060
rect 111740 56004 111796 56060
rect 111796 56004 111800 56060
rect 111736 56000 111800 56004
rect 111816 56060 111880 56064
rect 111816 56004 111820 56060
rect 111820 56004 111876 56060
rect 111876 56004 111880 56060
rect 111816 56000 111880 56004
rect 111896 56060 111960 56064
rect 111896 56004 111900 56060
rect 111900 56004 111956 56060
rect 111956 56004 111960 56060
rect 111896 56000 111960 56004
rect 111976 56060 112040 56064
rect 111976 56004 111980 56060
rect 111980 56004 112036 56060
rect 112036 56004 112040 56060
rect 111976 56000 112040 56004
rect 142456 56060 142520 56064
rect 142456 56004 142460 56060
rect 142460 56004 142516 56060
rect 142516 56004 142520 56060
rect 142456 56000 142520 56004
rect 142536 56060 142600 56064
rect 142536 56004 142540 56060
rect 142540 56004 142596 56060
rect 142596 56004 142600 56060
rect 142536 56000 142600 56004
rect 142616 56060 142680 56064
rect 142616 56004 142620 56060
rect 142620 56004 142676 56060
rect 142676 56004 142680 56060
rect 142616 56000 142680 56004
rect 142696 56060 142760 56064
rect 142696 56004 142700 56060
rect 142700 56004 142756 56060
rect 142756 56004 142760 56060
rect 142696 56000 142760 56004
rect 173176 56060 173240 56064
rect 173176 56004 173180 56060
rect 173180 56004 173236 56060
rect 173236 56004 173240 56060
rect 173176 56000 173240 56004
rect 173256 56060 173320 56064
rect 173256 56004 173260 56060
rect 173260 56004 173316 56060
rect 173316 56004 173320 56060
rect 173256 56000 173320 56004
rect 173336 56060 173400 56064
rect 173336 56004 173340 56060
rect 173340 56004 173396 56060
rect 173396 56004 173400 56060
rect 173336 56000 173400 56004
rect 173416 56060 173480 56064
rect 173416 56004 173420 56060
rect 173420 56004 173476 56060
rect 173476 56004 173480 56060
rect 173416 56000 173480 56004
rect 4216 55516 4280 55520
rect 4216 55460 4220 55516
rect 4220 55460 4276 55516
rect 4276 55460 4280 55516
rect 4216 55456 4280 55460
rect 4296 55516 4360 55520
rect 4296 55460 4300 55516
rect 4300 55460 4356 55516
rect 4356 55460 4360 55516
rect 4296 55456 4360 55460
rect 4376 55516 4440 55520
rect 4376 55460 4380 55516
rect 4380 55460 4436 55516
rect 4436 55460 4440 55516
rect 4376 55456 4440 55460
rect 4456 55516 4520 55520
rect 4456 55460 4460 55516
rect 4460 55460 4516 55516
rect 4516 55460 4520 55516
rect 4456 55456 4520 55460
rect 34936 55516 35000 55520
rect 34936 55460 34940 55516
rect 34940 55460 34996 55516
rect 34996 55460 35000 55516
rect 34936 55456 35000 55460
rect 35016 55516 35080 55520
rect 35016 55460 35020 55516
rect 35020 55460 35076 55516
rect 35076 55460 35080 55516
rect 35016 55456 35080 55460
rect 35096 55516 35160 55520
rect 35096 55460 35100 55516
rect 35100 55460 35156 55516
rect 35156 55460 35160 55516
rect 35096 55456 35160 55460
rect 35176 55516 35240 55520
rect 35176 55460 35180 55516
rect 35180 55460 35236 55516
rect 35236 55460 35240 55516
rect 35176 55456 35240 55460
rect 65656 55516 65720 55520
rect 65656 55460 65660 55516
rect 65660 55460 65716 55516
rect 65716 55460 65720 55516
rect 65656 55456 65720 55460
rect 65736 55516 65800 55520
rect 65736 55460 65740 55516
rect 65740 55460 65796 55516
rect 65796 55460 65800 55516
rect 65736 55456 65800 55460
rect 65816 55516 65880 55520
rect 65816 55460 65820 55516
rect 65820 55460 65876 55516
rect 65876 55460 65880 55516
rect 65816 55456 65880 55460
rect 65896 55516 65960 55520
rect 65896 55460 65900 55516
rect 65900 55460 65956 55516
rect 65956 55460 65960 55516
rect 65896 55456 65960 55460
rect 96376 55516 96440 55520
rect 96376 55460 96380 55516
rect 96380 55460 96436 55516
rect 96436 55460 96440 55516
rect 96376 55456 96440 55460
rect 96456 55516 96520 55520
rect 96456 55460 96460 55516
rect 96460 55460 96516 55516
rect 96516 55460 96520 55516
rect 96456 55456 96520 55460
rect 96536 55516 96600 55520
rect 96536 55460 96540 55516
rect 96540 55460 96596 55516
rect 96596 55460 96600 55516
rect 96536 55456 96600 55460
rect 96616 55516 96680 55520
rect 96616 55460 96620 55516
rect 96620 55460 96676 55516
rect 96676 55460 96680 55516
rect 96616 55456 96680 55460
rect 127096 55516 127160 55520
rect 127096 55460 127100 55516
rect 127100 55460 127156 55516
rect 127156 55460 127160 55516
rect 127096 55456 127160 55460
rect 127176 55516 127240 55520
rect 127176 55460 127180 55516
rect 127180 55460 127236 55516
rect 127236 55460 127240 55516
rect 127176 55456 127240 55460
rect 127256 55516 127320 55520
rect 127256 55460 127260 55516
rect 127260 55460 127316 55516
rect 127316 55460 127320 55516
rect 127256 55456 127320 55460
rect 127336 55516 127400 55520
rect 127336 55460 127340 55516
rect 127340 55460 127396 55516
rect 127396 55460 127400 55516
rect 127336 55456 127400 55460
rect 157816 55516 157880 55520
rect 157816 55460 157820 55516
rect 157820 55460 157876 55516
rect 157876 55460 157880 55516
rect 157816 55456 157880 55460
rect 157896 55516 157960 55520
rect 157896 55460 157900 55516
rect 157900 55460 157956 55516
rect 157956 55460 157960 55516
rect 157896 55456 157960 55460
rect 157976 55516 158040 55520
rect 157976 55460 157980 55516
rect 157980 55460 158036 55516
rect 158036 55460 158040 55516
rect 157976 55456 158040 55460
rect 158056 55516 158120 55520
rect 158056 55460 158060 55516
rect 158060 55460 158116 55516
rect 158116 55460 158120 55516
rect 158056 55456 158120 55460
rect 19576 54972 19640 54976
rect 19576 54916 19580 54972
rect 19580 54916 19636 54972
rect 19636 54916 19640 54972
rect 19576 54912 19640 54916
rect 19656 54972 19720 54976
rect 19656 54916 19660 54972
rect 19660 54916 19716 54972
rect 19716 54916 19720 54972
rect 19656 54912 19720 54916
rect 19736 54972 19800 54976
rect 19736 54916 19740 54972
rect 19740 54916 19796 54972
rect 19796 54916 19800 54972
rect 19736 54912 19800 54916
rect 19816 54972 19880 54976
rect 19816 54916 19820 54972
rect 19820 54916 19876 54972
rect 19876 54916 19880 54972
rect 19816 54912 19880 54916
rect 50296 54972 50360 54976
rect 50296 54916 50300 54972
rect 50300 54916 50356 54972
rect 50356 54916 50360 54972
rect 50296 54912 50360 54916
rect 50376 54972 50440 54976
rect 50376 54916 50380 54972
rect 50380 54916 50436 54972
rect 50436 54916 50440 54972
rect 50376 54912 50440 54916
rect 50456 54972 50520 54976
rect 50456 54916 50460 54972
rect 50460 54916 50516 54972
rect 50516 54916 50520 54972
rect 50456 54912 50520 54916
rect 50536 54972 50600 54976
rect 50536 54916 50540 54972
rect 50540 54916 50596 54972
rect 50596 54916 50600 54972
rect 50536 54912 50600 54916
rect 81016 54972 81080 54976
rect 81016 54916 81020 54972
rect 81020 54916 81076 54972
rect 81076 54916 81080 54972
rect 81016 54912 81080 54916
rect 81096 54972 81160 54976
rect 81096 54916 81100 54972
rect 81100 54916 81156 54972
rect 81156 54916 81160 54972
rect 81096 54912 81160 54916
rect 81176 54972 81240 54976
rect 81176 54916 81180 54972
rect 81180 54916 81236 54972
rect 81236 54916 81240 54972
rect 81176 54912 81240 54916
rect 81256 54972 81320 54976
rect 81256 54916 81260 54972
rect 81260 54916 81316 54972
rect 81316 54916 81320 54972
rect 81256 54912 81320 54916
rect 111736 54972 111800 54976
rect 111736 54916 111740 54972
rect 111740 54916 111796 54972
rect 111796 54916 111800 54972
rect 111736 54912 111800 54916
rect 111816 54972 111880 54976
rect 111816 54916 111820 54972
rect 111820 54916 111876 54972
rect 111876 54916 111880 54972
rect 111816 54912 111880 54916
rect 111896 54972 111960 54976
rect 111896 54916 111900 54972
rect 111900 54916 111956 54972
rect 111956 54916 111960 54972
rect 111896 54912 111960 54916
rect 111976 54972 112040 54976
rect 111976 54916 111980 54972
rect 111980 54916 112036 54972
rect 112036 54916 112040 54972
rect 111976 54912 112040 54916
rect 142456 54972 142520 54976
rect 142456 54916 142460 54972
rect 142460 54916 142516 54972
rect 142516 54916 142520 54972
rect 142456 54912 142520 54916
rect 142536 54972 142600 54976
rect 142536 54916 142540 54972
rect 142540 54916 142596 54972
rect 142596 54916 142600 54972
rect 142536 54912 142600 54916
rect 142616 54972 142680 54976
rect 142616 54916 142620 54972
rect 142620 54916 142676 54972
rect 142676 54916 142680 54972
rect 142616 54912 142680 54916
rect 142696 54972 142760 54976
rect 142696 54916 142700 54972
rect 142700 54916 142756 54972
rect 142756 54916 142760 54972
rect 142696 54912 142760 54916
rect 173176 54972 173240 54976
rect 173176 54916 173180 54972
rect 173180 54916 173236 54972
rect 173236 54916 173240 54972
rect 173176 54912 173240 54916
rect 173256 54972 173320 54976
rect 173256 54916 173260 54972
rect 173260 54916 173316 54972
rect 173316 54916 173320 54972
rect 173256 54912 173320 54916
rect 173336 54972 173400 54976
rect 173336 54916 173340 54972
rect 173340 54916 173396 54972
rect 173396 54916 173400 54972
rect 173336 54912 173400 54916
rect 173416 54972 173480 54976
rect 173416 54916 173420 54972
rect 173420 54916 173476 54972
rect 173476 54916 173480 54972
rect 173416 54912 173480 54916
rect 4216 54428 4280 54432
rect 4216 54372 4220 54428
rect 4220 54372 4276 54428
rect 4276 54372 4280 54428
rect 4216 54368 4280 54372
rect 4296 54428 4360 54432
rect 4296 54372 4300 54428
rect 4300 54372 4356 54428
rect 4356 54372 4360 54428
rect 4296 54368 4360 54372
rect 4376 54428 4440 54432
rect 4376 54372 4380 54428
rect 4380 54372 4436 54428
rect 4436 54372 4440 54428
rect 4376 54368 4440 54372
rect 4456 54428 4520 54432
rect 4456 54372 4460 54428
rect 4460 54372 4516 54428
rect 4516 54372 4520 54428
rect 4456 54368 4520 54372
rect 34936 54428 35000 54432
rect 34936 54372 34940 54428
rect 34940 54372 34996 54428
rect 34996 54372 35000 54428
rect 34936 54368 35000 54372
rect 35016 54428 35080 54432
rect 35016 54372 35020 54428
rect 35020 54372 35076 54428
rect 35076 54372 35080 54428
rect 35016 54368 35080 54372
rect 35096 54428 35160 54432
rect 35096 54372 35100 54428
rect 35100 54372 35156 54428
rect 35156 54372 35160 54428
rect 35096 54368 35160 54372
rect 35176 54428 35240 54432
rect 35176 54372 35180 54428
rect 35180 54372 35236 54428
rect 35236 54372 35240 54428
rect 35176 54368 35240 54372
rect 65656 54428 65720 54432
rect 65656 54372 65660 54428
rect 65660 54372 65716 54428
rect 65716 54372 65720 54428
rect 65656 54368 65720 54372
rect 65736 54428 65800 54432
rect 65736 54372 65740 54428
rect 65740 54372 65796 54428
rect 65796 54372 65800 54428
rect 65736 54368 65800 54372
rect 65816 54428 65880 54432
rect 65816 54372 65820 54428
rect 65820 54372 65876 54428
rect 65876 54372 65880 54428
rect 65816 54368 65880 54372
rect 65896 54428 65960 54432
rect 65896 54372 65900 54428
rect 65900 54372 65956 54428
rect 65956 54372 65960 54428
rect 65896 54368 65960 54372
rect 96376 54428 96440 54432
rect 96376 54372 96380 54428
rect 96380 54372 96436 54428
rect 96436 54372 96440 54428
rect 96376 54368 96440 54372
rect 96456 54428 96520 54432
rect 96456 54372 96460 54428
rect 96460 54372 96516 54428
rect 96516 54372 96520 54428
rect 96456 54368 96520 54372
rect 96536 54428 96600 54432
rect 96536 54372 96540 54428
rect 96540 54372 96596 54428
rect 96596 54372 96600 54428
rect 96536 54368 96600 54372
rect 96616 54428 96680 54432
rect 96616 54372 96620 54428
rect 96620 54372 96676 54428
rect 96676 54372 96680 54428
rect 96616 54368 96680 54372
rect 127096 54428 127160 54432
rect 127096 54372 127100 54428
rect 127100 54372 127156 54428
rect 127156 54372 127160 54428
rect 127096 54368 127160 54372
rect 127176 54428 127240 54432
rect 127176 54372 127180 54428
rect 127180 54372 127236 54428
rect 127236 54372 127240 54428
rect 127176 54368 127240 54372
rect 127256 54428 127320 54432
rect 127256 54372 127260 54428
rect 127260 54372 127316 54428
rect 127316 54372 127320 54428
rect 127256 54368 127320 54372
rect 127336 54428 127400 54432
rect 127336 54372 127340 54428
rect 127340 54372 127396 54428
rect 127396 54372 127400 54428
rect 127336 54368 127400 54372
rect 157816 54428 157880 54432
rect 157816 54372 157820 54428
rect 157820 54372 157876 54428
rect 157876 54372 157880 54428
rect 157816 54368 157880 54372
rect 157896 54428 157960 54432
rect 157896 54372 157900 54428
rect 157900 54372 157956 54428
rect 157956 54372 157960 54428
rect 157896 54368 157960 54372
rect 157976 54428 158040 54432
rect 157976 54372 157980 54428
rect 157980 54372 158036 54428
rect 158036 54372 158040 54428
rect 157976 54368 158040 54372
rect 158056 54428 158120 54432
rect 158056 54372 158060 54428
rect 158060 54372 158116 54428
rect 158116 54372 158120 54428
rect 158056 54368 158120 54372
rect 19576 53884 19640 53888
rect 19576 53828 19580 53884
rect 19580 53828 19636 53884
rect 19636 53828 19640 53884
rect 19576 53824 19640 53828
rect 19656 53884 19720 53888
rect 19656 53828 19660 53884
rect 19660 53828 19716 53884
rect 19716 53828 19720 53884
rect 19656 53824 19720 53828
rect 19736 53884 19800 53888
rect 19736 53828 19740 53884
rect 19740 53828 19796 53884
rect 19796 53828 19800 53884
rect 19736 53824 19800 53828
rect 19816 53884 19880 53888
rect 19816 53828 19820 53884
rect 19820 53828 19876 53884
rect 19876 53828 19880 53884
rect 19816 53824 19880 53828
rect 50296 53884 50360 53888
rect 50296 53828 50300 53884
rect 50300 53828 50356 53884
rect 50356 53828 50360 53884
rect 50296 53824 50360 53828
rect 50376 53884 50440 53888
rect 50376 53828 50380 53884
rect 50380 53828 50436 53884
rect 50436 53828 50440 53884
rect 50376 53824 50440 53828
rect 50456 53884 50520 53888
rect 50456 53828 50460 53884
rect 50460 53828 50516 53884
rect 50516 53828 50520 53884
rect 50456 53824 50520 53828
rect 50536 53884 50600 53888
rect 50536 53828 50540 53884
rect 50540 53828 50596 53884
rect 50596 53828 50600 53884
rect 50536 53824 50600 53828
rect 81016 53884 81080 53888
rect 81016 53828 81020 53884
rect 81020 53828 81076 53884
rect 81076 53828 81080 53884
rect 81016 53824 81080 53828
rect 81096 53884 81160 53888
rect 81096 53828 81100 53884
rect 81100 53828 81156 53884
rect 81156 53828 81160 53884
rect 81096 53824 81160 53828
rect 81176 53884 81240 53888
rect 81176 53828 81180 53884
rect 81180 53828 81236 53884
rect 81236 53828 81240 53884
rect 81176 53824 81240 53828
rect 81256 53884 81320 53888
rect 81256 53828 81260 53884
rect 81260 53828 81316 53884
rect 81316 53828 81320 53884
rect 81256 53824 81320 53828
rect 111736 53884 111800 53888
rect 111736 53828 111740 53884
rect 111740 53828 111796 53884
rect 111796 53828 111800 53884
rect 111736 53824 111800 53828
rect 111816 53884 111880 53888
rect 111816 53828 111820 53884
rect 111820 53828 111876 53884
rect 111876 53828 111880 53884
rect 111816 53824 111880 53828
rect 111896 53884 111960 53888
rect 111896 53828 111900 53884
rect 111900 53828 111956 53884
rect 111956 53828 111960 53884
rect 111896 53824 111960 53828
rect 111976 53884 112040 53888
rect 111976 53828 111980 53884
rect 111980 53828 112036 53884
rect 112036 53828 112040 53884
rect 111976 53824 112040 53828
rect 142456 53884 142520 53888
rect 142456 53828 142460 53884
rect 142460 53828 142516 53884
rect 142516 53828 142520 53884
rect 142456 53824 142520 53828
rect 142536 53884 142600 53888
rect 142536 53828 142540 53884
rect 142540 53828 142596 53884
rect 142596 53828 142600 53884
rect 142536 53824 142600 53828
rect 142616 53884 142680 53888
rect 142616 53828 142620 53884
rect 142620 53828 142676 53884
rect 142676 53828 142680 53884
rect 142616 53824 142680 53828
rect 142696 53884 142760 53888
rect 142696 53828 142700 53884
rect 142700 53828 142756 53884
rect 142756 53828 142760 53884
rect 142696 53824 142760 53828
rect 173176 53884 173240 53888
rect 173176 53828 173180 53884
rect 173180 53828 173236 53884
rect 173236 53828 173240 53884
rect 173176 53824 173240 53828
rect 173256 53884 173320 53888
rect 173256 53828 173260 53884
rect 173260 53828 173316 53884
rect 173316 53828 173320 53884
rect 173256 53824 173320 53828
rect 173336 53884 173400 53888
rect 173336 53828 173340 53884
rect 173340 53828 173396 53884
rect 173396 53828 173400 53884
rect 173336 53824 173400 53828
rect 173416 53884 173480 53888
rect 173416 53828 173420 53884
rect 173420 53828 173476 53884
rect 173476 53828 173480 53884
rect 173416 53824 173480 53828
rect 4216 53340 4280 53344
rect 4216 53284 4220 53340
rect 4220 53284 4276 53340
rect 4276 53284 4280 53340
rect 4216 53280 4280 53284
rect 4296 53340 4360 53344
rect 4296 53284 4300 53340
rect 4300 53284 4356 53340
rect 4356 53284 4360 53340
rect 4296 53280 4360 53284
rect 4376 53340 4440 53344
rect 4376 53284 4380 53340
rect 4380 53284 4436 53340
rect 4436 53284 4440 53340
rect 4376 53280 4440 53284
rect 4456 53340 4520 53344
rect 4456 53284 4460 53340
rect 4460 53284 4516 53340
rect 4516 53284 4520 53340
rect 4456 53280 4520 53284
rect 34936 53340 35000 53344
rect 34936 53284 34940 53340
rect 34940 53284 34996 53340
rect 34996 53284 35000 53340
rect 34936 53280 35000 53284
rect 35016 53340 35080 53344
rect 35016 53284 35020 53340
rect 35020 53284 35076 53340
rect 35076 53284 35080 53340
rect 35016 53280 35080 53284
rect 35096 53340 35160 53344
rect 35096 53284 35100 53340
rect 35100 53284 35156 53340
rect 35156 53284 35160 53340
rect 35096 53280 35160 53284
rect 35176 53340 35240 53344
rect 35176 53284 35180 53340
rect 35180 53284 35236 53340
rect 35236 53284 35240 53340
rect 35176 53280 35240 53284
rect 65656 53340 65720 53344
rect 65656 53284 65660 53340
rect 65660 53284 65716 53340
rect 65716 53284 65720 53340
rect 65656 53280 65720 53284
rect 65736 53340 65800 53344
rect 65736 53284 65740 53340
rect 65740 53284 65796 53340
rect 65796 53284 65800 53340
rect 65736 53280 65800 53284
rect 65816 53340 65880 53344
rect 65816 53284 65820 53340
rect 65820 53284 65876 53340
rect 65876 53284 65880 53340
rect 65816 53280 65880 53284
rect 65896 53340 65960 53344
rect 65896 53284 65900 53340
rect 65900 53284 65956 53340
rect 65956 53284 65960 53340
rect 65896 53280 65960 53284
rect 96376 53340 96440 53344
rect 96376 53284 96380 53340
rect 96380 53284 96436 53340
rect 96436 53284 96440 53340
rect 96376 53280 96440 53284
rect 96456 53340 96520 53344
rect 96456 53284 96460 53340
rect 96460 53284 96516 53340
rect 96516 53284 96520 53340
rect 96456 53280 96520 53284
rect 96536 53340 96600 53344
rect 96536 53284 96540 53340
rect 96540 53284 96596 53340
rect 96596 53284 96600 53340
rect 96536 53280 96600 53284
rect 96616 53340 96680 53344
rect 96616 53284 96620 53340
rect 96620 53284 96676 53340
rect 96676 53284 96680 53340
rect 96616 53280 96680 53284
rect 127096 53340 127160 53344
rect 127096 53284 127100 53340
rect 127100 53284 127156 53340
rect 127156 53284 127160 53340
rect 127096 53280 127160 53284
rect 127176 53340 127240 53344
rect 127176 53284 127180 53340
rect 127180 53284 127236 53340
rect 127236 53284 127240 53340
rect 127176 53280 127240 53284
rect 127256 53340 127320 53344
rect 127256 53284 127260 53340
rect 127260 53284 127316 53340
rect 127316 53284 127320 53340
rect 127256 53280 127320 53284
rect 127336 53340 127400 53344
rect 127336 53284 127340 53340
rect 127340 53284 127396 53340
rect 127396 53284 127400 53340
rect 127336 53280 127400 53284
rect 157816 53340 157880 53344
rect 157816 53284 157820 53340
rect 157820 53284 157876 53340
rect 157876 53284 157880 53340
rect 157816 53280 157880 53284
rect 157896 53340 157960 53344
rect 157896 53284 157900 53340
rect 157900 53284 157956 53340
rect 157956 53284 157960 53340
rect 157896 53280 157960 53284
rect 157976 53340 158040 53344
rect 157976 53284 157980 53340
rect 157980 53284 158036 53340
rect 158036 53284 158040 53340
rect 157976 53280 158040 53284
rect 158056 53340 158120 53344
rect 158056 53284 158060 53340
rect 158060 53284 158116 53340
rect 158116 53284 158120 53340
rect 158056 53280 158120 53284
rect 19576 52796 19640 52800
rect 19576 52740 19580 52796
rect 19580 52740 19636 52796
rect 19636 52740 19640 52796
rect 19576 52736 19640 52740
rect 19656 52796 19720 52800
rect 19656 52740 19660 52796
rect 19660 52740 19716 52796
rect 19716 52740 19720 52796
rect 19656 52736 19720 52740
rect 19736 52796 19800 52800
rect 19736 52740 19740 52796
rect 19740 52740 19796 52796
rect 19796 52740 19800 52796
rect 19736 52736 19800 52740
rect 19816 52796 19880 52800
rect 19816 52740 19820 52796
rect 19820 52740 19876 52796
rect 19876 52740 19880 52796
rect 19816 52736 19880 52740
rect 50296 52796 50360 52800
rect 50296 52740 50300 52796
rect 50300 52740 50356 52796
rect 50356 52740 50360 52796
rect 50296 52736 50360 52740
rect 50376 52796 50440 52800
rect 50376 52740 50380 52796
rect 50380 52740 50436 52796
rect 50436 52740 50440 52796
rect 50376 52736 50440 52740
rect 50456 52796 50520 52800
rect 50456 52740 50460 52796
rect 50460 52740 50516 52796
rect 50516 52740 50520 52796
rect 50456 52736 50520 52740
rect 50536 52796 50600 52800
rect 50536 52740 50540 52796
rect 50540 52740 50596 52796
rect 50596 52740 50600 52796
rect 50536 52736 50600 52740
rect 81016 52796 81080 52800
rect 81016 52740 81020 52796
rect 81020 52740 81076 52796
rect 81076 52740 81080 52796
rect 81016 52736 81080 52740
rect 81096 52796 81160 52800
rect 81096 52740 81100 52796
rect 81100 52740 81156 52796
rect 81156 52740 81160 52796
rect 81096 52736 81160 52740
rect 81176 52796 81240 52800
rect 81176 52740 81180 52796
rect 81180 52740 81236 52796
rect 81236 52740 81240 52796
rect 81176 52736 81240 52740
rect 81256 52796 81320 52800
rect 81256 52740 81260 52796
rect 81260 52740 81316 52796
rect 81316 52740 81320 52796
rect 81256 52736 81320 52740
rect 111736 52796 111800 52800
rect 111736 52740 111740 52796
rect 111740 52740 111796 52796
rect 111796 52740 111800 52796
rect 111736 52736 111800 52740
rect 111816 52796 111880 52800
rect 111816 52740 111820 52796
rect 111820 52740 111876 52796
rect 111876 52740 111880 52796
rect 111816 52736 111880 52740
rect 111896 52796 111960 52800
rect 111896 52740 111900 52796
rect 111900 52740 111956 52796
rect 111956 52740 111960 52796
rect 111896 52736 111960 52740
rect 111976 52796 112040 52800
rect 111976 52740 111980 52796
rect 111980 52740 112036 52796
rect 112036 52740 112040 52796
rect 111976 52736 112040 52740
rect 142456 52796 142520 52800
rect 142456 52740 142460 52796
rect 142460 52740 142516 52796
rect 142516 52740 142520 52796
rect 142456 52736 142520 52740
rect 142536 52796 142600 52800
rect 142536 52740 142540 52796
rect 142540 52740 142596 52796
rect 142596 52740 142600 52796
rect 142536 52736 142600 52740
rect 142616 52796 142680 52800
rect 142616 52740 142620 52796
rect 142620 52740 142676 52796
rect 142676 52740 142680 52796
rect 142616 52736 142680 52740
rect 142696 52796 142760 52800
rect 142696 52740 142700 52796
rect 142700 52740 142756 52796
rect 142756 52740 142760 52796
rect 142696 52736 142760 52740
rect 173176 52796 173240 52800
rect 173176 52740 173180 52796
rect 173180 52740 173236 52796
rect 173236 52740 173240 52796
rect 173176 52736 173240 52740
rect 173256 52796 173320 52800
rect 173256 52740 173260 52796
rect 173260 52740 173316 52796
rect 173316 52740 173320 52796
rect 173256 52736 173320 52740
rect 173336 52796 173400 52800
rect 173336 52740 173340 52796
rect 173340 52740 173396 52796
rect 173396 52740 173400 52796
rect 173336 52736 173400 52740
rect 173416 52796 173480 52800
rect 173416 52740 173420 52796
rect 173420 52740 173476 52796
rect 173476 52740 173480 52796
rect 173416 52736 173480 52740
rect 4216 52252 4280 52256
rect 4216 52196 4220 52252
rect 4220 52196 4276 52252
rect 4276 52196 4280 52252
rect 4216 52192 4280 52196
rect 4296 52252 4360 52256
rect 4296 52196 4300 52252
rect 4300 52196 4356 52252
rect 4356 52196 4360 52252
rect 4296 52192 4360 52196
rect 4376 52252 4440 52256
rect 4376 52196 4380 52252
rect 4380 52196 4436 52252
rect 4436 52196 4440 52252
rect 4376 52192 4440 52196
rect 4456 52252 4520 52256
rect 4456 52196 4460 52252
rect 4460 52196 4516 52252
rect 4516 52196 4520 52252
rect 4456 52192 4520 52196
rect 34936 52252 35000 52256
rect 34936 52196 34940 52252
rect 34940 52196 34996 52252
rect 34996 52196 35000 52252
rect 34936 52192 35000 52196
rect 35016 52252 35080 52256
rect 35016 52196 35020 52252
rect 35020 52196 35076 52252
rect 35076 52196 35080 52252
rect 35016 52192 35080 52196
rect 35096 52252 35160 52256
rect 35096 52196 35100 52252
rect 35100 52196 35156 52252
rect 35156 52196 35160 52252
rect 35096 52192 35160 52196
rect 35176 52252 35240 52256
rect 35176 52196 35180 52252
rect 35180 52196 35236 52252
rect 35236 52196 35240 52252
rect 35176 52192 35240 52196
rect 65656 52252 65720 52256
rect 65656 52196 65660 52252
rect 65660 52196 65716 52252
rect 65716 52196 65720 52252
rect 65656 52192 65720 52196
rect 65736 52252 65800 52256
rect 65736 52196 65740 52252
rect 65740 52196 65796 52252
rect 65796 52196 65800 52252
rect 65736 52192 65800 52196
rect 65816 52252 65880 52256
rect 65816 52196 65820 52252
rect 65820 52196 65876 52252
rect 65876 52196 65880 52252
rect 65816 52192 65880 52196
rect 65896 52252 65960 52256
rect 65896 52196 65900 52252
rect 65900 52196 65956 52252
rect 65956 52196 65960 52252
rect 65896 52192 65960 52196
rect 96376 52252 96440 52256
rect 96376 52196 96380 52252
rect 96380 52196 96436 52252
rect 96436 52196 96440 52252
rect 96376 52192 96440 52196
rect 96456 52252 96520 52256
rect 96456 52196 96460 52252
rect 96460 52196 96516 52252
rect 96516 52196 96520 52252
rect 96456 52192 96520 52196
rect 96536 52252 96600 52256
rect 96536 52196 96540 52252
rect 96540 52196 96596 52252
rect 96596 52196 96600 52252
rect 96536 52192 96600 52196
rect 96616 52252 96680 52256
rect 96616 52196 96620 52252
rect 96620 52196 96676 52252
rect 96676 52196 96680 52252
rect 96616 52192 96680 52196
rect 127096 52252 127160 52256
rect 127096 52196 127100 52252
rect 127100 52196 127156 52252
rect 127156 52196 127160 52252
rect 127096 52192 127160 52196
rect 127176 52252 127240 52256
rect 127176 52196 127180 52252
rect 127180 52196 127236 52252
rect 127236 52196 127240 52252
rect 127176 52192 127240 52196
rect 127256 52252 127320 52256
rect 127256 52196 127260 52252
rect 127260 52196 127316 52252
rect 127316 52196 127320 52252
rect 127256 52192 127320 52196
rect 127336 52252 127400 52256
rect 127336 52196 127340 52252
rect 127340 52196 127396 52252
rect 127396 52196 127400 52252
rect 127336 52192 127400 52196
rect 157816 52252 157880 52256
rect 157816 52196 157820 52252
rect 157820 52196 157876 52252
rect 157876 52196 157880 52252
rect 157816 52192 157880 52196
rect 157896 52252 157960 52256
rect 157896 52196 157900 52252
rect 157900 52196 157956 52252
rect 157956 52196 157960 52252
rect 157896 52192 157960 52196
rect 157976 52252 158040 52256
rect 157976 52196 157980 52252
rect 157980 52196 158036 52252
rect 158036 52196 158040 52252
rect 157976 52192 158040 52196
rect 158056 52252 158120 52256
rect 158056 52196 158060 52252
rect 158060 52196 158116 52252
rect 158116 52196 158120 52252
rect 158056 52192 158120 52196
rect 19576 51708 19640 51712
rect 19576 51652 19580 51708
rect 19580 51652 19636 51708
rect 19636 51652 19640 51708
rect 19576 51648 19640 51652
rect 19656 51708 19720 51712
rect 19656 51652 19660 51708
rect 19660 51652 19716 51708
rect 19716 51652 19720 51708
rect 19656 51648 19720 51652
rect 19736 51708 19800 51712
rect 19736 51652 19740 51708
rect 19740 51652 19796 51708
rect 19796 51652 19800 51708
rect 19736 51648 19800 51652
rect 19816 51708 19880 51712
rect 19816 51652 19820 51708
rect 19820 51652 19876 51708
rect 19876 51652 19880 51708
rect 19816 51648 19880 51652
rect 50296 51708 50360 51712
rect 50296 51652 50300 51708
rect 50300 51652 50356 51708
rect 50356 51652 50360 51708
rect 50296 51648 50360 51652
rect 50376 51708 50440 51712
rect 50376 51652 50380 51708
rect 50380 51652 50436 51708
rect 50436 51652 50440 51708
rect 50376 51648 50440 51652
rect 50456 51708 50520 51712
rect 50456 51652 50460 51708
rect 50460 51652 50516 51708
rect 50516 51652 50520 51708
rect 50456 51648 50520 51652
rect 50536 51708 50600 51712
rect 50536 51652 50540 51708
rect 50540 51652 50596 51708
rect 50596 51652 50600 51708
rect 50536 51648 50600 51652
rect 81016 51708 81080 51712
rect 81016 51652 81020 51708
rect 81020 51652 81076 51708
rect 81076 51652 81080 51708
rect 81016 51648 81080 51652
rect 81096 51708 81160 51712
rect 81096 51652 81100 51708
rect 81100 51652 81156 51708
rect 81156 51652 81160 51708
rect 81096 51648 81160 51652
rect 81176 51708 81240 51712
rect 81176 51652 81180 51708
rect 81180 51652 81236 51708
rect 81236 51652 81240 51708
rect 81176 51648 81240 51652
rect 81256 51708 81320 51712
rect 81256 51652 81260 51708
rect 81260 51652 81316 51708
rect 81316 51652 81320 51708
rect 81256 51648 81320 51652
rect 111736 51708 111800 51712
rect 111736 51652 111740 51708
rect 111740 51652 111796 51708
rect 111796 51652 111800 51708
rect 111736 51648 111800 51652
rect 111816 51708 111880 51712
rect 111816 51652 111820 51708
rect 111820 51652 111876 51708
rect 111876 51652 111880 51708
rect 111816 51648 111880 51652
rect 111896 51708 111960 51712
rect 111896 51652 111900 51708
rect 111900 51652 111956 51708
rect 111956 51652 111960 51708
rect 111896 51648 111960 51652
rect 111976 51708 112040 51712
rect 111976 51652 111980 51708
rect 111980 51652 112036 51708
rect 112036 51652 112040 51708
rect 111976 51648 112040 51652
rect 142456 51708 142520 51712
rect 142456 51652 142460 51708
rect 142460 51652 142516 51708
rect 142516 51652 142520 51708
rect 142456 51648 142520 51652
rect 142536 51708 142600 51712
rect 142536 51652 142540 51708
rect 142540 51652 142596 51708
rect 142596 51652 142600 51708
rect 142536 51648 142600 51652
rect 142616 51708 142680 51712
rect 142616 51652 142620 51708
rect 142620 51652 142676 51708
rect 142676 51652 142680 51708
rect 142616 51648 142680 51652
rect 142696 51708 142760 51712
rect 142696 51652 142700 51708
rect 142700 51652 142756 51708
rect 142756 51652 142760 51708
rect 142696 51648 142760 51652
rect 173176 51708 173240 51712
rect 173176 51652 173180 51708
rect 173180 51652 173236 51708
rect 173236 51652 173240 51708
rect 173176 51648 173240 51652
rect 173256 51708 173320 51712
rect 173256 51652 173260 51708
rect 173260 51652 173316 51708
rect 173316 51652 173320 51708
rect 173256 51648 173320 51652
rect 173336 51708 173400 51712
rect 173336 51652 173340 51708
rect 173340 51652 173396 51708
rect 173396 51652 173400 51708
rect 173336 51648 173400 51652
rect 173416 51708 173480 51712
rect 173416 51652 173420 51708
rect 173420 51652 173476 51708
rect 173476 51652 173480 51708
rect 173416 51648 173480 51652
rect 4216 51164 4280 51168
rect 4216 51108 4220 51164
rect 4220 51108 4276 51164
rect 4276 51108 4280 51164
rect 4216 51104 4280 51108
rect 4296 51164 4360 51168
rect 4296 51108 4300 51164
rect 4300 51108 4356 51164
rect 4356 51108 4360 51164
rect 4296 51104 4360 51108
rect 4376 51164 4440 51168
rect 4376 51108 4380 51164
rect 4380 51108 4436 51164
rect 4436 51108 4440 51164
rect 4376 51104 4440 51108
rect 4456 51164 4520 51168
rect 4456 51108 4460 51164
rect 4460 51108 4516 51164
rect 4516 51108 4520 51164
rect 4456 51104 4520 51108
rect 34936 51164 35000 51168
rect 34936 51108 34940 51164
rect 34940 51108 34996 51164
rect 34996 51108 35000 51164
rect 34936 51104 35000 51108
rect 35016 51164 35080 51168
rect 35016 51108 35020 51164
rect 35020 51108 35076 51164
rect 35076 51108 35080 51164
rect 35016 51104 35080 51108
rect 35096 51164 35160 51168
rect 35096 51108 35100 51164
rect 35100 51108 35156 51164
rect 35156 51108 35160 51164
rect 35096 51104 35160 51108
rect 35176 51164 35240 51168
rect 35176 51108 35180 51164
rect 35180 51108 35236 51164
rect 35236 51108 35240 51164
rect 35176 51104 35240 51108
rect 65656 51164 65720 51168
rect 65656 51108 65660 51164
rect 65660 51108 65716 51164
rect 65716 51108 65720 51164
rect 65656 51104 65720 51108
rect 65736 51164 65800 51168
rect 65736 51108 65740 51164
rect 65740 51108 65796 51164
rect 65796 51108 65800 51164
rect 65736 51104 65800 51108
rect 65816 51164 65880 51168
rect 65816 51108 65820 51164
rect 65820 51108 65876 51164
rect 65876 51108 65880 51164
rect 65816 51104 65880 51108
rect 65896 51164 65960 51168
rect 65896 51108 65900 51164
rect 65900 51108 65956 51164
rect 65956 51108 65960 51164
rect 65896 51104 65960 51108
rect 96376 51164 96440 51168
rect 96376 51108 96380 51164
rect 96380 51108 96436 51164
rect 96436 51108 96440 51164
rect 96376 51104 96440 51108
rect 96456 51164 96520 51168
rect 96456 51108 96460 51164
rect 96460 51108 96516 51164
rect 96516 51108 96520 51164
rect 96456 51104 96520 51108
rect 96536 51164 96600 51168
rect 96536 51108 96540 51164
rect 96540 51108 96596 51164
rect 96596 51108 96600 51164
rect 96536 51104 96600 51108
rect 96616 51164 96680 51168
rect 96616 51108 96620 51164
rect 96620 51108 96676 51164
rect 96676 51108 96680 51164
rect 96616 51104 96680 51108
rect 127096 51164 127160 51168
rect 127096 51108 127100 51164
rect 127100 51108 127156 51164
rect 127156 51108 127160 51164
rect 127096 51104 127160 51108
rect 127176 51164 127240 51168
rect 127176 51108 127180 51164
rect 127180 51108 127236 51164
rect 127236 51108 127240 51164
rect 127176 51104 127240 51108
rect 127256 51164 127320 51168
rect 127256 51108 127260 51164
rect 127260 51108 127316 51164
rect 127316 51108 127320 51164
rect 127256 51104 127320 51108
rect 127336 51164 127400 51168
rect 127336 51108 127340 51164
rect 127340 51108 127396 51164
rect 127396 51108 127400 51164
rect 127336 51104 127400 51108
rect 157816 51164 157880 51168
rect 157816 51108 157820 51164
rect 157820 51108 157876 51164
rect 157876 51108 157880 51164
rect 157816 51104 157880 51108
rect 157896 51164 157960 51168
rect 157896 51108 157900 51164
rect 157900 51108 157956 51164
rect 157956 51108 157960 51164
rect 157896 51104 157960 51108
rect 157976 51164 158040 51168
rect 157976 51108 157980 51164
rect 157980 51108 158036 51164
rect 158036 51108 158040 51164
rect 157976 51104 158040 51108
rect 158056 51164 158120 51168
rect 158056 51108 158060 51164
rect 158060 51108 158116 51164
rect 158116 51108 158120 51164
rect 158056 51104 158120 51108
rect 19576 50620 19640 50624
rect 19576 50564 19580 50620
rect 19580 50564 19636 50620
rect 19636 50564 19640 50620
rect 19576 50560 19640 50564
rect 19656 50620 19720 50624
rect 19656 50564 19660 50620
rect 19660 50564 19716 50620
rect 19716 50564 19720 50620
rect 19656 50560 19720 50564
rect 19736 50620 19800 50624
rect 19736 50564 19740 50620
rect 19740 50564 19796 50620
rect 19796 50564 19800 50620
rect 19736 50560 19800 50564
rect 19816 50620 19880 50624
rect 19816 50564 19820 50620
rect 19820 50564 19876 50620
rect 19876 50564 19880 50620
rect 19816 50560 19880 50564
rect 50296 50620 50360 50624
rect 50296 50564 50300 50620
rect 50300 50564 50356 50620
rect 50356 50564 50360 50620
rect 50296 50560 50360 50564
rect 50376 50620 50440 50624
rect 50376 50564 50380 50620
rect 50380 50564 50436 50620
rect 50436 50564 50440 50620
rect 50376 50560 50440 50564
rect 50456 50620 50520 50624
rect 50456 50564 50460 50620
rect 50460 50564 50516 50620
rect 50516 50564 50520 50620
rect 50456 50560 50520 50564
rect 50536 50620 50600 50624
rect 50536 50564 50540 50620
rect 50540 50564 50596 50620
rect 50596 50564 50600 50620
rect 50536 50560 50600 50564
rect 81016 50620 81080 50624
rect 81016 50564 81020 50620
rect 81020 50564 81076 50620
rect 81076 50564 81080 50620
rect 81016 50560 81080 50564
rect 81096 50620 81160 50624
rect 81096 50564 81100 50620
rect 81100 50564 81156 50620
rect 81156 50564 81160 50620
rect 81096 50560 81160 50564
rect 81176 50620 81240 50624
rect 81176 50564 81180 50620
rect 81180 50564 81236 50620
rect 81236 50564 81240 50620
rect 81176 50560 81240 50564
rect 81256 50620 81320 50624
rect 81256 50564 81260 50620
rect 81260 50564 81316 50620
rect 81316 50564 81320 50620
rect 81256 50560 81320 50564
rect 111736 50620 111800 50624
rect 111736 50564 111740 50620
rect 111740 50564 111796 50620
rect 111796 50564 111800 50620
rect 111736 50560 111800 50564
rect 111816 50620 111880 50624
rect 111816 50564 111820 50620
rect 111820 50564 111876 50620
rect 111876 50564 111880 50620
rect 111816 50560 111880 50564
rect 111896 50620 111960 50624
rect 111896 50564 111900 50620
rect 111900 50564 111956 50620
rect 111956 50564 111960 50620
rect 111896 50560 111960 50564
rect 111976 50620 112040 50624
rect 111976 50564 111980 50620
rect 111980 50564 112036 50620
rect 112036 50564 112040 50620
rect 111976 50560 112040 50564
rect 142456 50620 142520 50624
rect 142456 50564 142460 50620
rect 142460 50564 142516 50620
rect 142516 50564 142520 50620
rect 142456 50560 142520 50564
rect 142536 50620 142600 50624
rect 142536 50564 142540 50620
rect 142540 50564 142596 50620
rect 142596 50564 142600 50620
rect 142536 50560 142600 50564
rect 142616 50620 142680 50624
rect 142616 50564 142620 50620
rect 142620 50564 142676 50620
rect 142676 50564 142680 50620
rect 142616 50560 142680 50564
rect 142696 50620 142760 50624
rect 142696 50564 142700 50620
rect 142700 50564 142756 50620
rect 142756 50564 142760 50620
rect 142696 50560 142760 50564
rect 173176 50620 173240 50624
rect 173176 50564 173180 50620
rect 173180 50564 173236 50620
rect 173236 50564 173240 50620
rect 173176 50560 173240 50564
rect 173256 50620 173320 50624
rect 173256 50564 173260 50620
rect 173260 50564 173316 50620
rect 173316 50564 173320 50620
rect 173256 50560 173320 50564
rect 173336 50620 173400 50624
rect 173336 50564 173340 50620
rect 173340 50564 173396 50620
rect 173396 50564 173400 50620
rect 173336 50560 173400 50564
rect 173416 50620 173480 50624
rect 173416 50564 173420 50620
rect 173420 50564 173476 50620
rect 173476 50564 173480 50620
rect 173416 50560 173480 50564
rect 4216 50076 4280 50080
rect 4216 50020 4220 50076
rect 4220 50020 4276 50076
rect 4276 50020 4280 50076
rect 4216 50016 4280 50020
rect 4296 50076 4360 50080
rect 4296 50020 4300 50076
rect 4300 50020 4356 50076
rect 4356 50020 4360 50076
rect 4296 50016 4360 50020
rect 4376 50076 4440 50080
rect 4376 50020 4380 50076
rect 4380 50020 4436 50076
rect 4436 50020 4440 50076
rect 4376 50016 4440 50020
rect 4456 50076 4520 50080
rect 4456 50020 4460 50076
rect 4460 50020 4516 50076
rect 4516 50020 4520 50076
rect 4456 50016 4520 50020
rect 34936 50076 35000 50080
rect 34936 50020 34940 50076
rect 34940 50020 34996 50076
rect 34996 50020 35000 50076
rect 34936 50016 35000 50020
rect 35016 50076 35080 50080
rect 35016 50020 35020 50076
rect 35020 50020 35076 50076
rect 35076 50020 35080 50076
rect 35016 50016 35080 50020
rect 35096 50076 35160 50080
rect 35096 50020 35100 50076
rect 35100 50020 35156 50076
rect 35156 50020 35160 50076
rect 35096 50016 35160 50020
rect 35176 50076 35240 50080
rect 35176 50020 35180 50076
rect 35180 50020 35236 50076
rect 35236 50020 35240 50076
rect 35176 50016 35240 50020
rect 65656 50076 65720 50080
rect 65656 50020 65660 50076
rect 65660 50020 65716 50076
rect 65716 50020 65720 50076
rect 65656 50016 65720 50020
rect 65736 50076 65800 50080
rect 65736 50020 65740 50076
rect 65740 50020 65796 50076
rect 65796 50020 65800 50076
rect 65736 50016 65800 50020
rect 65816 50076 65880 50080
rect 65816 50020 65820 50076
rect 65820 50020 65876 50076
rect 65876 50020 65880 50076
rect 65816 50016 65880 50020
rect 65896 50076 65960 50080
rect 65896 50020 65900 50076
rect 65900 50020 65956 50076
rect 65956 50020 65960 50076
rect 65896 50016 65960 50020
rect 96376 50076 96440 50080
rect 96376 50020 96380 50076
rect 96380 50020 96436 50076
rect 96436 50020 96440 50076
rect 96376 50016 96440 50020
rect 96456 50076 96520 50080
rect 96456 50020 96460 50076
rect 96460 50020 96516 50076
rect 96516 50020 96520 50076
rect 96456 50016 96520 50020
rect 96536 50076 96600 50080
rect 96536 50020 96540 50076
rect 96540 50020 96596 50076
rect 96596 50020 96600 50076
rect 96536 50016 96600 50020
rect 96616 50076 96680 50080
rect 96616 50020 96620 50076
rect 96620 50020 96676 50076
rect 96676 50020 96680 50076
rect 96616 50016 96680 50020
rect 127096 50076 127160 50080
rect 127096 50020 127100 50076
rect 127100 50020 127156 50076
rect 127156 50020 127160 50076
rect 127096 50016 127160 50020
rect 127176 50076 127240 50080
rect 127176 50020 127180 50076
rect 127180 50020 127236 50076
rect 127236 50020 127240 50076
rect 127176 50016 127240 50020
rect 127256 50076 127320 50080
rect 127256 50020 127260 50076
rect 127260 50020 127316 50076
rect 127316 50020 127320 50076
rect 127256 50016 127320 50020
rect 127336 50076 127400 50080
rect 127336 50020 127340 50076
rect 127340 50020 127396 50076
rect 127396 50020 127400 50076
rect 127336 50016 127400 50020
rect 157816 50076 157880 50080
rect 157816 50020 157820 50076
rect 157820 50020 157876 50076
rect 157876 50020 157880 50076
rect 157816 50016 157880 50020
rect 157896 50076 157960 50080
rect 157896 50020 157900 50076
rect 157900 50020 157956 50076
rect 157956 50020 157960 50076
rect 157896 50016 157960 50020
rect 157976 50076 158040 50080
rect 157976 50020 157980 50076
rect 157980 50020 158036 50076
rect 158036 50020 158040 50076
rect 157976 50016 158040 50020
rect 158056 50076 158120 50080
rect 158056 50020 158060 50076
rect 158060 50020 158116 50076
rect 158116 50020 158120 50076
rect 158056 50016 158120 50020
rect 19576 49532 19640 49536
rect 19576 49476 19580 49532
rect 19580 49476 19636 49532
rect 19636 49476 19640 49532
rect 19576 49472 19640 49476
rect 19656 49532 19720 49536
rect 19656 49476 19660 49532
rect 19660 49476 19716 49532
rect 19716 49476 19720 49532
rect 19656 49472 19720 49476
rect 19736 49532 19800 49536
rect 19736 49476 19740 49532
rect 19740 49476 19796 49532
rect 19796 49476 19800 49532
rect 19736 49472 19800 49476
rect 19816 49532 19880 49536
rect 19816 49476 19820 49532
rect 19820 49476 19876 49532
rect 19876 49476 19880 49532
rect 19816 49472 19880 49476
rect 50296 49532 50360 49536
rect 50296 49476 50300 49532
rect 50300 49476 50356 49532
rect 50356 49476 50360 49532
rect 50296 49472 50360 49476
rect 50376 49532 50440 49536
rect 50376 49476 50380 49532
rect 50380 49476 50436 49532
rect 50436 49476 50440 49532
rect 50376 49472 50440 49476
rect 50456 49532 50520 49536
rect 50456 49476 50460 49532
rect 50460 49476 50516 49532
rect 50516 49476 50520 49532
rect 50456 49472 50520 49476
rect 50536 49532 50600 49536
rect 50536 49476 50540 49532
rect 50540 49476 50596 49532
rect 50596 49476 50600 49532
rect 50536 49472 50600 49476
rect 81016 49532 81080 49536
rect 81016 49476 81020 49532
rect 81020 49476 81076 49532
rect 81076 49476 81080 49532
rect 81016 49472 81080 49476
rect 81096 49532 81160 49536
rect 81096 49476 81100 49532
rect 81100 49476 81156 49532
rect 81156 49476 81160 49532
rect 81096 49472 81160 49476
rect 81176 49532 81240 49536
rect 81176 49476 81180 49532
rect 81180 49476 81236 49532
rect 81236 49476 81240 49532
rect 81176 49472 81240 49476
rect 81256 49532 81320 49536
rect 81256 49476 81260 49532
rect 81260 49476 81316 49532
rect 81316 49476 81320 49532
rect 81256 49472 81320 49476
rect 111736 49532 111800 49536
rect 111736 49476 111740 49532
rect 111740 49476 111796 49532
rect 111796 49476 111800 49532
rect 111736 49472 111800 49476
rect 111816 49532 111880 49536
rect 111816 49476 111820 49532
rect 111820 49476 111876 49532
rect 111876 49476 111880 49532
rect 111816 49472 111880 49476
rect 111896 49532 111960 49536
rect 111896 49476 111900 49532
rect 111900 49476 111956 49532
rect 111956 49476 111960 49532
rect 111896 49472 111960 49476
rect 111976 49532 112040 49536
rect 111976 49476 111980 49532
rect 111980 49476 112036 49532
rect 112036 49476 112040 49532
rect 111976 49472 112040 49476
rect 142456 49532 142520 49536
rect 142456 49476 142460 49532
rect 142460 49476 142516 49532
rect 142516 49476 142520 49532
rect 142456 49472 142520 49476
rect 142536 49532 142600 49536
rect 142536 49476 142540 49532
rect 142540 49476 142596 49532
rect 142596 49476 142600 49532
rect 142536 49472 142600 49476
rect 142616 49532 142680 49536
rect 142616 49476 142620 49532
rect 142620 49476 142676 49532
rect 142676 49476 142680 49532
rect 142616 49472 142680 49476
rect 142696 49532 142760 49536
rect 142696 49476 142700 49532
rect 142700 49476 142756 49532
rect 142756 49476 142760 49532
rect 142696 49472 142760 49476
rect 173176 49532 173240 49536
rect 173176 49476 173180 49532
rect 173180 49476 173236 49532
rect 173236 49476 173240 49532
rect 173176 49472 173240 49476
rect 173256 49532 173320 49536
rect 173256 49476 173260 49532
rect 173260 49476 173316 49532
rect 173316 49476 173320 49532
rect 173256 49472 173320 49476
rect 173336 49532 173400 49536
rect 173336 49476 173340 49532
rect 173340 49476 173396 49532
rect 173396 49476 173400 49532
rect 173336 49472 173400 49476
rect 173416 49532 173480 49536
rect 173416 49476 173420 49532
rect 173420 49476 173476 49532
rect 173476 49476 173480 49532
rect 173416 49472 173480 49476
rect 4216 48988 4280 48992
rect 4216 48932 4220 48988
rect 4220 48932 4276 48988
rect 4276 48932 4280 48988
rect 4216 48928 4280 48932
rect 4296 48988 4360 48992
rect 4296 48932 4300 48988
rect 4300 48932 4356 48988
rect 4356 48932 4360 48988
rect 4296 48928 4360 48932
rect 4376 48988 4440 48992
rect 4376 48932 4380 48988
rect 4380 48932 4436 48988
rect 4436 48932 4440 48988
rect 4376 48928 4440 48932
rect 4456 48988 4520 48992
rect 4456 48932 4460 48988
rect 4460 48932 4516 48988
rect 4516 48932 4520 48988
rect 4456 48928 4520 48932
rect 34936 48988 35000 48992
rect 34936 48932 34940 48988
rect 34940 48932 34996 48988
rect 34996 48932 35000 48988
rect 34936 48928 35000 48932
rect 35016 48988 35080 48992
rect 35016 48932 35020 48988
rect 35020 48932 35076 48988
rect 35076 48932 35080 48988
rect 35016 48928 35080 48932
rect 35096 48988 35160 48992
rect 35096 48932 35100 48988
rect 35100 48932 35156 48988
rect 35156 48932 35160 48988
rect 35096 48928 35160 48932
rect 35176 48988 35240 48992
rect 35176 48932 35180 48988
rect 35180 48932 35236 48988
rect 35236 48932 35240 48988
rect 35176 48928 35240 48932
rect 65656 48988 65720 48992
rect 65656 48932 65660 48988
rect 65660 48932 65716 48988
rect 65716 48932 65720 48988
rect 65656 48928 65720 48932
rect 65736 48988 65800 48992
rect 65736 48932 65740 48988
rect 65740 48932 65796 48988
rect 65796 48932 65800 48988
rect 65736 48928 65800 48932
rect 65816 48988 65880 48992
rect 65816 48932 65820 48988
rect 65820 48932 65876 48988
rect 65876 48932 65880 48988
rect 65816 48928 65880 48932
rect 65896 48988 65960 48992
rect 65896 48932 65900 48988
rect 65900 48932 65956 48988
rect 65956 48932 65960 48988
rect 65896 48928 65960 48932
rect 96376 48988 96440 48992
rect 96376 48932 96380 48988
rect 96380 48932 96436 48988
rect 96436 48932 96440 48988
rect 96376 48928 96440 48932
rect 96456 48988 96520 48992
rect 96456 48932 96460 48988
rect 96460 48932 96516 48988
rect 96516 48932 96520 48988
rect 96456 48928 96520 48932
rect 96536 48988 96600 48992
rect 96536 48932 96540 48988
rect 96540 48932 96596 48988
rect 96596 48932 96600 48988
rect 96536 48928 96600 48932
rect 96616 48988 96680 48992
rect 96616 48932 96620 48988
rect 96620 48932 96676 48988
rect 96676 48932 96680 48988
rect 96616 48928 96680 48932
rect 127096 48988 127160 48992
rect 127096 48932 127100 48988
rect 127100 48932 127156 48988
rect 127156 48932 127160 48988
rect 127096 48928 127160 48932
rect 127176 48988 127240 48992
rect 127176 48932 127180 48988
rect 127180 48932 127236 48988
rect 127236 48932 127240 48988
rect 127176 48928 127240 48932
rect 127256 48988 127320 48992
rect 127256 48932 127260 48988
rect 127260 48932 127316 48988
rect 127316 48932 127320 48988
rect 127256 48928 127320 48932
rect 127336 48988 127400 48992
rect 127336 48932 127340 48988
rect 127340 48932 127396 48988
rect 127396 48932 127400 48988
rect 127336 48928 127400 48932
rect 157816 48988 157880 48992
rect 157816 48932 157820 48988
rect 157820 48932 157876 48988
rect 157876 48932 157880 48988
rect 157816 48928 157880 48932
rect 157896 48988 157960 48992
rect 157896 48932 157900 48988
rect 157900 48932 157956 48988
rect 157956 48932 157960 48988
rect 157896 48928 157960 48932
rect 157976 48988 158040 48992
rect 157976 48932 157980 48988
rect 157980 48932 158036 48988
rect 158036 48932 158040 48988
rect 157976 48928 158040 48932
rect 158056 48988 158120 48992
rect 158056 48932 158060 48988
rect 158060 48932 158116 48988
rect 158116 48932 158120 48988
rect 158056 48928 158120 48932
rect 19576 48444 19640 48448
rect 19576 48388 19580 48444
rect 19580 48388 19636 48444
rect 19636 48388 19640 48444
rect 19576 48384 19640 48388
rect 19656 48444 19720 48448
rect 19656 48388 19660 48444
rect 19660 48388 19716 48444
rect 19716 48388 19720 48444
rect 19656 48384 19720 48388
rect 19736 48444 19800 48448
rect 19736 48388 19740 48444
rect 19740 48388 19796 48444
rect 19796 48388 19800 48444
rect 19736 48384 19800 48388
rect 19816 48444 19880 48448
rect 19816 48388 19820 48444
rect 19820 48388 19876 48444
rect 19876 48388 19880 48444
rect 19816 48384 19880 48388
rect 50296 48444 50360 48448
rect 50296 48388 50300 48444
rect 50300 48388 50356 48444
rect 50356 48388 50360 48444
rect 50296 48384 50360 48388
rect 50376 48444 50440 48448
rect 50376 48388 50380 48444
rect 50380 48388 50436 48444
rect 50436 48388 50440 48444
rect 50376 48384 50440 48388
rect 50456 48444 50520 48448
rect 50456 48388 50460 48444
rect 50460 48388 50516 48444
rect 50516 48388 50520 48444
rect 50456 48384 50520 48388
rect 50536 48444 50600 48448
rect 50536 48388 50540 48444
rect 50540 48388 50596 48444
rect 50596 48388 50600 48444
rect 50536 48384 50600 48388
rect 81016 48444 81080 48448
rect 81016 48388 81020 48444
rect 81020 48388 81076 48444
rect 81076 48388 81080 48444
rect 81016 48384 81080 48388
rect 81096 48444 81160 48448
rect 81096 48388 81100 48444
rect 81100 48388 81156 48444
rect 81156 48388 81160 48444
rect 81096 48384 81160 48388
rect 81176 48444 81240 48448
rect 81176 48388 81180 48444
rect 81180 48388 81236 48444
rect 81236 48388 81240 48444
rect 81176 48384 81240 48388
rect 81256 48444 81320 48448
rect 81256 48388 81260 48444
rect 81260 48388 81316 48444
rect 81316 48388 81320 48444
rect 81256 48384 81320 48388
rect 111736 48444 111800 48448
rect 111736 48388 111740 48444
rect 111740 48388 111796 48444
rect 111796 48388 111800 48444
rect 111736 48384 111800 48388
rect 111816 48444 111880 48448
rect 111816 48388 111820 48444
rect 111820 48388 111876 48444
rect 111876 48388 111880 48444
rect 111816 48384 111880 48388
rect 111896 48444 111960 48448
rect 111896 48388 111900 48444
rect 111900 48388 111956 48444
rect 111956 48388 111960 48444
rect 111896 48384 111960 48388
rect 111976 48444 112040 48448
rect 111976 48388 111980 48444
rect 111980 48388 112036 48444
rect 112036 48388 112040 48444
rect 111976 48384 112040 48388
rect 142456 48444 142520 48448
rect 142456 48388 142460 48444
rect 142460 48388 142516 48444
rect 142516 48388 142520 48444
rect 142456 48384 142520 48388
rect 142536 48444 142600 48448
rect 142536 48388 142540 48444
rect 142540 48388 142596 48444
rect 142596 48388 142600 48444
rect 142536 48384 142600 48388
rect 142616 48444 142680 48448
rect 142616 48388 142620 48444
rect 142620 48388 142676 48444
rect 142676 48388 142680 48444
rect 142616 48384 142680 48388
rect 142696 48444 142760 48448
rect 142696 48388 142700 48444
rect 142700 48388 142756 48444
rect 142756 48388 142760 48444
rect 142696 48384 142760 48388
rect 173176 48444 173240 48448
rect 173176 48388 173180 48444
rect 173180 48388 173236 48444
rect 173236 48388 173240 48444
rect 173176 48384 173240 48388
rect 173256 48444 173320 48448
rect 173256 48388 173260 48444
rect 173260 48388 173316 48444
rect 173316 48388 173320 48444
rect 173256 48384 173320 48388
rect 173336 48444 173400 48448
rect 173336 48388 173340 48444
rect 173340 48388 173396 48444
rect 173396 48388 173400 48444
rect 173336 48384 173400 48388
rect 173416 48444 173480 48448
rect 173416 48388 173420 48444
rect 173420 48388 173476 48444
rect 173476 48388 173480 48444
rect 173416 48384 173480 48388
rect 4216 47900 4280 47904
rect 4216 47844 4220 47900
rect 4220 47844 4276 47900
rect 4276 47844 4280 47900
rect 4216 47840 4280 47844
rect 4296 47900 4360 47904
rect 4296 47844 4300 47900
rect 4300 47844 4356 47900
rect 4356 47844 4360 47900
rect 4296 47840 4360 47844
rect 4376 47900 4440 47904
rect 4376 47844 4380 47900
rect 4380 47844 4436 47900
rect 4436 47844 4440 47900
rect 4376 47840 4440 47844
rect 4456 47900 4520 47904
rect 4456 47844 4460 47900
rect 4460 47844 4516 47900
rect 4516 47844 4520 47900
rect 4456 47840 4520 47844
rect 34936 47900 35000 47904
rect 34936 47844 34940 47900
rect 34940 47844 34996 47900
rect 34996 47844 35000 47900
rect 34936 47840 35000 47844
rect 35016 47900 35080 47904
rect 35016 47844 35020 47900
rect 35020 47844 35076 47900
rect 35076 47844 35080 47900
rect 35016 47840 35080 47844
rect 35096 47900 35160 47904
rect 35096 47844 35100 47900
rect 35100 47844 35156 47900
rect 35156 47844 35160 47900
rect 35096 47840 35160 47844
rect 35176 47900 35240 47904
rect 35176 47844 35180 47900
rect 35180 47844 35236 47900
rect 35236 47844 35240 47900
rect 35176 47840 35240 47844
rect 65656 47900 65720 47904
rect 65656 47844 65660 47900
rect 65660 47844 65716 47900
rect 65716 47844 65720 47900
rect 65656 47840 65720 47844
rect 65736 47900 65800 47904
rect 65736 47844 65740 47900
rect 65740 47844 65796 47900
rect 65796 47844 65800 47900
rect 65736 47840 65800 47844
rect 65816 47900 65880 47904
rect 65816 47844 65820 47900
rect 65820 47844 65876 47900
rect 65876 47844 65880 47900
rect 65816 47840 65880 47844
rect 65896 47900 65960 47904
rect 65896 47844 65900 47900
rect 65900 47844 65956 47900
rect 65956 47844 65960 47900
rect 65896 47840 65960 47844
rect 96376 47900 96440 47904
rect 96376 47844 96380 47900
rect 96380 47844 96436 47900
rect 96436 47844 96440 47900
rect 96376 47840 96440 47844
rect 96456 47900 96520 47904
rect 96456 47844 96460 47900
rect 96460 47844 96516 47900
rect 96516 47844 96520 47900
rect 96456 47840 96520 47844
rect 96536 47900 96600 47904
rect 96536 47844 96540 47900
rect 96540 47844 96596 47900
rect 96596 47844 96600 47900
rect 96536 47840 96600 47844
rect 96616 47900 96680 47904
rect 96616 47844 96620 47900
rect 96620 47844 96676 47900
rect 96676 47844 96680 47900
rect 96616 47840 96680 47844
rect 127096 47900 127160 47904
rect 127096 47844 127100 47900
rect 127100 47844 127156 47900
rect 127156 47844 127160 47900
rect 127096 47840 127160 47844
rect 127176 47900 127240 47904
rect 127176 47844 127180 47900
rect 127180 47844 127236 47900
rect 127236 47844 127240 47900
rect 127176 47840 127240 47844
rect 127256 47900 127320 47904
rect 127256 47844 127260 47900
rect 127260 47844 127316 47900
rect 127316 47844 127320 47900
rect 127256 47840 127320 47844
rect 127336 47900 127400 47904
rect 127336 47844 127340 47900
rect 127340 47844 127396 47900
rect 127396 47844 127400 47900
rect 127336 47840 127400 47844
rect 157816 47900 157880 47904
rect 157816 47844 157820 47900
rect 157820 47844 157876 47900
rect 157876 47844 157880 47900
rect 157816 47840 157880 47844
rect 157896 47900 157960 47904
rect 157896 47844 157900 47900
rect 157900 47844 157956 47900
rect 157956 47844 157960 47900
rect 157896 47840 157960 47844
rect 157976 47900 158040 47904
rect 157976 47844 157980 47900
rect 157980 47844 158036 47900
rect 158036 47844 158040 47900
rect 157976 47840 158040 47844
rect 158056 47900 158120 47904
rect 158056 47844 158060 47900
rect 158060 47844 158116 47900
rect 158116 47844 158120 47900
rect 158056 47840 158120 47844
rect 19576 47356 19640 47360
rect 19576 47300 19580 47356
rect 19580 47300 19636 47356
rect 19636 47300 19640 47356
rect 19576 47296 19640 47300
rect 19656 47356 19720 47360
rect 19656 47300 19660 47356
rect 19660 47300 19716 47356
rect 19716 47300 19720 47356
rect 19656 47296 19720 47300
rect 19736 47356 19800 47360
rect 19736 47300 19740 47356
rect 19740 47300 19796 47356
rect 19796 47300 19800 47356
rect 19736 47296 19800 47300
rect 19816 47356 19880 47360
rect 19816 47300 19820 47356
rect 19820 47300 19876 47356
rect 19876 47300 19880 47356
rect 19816 47296 19880 47300
rect 50296 47356 50360 47360
rect 50296 47300 50300 47356
rect 50300 47300 50356 47356
rect 50356 47300 50360 47356
rect 50296 47296 50360 47300
rect 50376 47356 50440 47360
rect 50376 47300 50380 47356
rect 50380 47300 50436 47356
rect 50436 47300 50440 47356
rect 50376 47296 50440 47300
rect 50456 47356 50520 47360
rect 50456 47300 50460 47356
rect 50460 47300 50516 47356
rect 50516 47300 50520 47356
rect 50456 47296 50520 47300
rect 50536 47356 50600 47360
rect 50536 47300 50540 47356
rect 50540 47300 50596 47356
rect 50596 47300 50600 47356
rect 50536 47296 50600 47300
rect 81016 47356 81080 47360
rect 81016 47300 81020 47356
rect 81020 47300 81076 47356
rect 81076 47300 81080 47356
rect 81016 47296 81080 47300
rect 81096 47356 81160 47360
rect 81096 47300 81100 47356
rect 81100 47300 81156 47356
rect 81156 47300 81160 47356
rect 81096 47296 81160 47300
rect 81176 47356 81240 47360
rect 81176 47300 81180 47356
rect 81180 47300 81236 47356
rect 81236 47300 81240 47356
rect 81176 47296 81240 47300
rect 81256 47356 81320 47360
rect 81256 47300 81260 47356
rect 81260 47300 81316 47356
rect 81316 47300 81320 47356
rect 81256 47296 81320 47300
rect 111736 47356 111800 47360
rect 111736 47300 111740 47356
rect 111740 47300 111796 47356
rect 111796 47300 111800 47356
rect 111736 47296 111800 47300
rect 111816 47356 111880 47360
rect 111816 47300 111820 47356
rect 111820 47300 111876 47356
rect 111876 47300 111880 47356
rect 111816 47296 111880 47300
rect 111896 47356 111960 47360
rect 111896 47300 111900 47356
rect 111900 47300 111956 47356
rect 111956 47300 111960 47356
rect 111896 47296 111960 47300
rect 111976 47356 112040 47360
rect 111976 47300 111980 47356
rect 111980 47300 112036 47356
rect 112036 47300 112040 47356
rect 111976 47296 112040 47300
rect 142456 47356 142520 47360
rect 142456 47300 142460 47356
rect 142460 47300 142516 47356
rect 142516 47300 142520 47356
rect 142456 47296 142520 47300
rect 142536 47356 142600 47360
rect 142536 47300 142540 47356
rect 142540 47300 142596 47356
rect 142596 47300 142600 47356
rect 142536 47296 142600 47300
rect 142616 47356 142680 47360
rect 142616 47300 142620 47356
rect 142620 47300 142676 47356
rect 142676 47300 142680 47356
rect 142616 47296 142680 47300
rect 142696 47356 142760 47360
rect 142696 47300 142700 47356
rect 142700 47300 142756 47356
rect 142756 47300 142760 47356
rect 142696 47296 142760 47300
rect 173176 47356 173240 47360
rect 173176 47300 173180 47356
rect 173180 47300 173236 47356
rect 173236 47300 173240 47356
rect 173176 47296 173240 47300
rect 173256 47356 173320 47360
rect 173256 47300 173260 47356
rect 173260 47300 173316 47356
rect 173316 47300 173320 47356
rect 173256 47296 173320 47300
rect 173336 47356 173400 47360
rect 173336 47300 173340 47356
rect 173340 47300 173396 47356
rect 173396 47300 173400 47356
rect 173336 47296 173400 47300
rect 173416 47356 173480 47360
rect 173416 47300 173420 47356
rect 173420 47300 173476 47356
rect 173476 47300 173480 47356
rect 173416 47296 173480 47300
rect 4216 46812 4280 46816
rect 4216 46756 4220 46812
rect 4220 46756 4276 46812
rect 4276 46756 4280 46812
rect 4216 46752 4280 46756
rect 4296 46812 4360 46816
rect 4296 46756 4300 46812
rect 4300 46756 4356 46812
rect 4356 46756 4360 46812
rect 4296 46752 4360 46756
rect 4376 46812 4440 46816
rect 4376 46756 4380 46812
rect 4380 46756 4436 46812
rect 4436 46756 4440 46812
rect 4376 46752 4440 46756
rect 4456 46812 4520 46816
rect 4456 46756 4460 46812
rect 4460 46756 4516 46812
rect 4516 46756 4520 46812
rect 4456 46752 4520 46756
rect 34936 46812 35000 46816
rect 34936 46756 34940 46812
rect 34940 46756 34996 46812
rect 34996 46756 35000 46812
rect 34936 46752 35000 46756
rect 35016 46812 35080 46816
rect 35016 46756 35020 46812
rect 35020 46756 35076 46812
rect 35076 46756 35080 46812
rect 35016 46752 35080 46756
rect 35096 46812 35160 46816
rect 35096 46756 35100 46812
rect 35100 46756 35156 46812
rect 35156 46756 35160 46812
rect 35096 46752 35160 46756
rect 35176 46812 35240 46816
rect 35176 46756 35180 46812
rect 35180 46756 35236 46812
rect 35236 46756 35240 46812
rect 35176 46752 35240 46756
rect 65656 46812 65720 46816
rect 65656 46756 65660 46812
rect 65660 46756 65716 46812
rect 65716 46756 65720 46812
rect 65656 46752 65720 46756
rect 65736 46812 65800 46816
rect 65736 46756 65740 46812
rect 65740 46756 65796 46812
rect 65796 46756 65800 46812
rect 65736 46752 65800 46756
rect 65816 46812 65880 46816
rect 65816 46756 65820 46812
rect 65820 46756 65876 46812
rect 65876 46756 65880 46812
rect 65816 46752 65880 46756
rect 65896 46812 65960 46816
rect 65896 46756 65900 46812
rect 65900 46756 65956 46812
rect 65956 46756 65960 46812
rect 65896 46752 65960 46756
rect 96376 46812 96440 46816
rect 96376 46756 96380 46812
rect 96380 46756 96436 46812
rect 96436 46756 96440 46812
rect 96376 46752 96440 46756
rect 96456 46812 96520 46816
rect 96456 46756 96460 46812
rect 96460 46756 96516 46812
rect 96516 46756 96520 46812
rect 96456 46752 96520 46756
rect 96536 46812 96600 46816
rect 96536 46756 96540 46812
rect 96540 46756 96596 46812
rect 96596 46756 96600 46812
rect 96536 46752 96600 46756
rect 96616 46812 96680 46816
rect 96616 46756 96620 46812
rect 96620 46756 96676 46812
rect 96676 46756 96680 46812
rect 96616 46752 96680 46756
rect 127096 46812 127160 46816
rect 127096 46756 127100 46812
rect 127100 46756 127156 46812
rect 127156 46756 127160 46812
rect 127096 46752 127160 46756
rect 127176 46812 127240 46816
rect 127176 46756 127180 46812
rect 127180 46756 127236 46812
rect 127236 46756 127240 46812
rect 127176 46752 127240 46756
rect 127256 46812 127320 46816
rect 127256 46756 127260 46812
rect 127260 46756 127316 46812
rect 127316 46756 127320 46812
rect 127256 46752 127320 46756
rect 127336 46812 127400 46816
rect 127336 46756 127340 46812
rect 127340 46756 127396 46812
rect 127396 46756 127400 46812
rect 127336 46752 127400 46756
rect 157816 46812 157880 46816
rect 157816 46756 157820 46812
rect 157820 46756 157876 46812
rect 157876 46756 157880 46812
rect 157816 46752 157880 46756
rect 157896 46812 157960 46816
rect 157896 46756 157900 46812
rect 157900 46756 157956 46812
rect 157956 46756 157960 46812
rect 157896 46752 157960 46756
rect 157976 46812 158040 46816
rect 157976 46756 157980 46812
rect 157980 46756 158036 46812
rect 158036 46756 158040 46812
rect 157976 46752 158040 46756
rect 158056 46812 158120 46816
rect 158056 46756 158060 46812
rect 158060 46756 158116 46812
rect 158116 46756 158120 46812
rect 158056 46752 158120 46756
rect 19576 46268 19640 46272
rect 19576 46212 19580 46268
rect 19580 46212 19636 46268
rect 19636 46212 19640 46268
rect 19576 46208 19640 46212
rect 19656 46268 19720 46272
rect 19656 46212 19660 46268
rect 19660 46212 19716 46268
rect 19716 46212 19720 46268
rect 19656 46208 19720 46212
rect 19736 46268 19800 46272
rect 19736 46212 19740 46268
rect 19740 46212 19796 46268
rect 19796 46212 19800 46268
rect 19736 46208 19800 46212
rect 19816 46268 19880 46272
rect 19816 46212 19820 46268
rect 19820 46212 19876 46268
rect 19876 46212 19880 46268
rect 19816 46208 19880 46212
rect 50296 46268 50360 46272
rect 50296 46212 50300 46268
rect 50300 46212 50356 46268
rect 50356 46212 50360 46268
rect 50296 46208 50360 46212
rect 50376 46268 50440 46272
rect 50376 46212 50380 46268
rect 50380 46212 50436 46268
rect 50436 46212 50440 46268
rect 50376 46208 50440 46212
rect 50456 46268 50520 46272
rect 50456 46212 50460 46268
rect 50460 46212 50516 46268
rect 50516 46212 50520 46268
rect 50456 46208 50520 46212
rect 50536 46268 50600 46272
rect 50536 46212 50540 46268
rect 50540 46212 50596 46268
rect 50596 46212 50600 46268
rect 50536 46208 50600 46212
rect 81016 46268 81080 46272
rect 81016 46212 81020 46268
rect 81020 46212 81076 46268
rect 81076 46212 81080 46268
rect 81016 46208 81080 46212
rect 81096 46268 81160 46272
rect 81096 46212 81100 46268
rect 81100 46212 81156 46268
rect 81156 46212 81160 46268
rect 81096 46208 81160 46212
rect 81176 46268 81240 46272
rect 81176 46212 81180 46268
rect 81180 46212 81236 46268
rect 81236 46212 81240 46268
rect 81176 46208 81240 46212
rect 81256 46268 81320 46272
rect 81256 46212 81260 46268
rect 81260 46212 81316 46268
rect 81316 46212 81320 46268
rect 81256 46208 81320 46212
rect 111736 46268 111800 46272
rect 111736 46212 111740 46268
rect 111740 46212 111796 46268
rect 111796 46212 111800 46268
rect 111736 46208 111800 46212
rect 111816 46268 111880 46272
rect 111816 46212 111820 46268
rect 111820 46212 111876 46268
rect 111876 46212 111880 46268
rect 111816 46208 111880 46212
rect 111896 46268 111960 46272
rect 111896 46212 111900 46268
rect 111900 46212 111956 46268
rect 111956 46212 111960 46268
rect 111896 46208 111960 46212
rect 111976 46268 112040 46272
rect 111976 46212 111980 46268
rect 111980 46212 112036 46268
rect 112036 46212 112040 46268
rect 111976 46208 112040 46212
rect 142456 46268 142520 46272
rect 142456 46212 142460 46268
rect 142460 46212 142516 46268
rect 142516 46212 142520 46268
rect 142456 46208 142520 46212
rect 142536 46268 142600 46272
rect 142536 46212 142540 46268
rect 142540 46212 142596 46268
rect 142596 46212 142600 46268
rect 142536 46208 142600 46212
rect 142616 46268 142680 46272
rect 142616 46212 142620 46268
rect 142620 46212 142676 46268
rect 142676 46212 142680 46268
rect 142616 46208 142680 46212
rect 142696 46268 142760 46272
rect 142696 46212 142700 46268
rect 142700 46212 142756 46268
rect 142756 46212 142760 46268
rect 142696 46208 142760 46212
rect 173176 46268 173240 46272
rect 173176 46212 173180 46268
rect 173180 46212 173236 46268
rect 173236 46212 173240 46268
rect 173176 46208 173240 46212
rect 173256 46268 173320 46272
rect 173256 46212 173260 46268
rect 173260 46212 173316 46268
rect 173316 46212 173320 46268
rect 173256 46208 173320 46212
rect 173336 46268 173400 46272
rect 173336 46212 173340 46268
rect 173340 46212 173396 46268
rect 173396 46212 173400 46268
rect 173336 46208 173400 46212
rect 173416 46268 173480 46272
rect 173416 46212 173420 46268
rect 173420 46212 173476 46268
rect 173476 46212 173480 46268
rect 173416 46208 173480 46212
rect 4216 45724 4280 45728
rect 4216 45668 4220 45724
rect 4220 45668 4276 45724
rect 4276 45668 4280 45724
rect 4216 45664 4280 45668
rect 4296 45724 4360 45728
rect 4296 45668 4300 45724
rect 4300 45668 4356 45724
rect 4356 45668 4360 45724
rect 4296 45664 4360 45668
rect 4376 45724 4440 45728
rect 4376 45668 4380 45724
rect 4380 45668 4436 45724
rect 4436 45668 4440 45724
rect 4376 45664 4440 45668
rect 4456 45724 4520 45728
rect 4456 45668 4460 45724
rect 4460 45668 4516 45724
rect 4516 45668 4520 45724
rect 4456 45664 4520 45668
rect 34936 45724 35000 45728
rect 34936 45668 34940 45724
rect 34940 45668 34996 45724
rect 34996 45668 35000 45724
rect 34936 45664 35000 45668
rect 35016 45724 35080 45728
rect 35016 45668 35020 45724
rect 35020 45668 35076 45724
rect 35076 45668 35080 45724
rect 35016 45664 35080 45668
rect 35096 45724 35160 45728
rect 35096 45668 35100 45724
rect 35100 45668 35156 45724
rect 35156 45668 35160 45724
rect 35096 45664 35160 45668
rect 35176 45724 35240 45728
rect 35176 45668 35180 45724
rect 35180 45668 35236 45724
rect 35236 45668 35240 45724
rect 35176 45664 35240 45668
rect 65656 45724 65720 45728
rect 65656 45668 65660 45724
rect 65660 45668 65716 45724
rect 65716 45668 65720 45724
rect 65656 45664 65720 45668
rect 65736 45724 65800 45728
rect 65736 45668 65740 45724
rect 65740 45668 65796 45724
rect 65796 45668 65800 45724
rect 65736 45664 65800 45668
rect 65816 45724 65880 45728
rect 65816 45668 65820 45724
rect 65820 45668 65876 45724
rect 65876 45668 65880 45724
rect 65816 45664 65880 45668
rect 65896 45724 65960 45728
rect 65896 45668 65900 45724
rect 65900 45668 65956 45724
rect 65956 45668 65960 45724
rect 65896 45664 65960 45668
rect 96376 45724 96440 45728
rect 96376 45668 96380 45724
rect 96380 45668 96436 45724
rect 96436 45668 96440 45724
rect 96376 45664 96440 45668
rect 96456 45724 96520 45728
rect 96456 45668 96460 45724
rect 96460 45668 96516 45724
rect 96516 45668 96520 45724
rect 96456 45664 96520 45668
rect 96536 45724 96600 45728
rect 96536 45668 96540 45724
rect 96540 45668 96596 45724
rect 96596 45668 96600 45724
rect 96536 45664 96600 45668
rect 96616 45724 96680 45728
rect 96616 45668 96620 45724
rect 96620 45668 96676 45724
rect 96676 45668 96680 45724
rect 96616 45664 96680 45668
rect 127096 45724 127160 45728
rect 127096 45668 127100 45724
rect 127100 45668 127156 45724
rect 127156 45668 127160 45724
rect 127096 45664 127160 45668
rect 127176 45724 127240 45728
rect 127176 45668 127180 45724
rect 127180 45668 127236 45724
rect 127236 45668 127240 45724
rect 127176 45664 127240 45668
rect 127256 45724 127320 45728
rect 127256 45668 127260 45724
rect 127260 45668 127316 45724
rect 127316 45668 127320 45724
rect 127256 45664 127320 45668
rect 127336 45724 127400 45728
rect 127336 45668 127340 45724
rect 127340 45668 127396 45724
rect 127396 45668 127400 45724
rect 127336 45664 127400 45668
rect 157816 45724 157880 45728
rect 157816 45668 157820 45724
rect 157820 45668 157876 45724
rect 157876 45668 157880 45724
rect 157816 45664 157880 45668
rect 157896 45724 157960 45728
rect 157896 45668 157900 45724
rect 157900 45668 157956 45724
rect 157956 45668 157960 45724
rect 157896 45664 157960 45668
rect 157976 45724 158040 45728
rect 157976 45668 157980 45724
rect 157980 45668 158036 45724
rect 158036 45668 158040 45724
rect 157976 45664 158040 45668
rect 158056 45724 158120 45728
rect 158056 45668 158060 45724
rect 158060 45668 158116 45724
rect 158116 45668 158120 45724
rect 158056 45664 158120 45668
rect 19576 45180 19640 45184
rect 19576 45124 19580 45180
rect 19580 45124 19636 45180
rect 19636 45124 19640 45180
rect 19576 45120 19640 45124
rect 19656 45180 19720 45184
rect 19656 45124 19660 45180
rect 19660 45124 19716 45180
rect 19716 45124 19720 45180
rect 19656 45120 19720 45124
rect 19736 45180 19800 45184
rect 19736 45124 19740 45180
rect 19740 45124 19796 45180
rect 19796 45124 19800 45180
rect 19736 45120 19800 45124
rect 19816 45180 19880 45184
rect 19816 45124 19820 45180
rect 19820 45124 19876 45180
rect 19876 45124 19880 45180
rect 19816 45120 19880 45124
rect 50296 45180 50360 45184
rect 50296 45124 50300 45180
rect 50300 45124 50356 45180
rect 50356 45124 50360 45180
rect 50296 45120 50360 45124
rect 50376 45180 50440 45184
rect 50376 45124 50380 45180
rect 50380 45124 50436 45180
rect 50436 45124 50440 45180
rect 50376 45120 50440 45124
rect 50456 45180 50520 45184
rect 50456 45124 50460 45180
rect 50460 45124 50516 45180
rect 50516 45124 50520 45180
rect 50456 45120 50520 45124
rect 50536 45180 50600 45184
rect 50536 45124 50540 45180
rect 50540 45124 50596 45180
rect 50596 45124 50600 45180
rect 50536 45120 50600 45124
rect 81016 45180 81080 45184
rect 81016 45124 81020 45180
rect 81020 45124 81076 45180
rect 81076 45124 81080 45180
rect 81016 45120 81080 45124
rect 81096 45180 81160 45184
rect 81096 45124 81100 45180
rect 81100 45124 81156 45180
rect 81156 45124 81160 45180
rect 81096 45120 81160 45124
rect 81176 45180 81240 45184
rect 81176 45124 81180 45180
rect 81180 45124 81236 45180
rect 81236 45124 81240 45180
rect 81176 45120 81240 45124
rect 81256 45180 81320 45184
rect 81256 45124 81260 45180
rect 81260 45124 81316 45180
rect 81316 45124 81320 45180
rect 81256 45120 81320 45124
rect 111736 45180 111800 45184
rect 111736 45124 111740 45180
rect 111740 45124 111796 45180
rect 111796 45124 111800 45180
rect 111736 45120 111800 45124
rect 111816 45180 111880 45184
rect 111816 45124 111820 45180
rect 111820 45124 111876 45180
rect 111876 45124 111880 45180
rect 111816 45120 111880 45124
rect 111896 45180 111960 45184
rect 111896 45124 111900 45180
rect 111900 45124 111956 45180
rect 111956 45124 111960 45180
rect 111896 45120 111960 45124
rect 111976 45180 112040 45184
rect 111976 45124 111980 45180
rect 111980 45124 112036 45180
rect 112036 45124 112040 45180
rect 111976 45120 112040 45124
rect 142456 45180 142520 45184
rect 142456 45124 142460 45180
rect 142460 45124 142516 45180
rect 142516 45124 142520 45180
rect 142456 45120 142520 45124
rect 142536 45180 142600 45184
rect 142536 45124 142540 45180
rect 142540 45124 142596 45180
rect 142596 45124 142600 45180
rect 142536 45120 142600 45124
rect 142616 45180 142680 45184
rect 142616 45124 142620 45180
rect 142620 45124 142676 45180
rect 142676 45124 142680 45180
rect 142616 45120 142680 45124
rect 142696 45180 142760 45184
rect 142696 45124 142700 45180
rect 142700 45124 142756 45180
rect 142756 45124 142760 45180
rect 142696 45120 142760 45124
rect 173176 45180 173240 45184
rect 173176 45124 173180 45180
rect 173180 45124 173236 45180
rect 173236 45124 173240 45180
rect 173176 45120 173240 45124
rect 173256 45180 173320 45184
rect 173256 45124 173260 45180
rect 173260 45124 173316 45180
rect 173316 45124 173320 45180
rect 173256 45120 173320 45124
rect 173336 45180 173400 45184
rect 173336 45124 173340 45180
rect 173340 45124 173396 45180
rect 173396 45124 173400 45180
rect 173336 45120 173400 45124
rect 173416 45180 173480 45184
rect 173416 45124 173420 45180
rect 173420 45124 173476 45180
rect 173476 45124 173480 45180
rect 173416 45120 173480 45124
rect 4216 44636 4280 44640
rect 4216 44580 4220 44636
rect 4220 44580 4276 44636
rect 4276 44580 4280 44636
rect 4216 44576 4280 44580
rect 4296 44636 4360 44640
rect 4296 44580 4300 44636
rect 4300 44580 4356 44636
rect 4356 44580 4360 44636
rect 4296 44576 4360 44580
rect 4376 44636 4440 44640
rect 4376 44580 4380 44636
rect 4380 44580 4436 44636
rect 4436 44580 4440 44636
rect 4376 44576 4440 44580
rect 4456 44636 4520 44640
rect 4456 44580 4460 44636
rect 4460 44580 4516 44636
rect 4516 44580 4520 44636
rect 4456 44576 4520 44580
rect 34936 44636 35000 44640
rect 34936 44580 34940 44636
rect 34940 44580 34996 44636
rect 34996 44580 35000 44636
rect 34936 44576 35000 44580
rect 35016 44636 35080 44640
rect 35016 44580 35020 44636
rect 35020 44580 35076 44636
rect 35076 44580 35080 44636
rect 35016 44576 35080 44580
rect 35096 44636 35160 44640
rect 35096 44580 35100 44636
rect 35100 44580 35156 44636
rect 35156 44580 35160 44636
rect 35096 44576 35160 44580
rect 35176 44636 35240 44640
rect 35176 44580 35180 44636
rect 35180 44580 35236 44636
rect 35236 44580 35240 44636
rect 35176 44576 35240 44580
rect 65656 44636 65720 44640
rect 65656 44580 65660 44636
rect 65660 44580 65716 44636
rect 65716 44580 65720 44636
rect 65656 44576 65720 44580
rect 65736 44636 65800 44640
rect 65736 44580 65740 44636
rect 65740 44580 65796 44636
rect 65796 44580 65800 44636
rect 65736 44576 65800 44580
rect 65816 44636 65880 44640
rect 65816 44580 65820 44636
rect 65820 44580 65876 44636
rect 65876 44580 65880 44636
rect 65816 44576 65880 44580
rect 65896 44636 65960 44640
rect 65896 44580 65900 44636
rect 65900 44580 65956 44636
rect 65956 44580 65960 44636
rect 65896 44576 65960 44580
rect 96376 44636 96440 44640
rect 96376 44580 96380 44636
rect 96380 44580 96436 44636
rect 96436 44580 96440 44636
rect 96376 44576 96440 44580
rect 96456 44636 96520 44640
rect 96456 44580 96460 44636
rect 96460 44580 96516 44636
rect 96516 44580 96520 44636
rect 96456 44576 96520 44580
rect 96536 44636 96600 44640
rect 96536 44580 96540 44636
rect 96540 44580 96596 44636
rect 96596 44580 96600 44636
rect 96536 44576 96600 44580
rect 96616 44636 96680 44640
rect 96616 44580 96620 44636
rect 96620 44580 96676 44636
rect 96676 44580 96680 44636
rect 96616 44576 96680 44580
rect 127096 44636 127160 44640
rect 127096 44580 127100 44636
rect 127100 44580 127156 44636
rect 127156 44580 127160 44636
rect 127096 44576 127160 44580
rect 127176 44636 127240 44640
rect 127176 44580 127180 44636
rect 127180 44580 127236 44636
rect 127236 44580 127240 44636
rect 127176 44576 127240 44580
rect 127256 44636 127320 44640
rect 127256 44580 127260 44636
rect 127260 44580 127316 44636
rect 127316 44580 127320 44636
rect 127256 44576 127320 44580
rect 127336 44636 127400 44640
rect 127336 44580 127340 44636
rect 127340 44580 127396 44636
rect 127396 44580 127400 44636
rect 127336 44576 127400 44580
rect 157816 44636 157880 44640
rect 157816 44580 157820 44636
rect 157820 44580 157876 44636
rect 157876 44580 157880 44636
rect 157816 44576 157880 44580
rect 157896 44636 157960 44640
rect 157896 44580 157900 44636
rect 157900 44580 157956 44636
rect 157956 44580 157960 44636
rect 157896 44576 157960 44580
rect 157976 44636 158040 44640
rect 157976 44580 157980 44636
rect 157980 44580 158036 44636
rect 158036 44580 158040 44636
rect 157976 44576 158040 44580
rect 158056 44636 158120 44640
rect 158056 44580 158060 44636
rect 158060 44580 158116 44636
rect 158116 44580 158120 44636
rect 158056 44576 158120 44580
rect 19576 44092 19640 44096
rect 19576 44036 19580 44092
rect 19580 44036 19636 44092
rect 19636 44036 19640 44092
rect 19576 44032 19640 44036
rect 19656 44092 19720 44096
rect 19656 44036 19660 44092
rect 19660 44036 19716 44092
rect 19716 44036 19720 44092
rect 19656 44032 19720 44036
rect 19736 44092 19800 44096
rect 19736 44036 19740 44092
rect 19740 44036 19796 44092
rect 19796 44036 19800 44092
rect 19736 44032 19800 44036
rect 19816 44092 19880 44096
rect 19816 44036 19820 44092
rect 19820 44036 19876 44092
rect 19876 44036 19880 44092
rect 19816 44032 19880 44036
rect 50296 44092 50360 44096
rect 50296 44036 50300 44092
rect 50300 44036 50356 44092
rect 50356 44036 50360 44092
rect 50296 44032 50360 44036
rect 50376 44092 50440 44096
rect 50376 44036 50380 44092
rect 50380 44036 50436 44092
rect 50436 44036 50440 44092
rect 50376 44032 50440 44036
rect 50456 44092 50520 44096
rect 50456 44036 50460 44092
rect 50460 44036 50516 44092
rect 50516 44036 50520 44092
rect 50456 44032 50520 44036
rect 50536 44092 50600 44096
rect 50536 44036 50540 44092
rect 50540 44036 50596 44092
rect 50596 44036 50600 44092
rect 50536 44032 50600 44036
rect 81016 44092 81080 44096
rect 81016 44036 81020 44092
rect 81020 44036 81076 44092
rect 81076 44036 81080 44092
rect 81016 44032 81080 44036
rect 81096 44092 81160 44096
rect 81096 44036 81100 44092
rect 81100 44036 81156 44092
rect 81156 44036 81160 44092
rect 81096 44032 81160 44036
rect 81176 44092 81240 44096
rect 81176 44036 81180 44092
rect 81180 44036 81236 44092
rect 81236 44036 81240 44092
rect 81176 44032 81240 44036
rect 81256 44092 81320 44096
rect 81256 44036 81260 44092
rect 81260 44036 81316 44092
rect 81316 44036 81320 44092
rect 81256 44032 81320 44036
rect 111736 44092 111800 44096
rect 111736 44036 111740 44092
rect 111740 44036 111796 44092
rect 111796 44036 111800 44092
rect 111736 44032 111800 44036
rect 111816 44092 111880 44096
rect 111816 44036 111820 44092
rect 111820 44036 111876 44092
rect 111876 44036 111880 44092
rect 111816 44032 111880 44036
rect 111896 44092 111960 44096
rect 111896 44036 111900 44092
rect 111900 44036 111956 44092
rect 111956 44036 111960 44092
rect 111896 44032 111960 44036
rect 111976 44092 112040 44096
rect 111976 44036 111980 44092
rect 111980 44036 112036 44092
rect 112036 44036 112040 44092
rect 111976 44032 112040 44036
rect 142456 44092 142520 44096
rect 142456 44036 142460 44092
rect 142460 44036 142516 44092
rect 142516 44036 142520 44092
rect 142456 44032 142520 44036
rect 142536 44092 142600 44096
rect 142536 44036 142540 44092
rect 142540 44036 142596 44092
rect 142596 44036 142600 44092
rect 142536 44032 142600 44036
rect 142616 44092 142680 44096
rect 142616 44036 142620 44092
rect 142620 44036 142676 44092
rect 142676 44036 142680 44092
rect 142616 44032 142680 44036
rect 142696 44092 142760 44096
rect 142696 44036 142700 44092
rect 142700 44036 142756 44092
rect 142756 44036 142760 44092
rect 142696 44032 142760 44036
rect 173176 44092 173240 44096
rect 173176 44036 173180 44092
rect 173180 44036 173236 44092
rect 173236 44036 173240 44092
rect 173176 44032 173240 44036
rect 173256 44092 173320 44096
rect 173256 44036 173260 44092
rect 173260 44036 173316 44092
rect 173316 44036 173320 44092
rect 173256 44032 173320 44036
rect 173336 44092 173400 44096
rect 173336 44036 173340 44092
rect 173340 44036 173396 44092
rect 173396 44036 173400 44092
rect 173336 44032 173400 44036
rect 173416 44092 173480 44096
rect 173416 44036 173420 44092
rect 173420 44036 173476 44092
rect 173476 44036 173480 44092
rect 173416 44032 173480 44036
rect 4216 43548 4280 43552
rect 4216 43492 4220 43548
rect 4220 43492 4276 43548
rect 4276 43492 4280 43548
rect 4216 43488 4280 43492
rect 4296 43548 4360 43552
rect 4296 43492 4300 43548
rect 4300 43492 4356 43548
rect 4356 43492 4360 43548
rect 4296 43488 4360 43492
rect 4376 43548 4440 43552
rect 4376 43492 4380 43548
rect 4380 43492 4436 43548
rect 4436 43492 4440 43548
rect 4376 43488 4440 43492
rect 4456 43548 4520 43552
rect 4456 43492 4460 43548
rect 4460 43492 4516 43548
rect 4516 43492 4520 43548
rect 4456 43488 4520 43492
rect 34936 43548 35000 43552
rect 34936 43492 34940 43548
rect 34940 43492 34996 43548
rect 34996 43492 35000 43548
rect 34936 43488 35000 43492
rect 35016 43548 35080 43552
rect 35016 43492 35020 43548
rect 35020 43492 35076 43548
rect 35076 43492 35080 43548
rect 35016 43488 35080 43492
rect 35096 43548 35160 43552
rect 35096 43492 35100 43548
rect 35100 43492 35156 43548
rect 35156 43492 35160 43548
rect 35096 43488 35160 43492
rect 35176 43548 35240 43552
rect 35176 43492 35180 43548
rect 35180 43492 35236 43548
rect 35236 43492 35240 43548
rect 35176 43488 35240 43492
rect 65656 43548 65720 43552
rect 65656 43492 65660 43548
rect 65660 43492 65716 43548
rect 65716 43492 65720 43548
rect 65656 43488 65720 43492
rect 65736 43548 65800 43552
rect 65736 43492 65740 43548
rect 65740 43492 65796 43548
rect 65796 43492 65800 43548
rect 65736 43488 65800 43492
rect 65816 43548 65880 43552
rect 65816 43492 65820 43548
rect 65820 43492 65876 43548
rect 65876 43492 65880 43548
rect 65816 43488 65880 43492
rect 65896 43548 65960 43552
rect 65896 43492 65900 43548
rect 65900 43492 65956 43548
rect 65956 43492 65960 43548
rect 65896 43488 65960 43492
rect 96376 43548 96440 43552
rect 96376 43492 96380 43548
rect 96380 43492 96436 43548
rect 96436 43492 96440 43548
rect 96376 43488 96440 43492
rect 96456 43548 96520 43552
rect 96456 43492 96460 43548
rect 96460 43492 96516 43548
rect 96516 43492 96520 43548
rect 96456 43488 96520 43492
rect 96536 43548 96600 43552
rect 96536 43492 96540 43548
rect 96540 43492 96596 43548
rect 96596 43492 96600 43548
rect 96536 43488 96600 43492
rect 96616 43548 96680 43552
rect 96616 43492 96620 43548
rect 96620 43492 96676 43548
rect 96676 43492 96680 43548
rect 96616 43488 96680 43492
rect 127096 43548 127160 43552
rect 127096 43492 127100 43548
rect 127100 43492 127156 43548
rect 127156 43492 127160 43548
rect 127096 43488 127160 43492
rect 127176 43548 127240 43552
rect 127176 43492 127180 43548
rect 127180 43492 127236 43548
rect 127236 43492 127240 43548
rect 127176 43488 127240 43492
rect 127256 43548 127320 43552
rect 127256 43492 127260 43548
rect 127260 43492 127316 43548
rect 127316 43492 127320 43548
rect 127256 43488 127320 43492
rect 127336 43548 127400 43552
rect 127336 43492 127340 43548
rect 127340 43492 127396 43548
rect 127396 43492 127400 43548
rect 127336 43488 127400 43492
rect 157816 43548 157880 43552
rect 157816 43492 157820 43548
rect 157820 43492 157876 43548
rect 157876 43492 157880 43548
rect 157816 43488 157880 43492
rect 157896 43548 157960 43552
rect 157896 43492 157900 43548
rect 157900 43492 157956 43548
rect 157956 43492 157960 43548
rect 157896 43488 157960 43492
rect 157976 43548 158040 43552
rect 157976 43492 157980 43548
rect 157980 43492 158036 43548
rect 158036 43492 158040 43548
rect 157976 43488 158040 43492
rect 158056 43548 158120 43552
rect 158056 43492 158060 43548
rect 158060 43492 158116 43548
rect 158116 43492 158120 43548
rect 158056 43488 158120 43492
rect 19576 43004 19640 43008
rect 19576 42948 19580 43004
rect 19580 42948 19636 43004
rect 19636 42948 19640 43004
rect 19576 42944 19640 42948
rect 19656 43004 19720 43008
rect 19656 42948 19660 43004
rect 19660 42948 19716 43004
rect 19716 42948 19720 43004
rect 19656 42944 19720 42948
rect 19736 43004 19800 43008
rect 19736 42948 19740 43004
rect 19740 42948 19796 43004
rect 19796 42948 19800 43004
rect 19736 42944 19800 42948
rect 19816 43004 19880 43008
rect 19816 42948 19820 43004
rect 19820 42948 19876 43004
rect 19876 42948 19880 43004
rect 19816 42944 19880 42948
rect 50296 43004 50360 43008
rect 50296 42948 50300 43004
rect 50300 42948 50356 43004
rect 50356 42948 50360 43004
rect 50296 42944 50360 42948
rect 50376 43004 50440 43008
rect 50376 42948 50380 43004
rect 50380 42948 50436 43004
rect 50436 42948 50440 43004
rect 50376 42944 50440 42948
rect 50456 43004 50520 43008
rect 50456 42948 50460 43004
rect 50460 42948 50516 43004
rect 50516 42948 50520 43004
rect 50456 42944 50520 42948
rect 50536 43004 50600 43008
rect 50536 42948 50540 43004
rect 50540 42948 50596 43004
rect 50596 42948 50600 43004
rect 50536 42944 50600 42948
rect 81016 43004 81080 43008
rect 81016 42948 81020 43004
rect 81020 42948 81076 43004
rect 81076 42948 81080 43004
rect 81016 42944 81080 42948
rect 81096 43004 81160 43008
rect 81096 42948 81100 43004
rect 81100 42948 81156 43004
rect 81156 42948 81160 43004
rect 81096 42944 81160 42948
rect 81176 43004 81240 43008
rect 81176 42948 81180 43004
rect 81180 42948 81236 43004
rect 81236 42948 81240 43004
rect 81176 42944 81240 42948
rect 81256 43004 81320 43008
rect 81256 42948 81260 43004
rect 81260 42948 81316 43004
rect 81316 42948 81320 43004
rect 81256 42944 81320 42948
rect 111736 43004 111800 43008
rect 111736 42948 111740 43004
rect 111740 42948 111796 43004
rect 111796 42948 111800 43004
rect 111736 42944 111800 42948
rect 111816 43004 111880 43008
rect 111816 42948 111820 43004
rect 111820 42948 111876 43004
rect 111876 42948 111880 43004
rect 111816 42944 111880 42948
rect 111896 43004 111960 43008
rect 111896 42948 111900 43004
rect 111900 42948 111956 43004
rect 111956 42948 111960 43004
rect 111896 42944 111960 42948
rect 111976 43004 112040 43008
rect 111976 42948 111980 43004
rect 111980 42948 112036 43004
rect 112036 42948 112040 43004
rect 111976 42944 112040 42948
rect 142456 43004 142520 43008
rect 142456 42948 142460 43004
rect 142460 42948 142516 43004
rect 142516 42948 142520 43004
rect 142456 42944 142520 42948
rect 142536 43004 142600 43008
rect 142536 42948 142540 43004
rect 142540 42948 142596 43004
rect 142596 42948 142600 43004
rect 142536 42944 142600 42948
rect 142616 43004 142680 43008
rect 142616 42948 142620 43004
rect 142620 42948 142676 43004
rect 142676 42948 142680 43004
rect 142616 42944 142680 42948
rect 142696 43004 142760 43008
rect 142696 42948 142700 43004
rect 142700 42948 142756 43004
rect 142756 42948 142760 43004
rect 142696 42944 142760 42948
rect 173176 43004 173240 43008
rect 173176 42948 173180 43004
rect 173180 42948 173236 43004
rect 173236 42948 173240 43004
rect 173176 42944 173240 42948
rect 173256 43004 173320 43008
rect 173256 42948 173260 43004
rect 173260 42948 173316 43004
rect 173316 42948 173320 43004
rect 173256 42944 173320 42948
rect 173336 43004 173400 43008
rect 173336 42948 173340 43004
rect 173340 42948 173396 43004
rect 173396 42948 173400 43004
rect 173336 42944 173400 42948
rect 173416 43004 173480 43008
rect 173416 42948 173420 43004
rect 173420 42948 173476 43004
rect 173476 42948 173480 43004
rect 173416 42944 173480 42948
rect 4216 42460 4280 42464
rect 4216 42404 4220 42460
rect 4220 42404 4276 42460
rect 4276 42404 4280 42460
rect 4216 42400 4280 42404
rect 4296 42460 4360 42464
rect 4296 42404 4300 42460
rect 4300 42404 4356 42460
rect 4356 42404 4360 42460
rect 4296 42400 4360 42404
rect 4376 42460 4440 42464
rect 4376 42404 4380 42460
rect 4380 42404 4436 42460
rect 4436 42404 4440 42460
rect 4376 42400 4440 42404
rect 4456 42460 4520 42464
rect 4456 42404 4460 42460
rect 4460 42404 4516 42460
rect 4516 42404 4520 42460
rect 4456 42400 4520 42404
rect 34936 42460 35000 42464
rect 34936 42404 34940 42460
rect 34940 42404 34996 42460
rect 34996 42404 35000 42460
rect 34936 42400 35000 42404
rect 35016 42460 35080 42464
rect 35016 42404 35020 42460
rect 35020 42404 35076 42460
rect 35076 42404 35080 42460
rect 35016 42400 35080 42404
rect 35096 42460 35160 42464
rect 35096 42404 35100 42460
rect 35100 42404 35156 42460
rect 35156 42404 35160 42460
rect 35096 42400 35160 42404
rect 35176 42460 35240 42464
rect 35176 42404 35180 42460
rect 35180 42404 35236 42460
rect 35236 42404 35240 42460
rect 35176 42400 35240 42404
rect 65656 42460 65720 42464
rect 65656 42404 65660 42460
rect 65660 42404 65716 42460
rect 65716 42404 65720 42460
rect 65656 42400 65720 42404
rect 65736 42460 65800 42464
rect 65736 42404 65740 42460
rect 65740 42404 65796 42460
rect 65796 42404 65800 42460
rect 65736 42400 65800 42404
rect 65816 42460 65880 42464
rect 65816 42404 65820 42460
rect 65820 42404 65876 42460
rect 65876 42404 65880 42460
rect 65816 42400 65880 42404
rect 65896 42460 65960 42464
rect 65896 42404 65900 42460
rect 65900 42404 65956 42460
rect 65956 42404 65960 42460
rect 65896 42400 65960 42404
rect 96376 42460 96440 42464
rect 96376 42404 96380 42460
rect 96380 42404 96436 42460
rect 96436 42404 96440 42460
rect 96376 42400 96440 42404
rect 96456 42460 96520 42464
rect 96456 42404 96460 42460
rect 96460 42404 96516 42460
rect 96516 42404 96520 42460
rect 96456 42400 96520 42404
rect 96536 42460 96600 42464
rect 96536 42404 96540 42460
rect 96540 42404 96596 42460
rect 96596 42404 96600 42460
rect 96536 42400 96600 42404
rect 96616 42460 96680 42464
rect 96616 42404 96620 42460
rect 96620 42404 96676 42460
rect 96676 42404 96680 42460
rect 96616 42400 96680 42404
rect 127096 42460 127160 42464
rect 127096 42404 127100 42460
rect 127100 42404 127156 42460
rect 127156 42404 127160 42460
rect 127096 42400 127160 42404
rect 127176 42460 127240 42464
rect 127176 42404 127180 42460
rect 127180 42404 127236 42460
rect 127236 42404 127240 42460
rect 127176 42400 127240 42404
rect 127256 42460 127320 42464
rect 127256 42404 127260 42460
rect 127260 42404 127316 42460
rect 127316 42404 127320 42460
rect 127256 42400 127320 42404
rect 127336 42460 127400 42464
rect 127336 42404 127340 42460
rect 127340 42404 127396 42460
rect 127396 42404 127400 42460
rect 127336 42400 127400 42404
rect 157816 42460 157880 42464
rect 157816 42404 157820 42460
rect 157820 42404 157876 42460
rect 157876 42404 157880 42460
rect 157816 42400 157880 42404
rect 157896 42460 157960 42464
rect 157896 42404 157900 42460
rect 157900 42404 157956 42460
rect 157956 42404 157960 42460
rect 157896 42400 157960 42404
rect 157976 42460 158040 42464
rect 157976 42404 157980 42460
rect 157980 42404 158036 42460
rect 158036 42404 158040 42460
rect 157976 42400 158040 42404
rect 158056 42460 158120 42464
rect 158056 42404 158060 42460
rect 158060 42404 158116 42460
rect 158116 42404 158120 42460
rect 158056 42400 158120 42404
rect 19576 41916 19640 41920
rect 19576 41860 19580 41916
rect 19580 41860 19636 41916
rect 19636 41860 19640 41916
rect 19576 41856 19640 41860
rect 19656 41916 19720 41920
rect 19656 41860 19660 41916
rect 19660 41860 19716 41916
rect 19716 41860 19720 41916
rect 19656 41856 19720 41860
rect 19736 41916 19800 41920
rect 19736 41860 19740 41916
rect 19740 41860 19796 41916
rect 19796 41860 19800 41916
rect 19736 41856 19800 41860
rect 19816 41916 19880 41920
rect 19816 41860 19820 41916
rect 19820 41860 19876 41916
rect 19876 41860 19880 41916
rect 19816 41856 19880 41860
rect 50296 41916 50360 41920
rect 50296 41860 50300 41916
rect 50300 41860 50356 41916
rect 50356 41860 50360 41916
rect 50296 41856 50360 41860
rect 50376 41916 50440 41920
rect 50376 41860 50380 41916
rect 50380 41860 50436 41916
rect 50436 41860 50440 41916
rect 50376 41856 50440 41860
rect 50456 41916 50520 41920
rect 50456 41860 50460 41916
rect 50460 41860 50516 41916
rect 50516 41860 50520 41916
rect 50456 41856 50520 41860
rect 50536 41916 50600 41920
rect 50536 41860 50540 41916
rect 50540 41860 50596 41916
rect 50596 41860 50600 41916
rect 50536 41856 50600 41860
rect 81016 41916 81080 41920
rect 81016 41860 81020 41916
rect 81020 41860 81076 41916
rect 81076 41860 81080 41916
rect 81016 41856 81080 41860
rect 81096 41916 81160 41920
rect 81096 41860 81100 41916
rect 81100 41860 81156 41916
rect 81156 41860 81160 41916
rect 81096 41856 81160 41860
rect 81176 41916 81240 41920
rect 81176 41860 81180 41916
rect 81180 41860 81236 41916
rect 81236 41860 81240 41916
rect 81176 41856 81240 41860
rect 81256 41916 81320 41920
rect 81256 41860 81260 41916
rect 81260 41860 81316 41916
rect 81316 41860 81320 41916
rect 81256 41856 81320 41860
rect 111736 41916 111800 41920
rect 111736 41860 111740 41916
rect 111740 41860 111796 41916
rect 111796 41860 111800 41916
rect 111736 41856 111800 41860
rect 111816 41916 111880 41920
rect 111816 41860 111820 41916
rect 111820 41860 111876 41916
rect 111876 41860 111880 41916
rect 111816 41856 111880 41860
rect 111896 41916 111960 41920
rect 111896 41860 111900 41916
rect 111900 41860 111956 41916
rect 111956 41860 111960 41916
rect 111896 41856 111960 41860
rect 111976 41916 112040 41920
rect 111976 41860 111980 41916
rect 111980 41860 112036 41916
rect 112036 41860 112040 41916
rect 111976 41856 112040 41860
rect 142456 41916 142520 41920
rect 142456 41860 142460 41916
rect 142460 41860 142516 41916
rect 142516 41860 142520 41916
rect 142456 41856 142520 41860
rect 142536 41916 142600 41920
rect 142536 41860 142540 41916
rect 142540 41860 142596 41916
rect 142596 41860 142600 41916
rect 142536 41856 142600 41860
rect 142616 41916 142680 41920
rect 142616 41860 142620 41916
rect 142620 41860 142676 41916
rect 142676 41860 142680 41916
rect 142616 41856 142680 41860
rect 142696 41916 142760 41920
rect 142696 41860 142700 41916
rect 142700 41860 142756 41916
rect 142756 41860 142760 41916
rect 142696 41856 142760 41860
rect 173176 41916 173240 41920
rect 173176 41860 173180 41916
rect 173180 41860 173236 41916
rect 173236 41860 173240 41916
rect 173176 41856 173240 41860
rect 173256 41916 173320 41920
rect 173256 41860 173260 41916
rect 173260 41860 173316 41916
rect 173316 41860 173320 41916
rect 173256 41856 173320 41860
rect 173336 41916 173400 41920
rect 173336 41860 173340 41916
rect 173340 41860 173396 41916
rect 173396 41860 173400 41916
rect 173336 41856 173400 41860
rect 173416 41916 173480 41920
rect 173416 41860 173420 41916
rect 173420 41860 173476 41916
rect 173476 41860 173480 41916
rect 173416 41856 173480 41860
rect 4216 41372 4280 41376
rect 4216 41316 4220 41372
rect 4220 41316 4276 41372
rect 4276 41316 4280 41372
rect 4216 41312 4280 41316
rect 4296 41372 4360 41376
rect 4296 41316 4300 41372
rect 4300 41316 4356 41372
rect 4356 41316 4360 41372
rect 4296 41312 4360 41316
rect 4376 41372 4440 41376
rect 4376 41316 4380 41372
rect 4380 41316 4436 41372
rect 4436 41316 4440 41372
rect 4376 41312 4440 41316
rect 4456 41372 4520 41376
rect 4456 41316 4460 41372
rect 4460 41316 4516 41372
rect 4516 41316 4520 41372
rect 4456 41312 4520 41316
rect 34936 41372 35000 41376
rect 34936 41316 34940 41372
rect 34940 41316 34996 41372
rect 34996 41316 35000 41372
rect 34936 41312 35000 41316
rect 35016 41372 35080 41376
rect 35016 41316 35020 41372
rect 35020 41316 35076 41372
rect 35076 41316 35080 41372
rect 35016 41312 35080 41316
rect 35096 41372 35160 41376
rect 35096 41316 35100 41372
rect 35100 41316 35156 41372
rect 35156 41316 35160 41372
rect 35096 41312 35160 41316
rect 35176 41372 35240 41376
rect 35176 41316 35180 41372
rect 35180 41316 35236 41372
rect 35236 41316 35240 41372
rect 35176 41312 35240 41316
rect 65656 41372 65720 41376
rect 65656 41316 65660 41372
rect 65660 41316 65716 41372
rect 65716 41316 65720 41372
rect 65656 41312 65720 41316
rect 65736 41372 65800 41376
rect 65736 41316 65740 41372
rect 65740 41316 65796 41372
rect 65796 41316 65800 41372
rect 65736 41312 65800 41316
rect 65816 41372 65880 41376
rect 65816 41316 65820 41372
rect 65820 41316 65876 41372
rect 65876 41316 65880 41372
rect 65816 41312 65880 41316
rect 65896 41372 65960 41376
rect 65896 41316 65900 41372
rect 65900 41316 65956 41372
rect 65956 41316 65960 41372
rect 65896 41312 65960 41316
rect 96376 41372 96440 41376
rect 96376 41316 96380 41372
rect 96380 41316 96436 41372
rect 96436 41316 96440 41372
rect 96376 41312 96440 41316
rect 96456 41372 96520 41376
rect 96456 41316 96460 41372
rect 96460 41316 96516 41372
rect 96516 41316 96520 41372
rect 96456 41312 96520 41316
rect 96536 41372 96600 41376
rect 96536 41316 96540 41372
rect 96540 41316 96596 41372
rect 96596 41316 96600 41372
rect 96536 41312 96600 41316
rect 96616 41372 96680 41376
rect 96616 41316 96620 41372
rect 96620 41316 96676 41372
rect 96676 41316 96680 41372
rect 96616 41312 96680 41316
rect 127096 41372 127160 41376
rect 127096 41316 127100 41372
rect 127100 41316 127156 41372
rect 127156 41316 127160 41372
rect 127096 41312 127160 41316
rect 127176 41372 127240 41376
rect 127176 41316 127180 41372
rect 127180 41316 127236 41372
rect 127236 41316 127240 41372
rect 127176 41312 127240 41316
rect 127256 41372 127320 41376
rect 127256 41316 127260 41372
rect 127260 41316 127316 41372
rect 127316 41316 127320 41372
rect 127256 41312 127320 41316
rect 127336 41372 127400 41376
rect 127336 41316 127340 41372
rect 127340 41316 127396 41372
rect 127396 41316 127400 41372
rect 127336 41312 127400 41316
rect 157816 41372 157880 41376
rect 157816 41316 157820 41372
rect 157820 41316 157876 41372
rect 157876 41316 157880 41372
rect 157816 41312 157880 41316
rect 157896 41372 157960 41376
rect 157896 41316 157900 41372
rect 157900 41316 157956 41372
rect 157956 41316 157960 41372
rect 157896 41312 157960 41316
rect 157976 41372 158040 41376
rect 157976 41316 157980 41372
rect 157980 41316 158036 41372
rect 158036 41316 158040 41372
rect 157976 41312 158040 41316
rect 158056 41372 158120 41376
rect 158056 41316 158060 41372
rect 158060 41316 158116 41372
rect 158116 41316 158120 41372
rect 158056 41312 158120 41316
rect 19576 40828 19640 40832
rect 19576 40772 19580 40828
rect 19580 40772 19636 40828
rect 19636 40772 19640 40828
rect 19576 40768 19640 40772
rect 19656 40828 19720 40832
rect 19656 40772 19660 40828
rect 19660 40772 19716 40828
rect 19716 40772 19720 40828
rect 19656 40768 19720 40772
rect 19736 40828 19800 40832
rect 19736 40772 19740 40828
rect 19740 40772 19796 40828
rect 19796 40772 19800 40828
rect 19736 40768 19800 40772
rect 19816 40828 19880 40832
rect 19816 40772 19820 40828
rect 19820 40772 19876 40828
rect 19876 40772 19880 40828
rect 19816 40768 19880 40772
rect 50296 40828 50360 40832
rect 50296 40772 50300 40828
rect 50300 40772 50356 40828
rect 50356 40772 50360 40828
rect 50296 40768 50360 40772
rect 50376 40828 50440 40832
rect 50376 40772 50380 40828
rect 50380 40772 50436 40828
rect 50436 40772 50440 40828
rect 50376 40768 50440 40772
rect 50456 40828 50520 40832
rect 50456 40772 50460 40828
rect 50460 40772 50516 40828
rect 50516 40772 50520 40828
rect 50456 40768 50520 40772
rect 50536 40828 50600 40832
rect 50536 40772 50540 40828
rect 50540 40772 50596 40828
rect 50596 40772 50600 40828
rect 50536 40768 50600 40772
rect 81016 40828 81080 40832
rect 81016 40772 81020 40828
rect 81020 40772 81076 40828
rect 81076 40772 81080 40828
rect 81016 40768 81080 40772
rect 81096 40828 81160 40832
rect 81096 40772 81100 40828
rect 81100 40772 81156 40828
rect 81156 40772 81160 40828
rect 81096 40768 81160 40772
rect 81176 40828 81240 40832
rect 81176 40772 81180 40828
rect 81180 40772 81236 40828
rect 81236 40772 81240 40828
rect 81176 40768 81240 40772
rect 81256 40828 81320 40832
rect 81256 40772 81260 40828
rect 81260 40772 81316 40828
rect 81316 40772 81320 40828
rect 81256 40768 81320 40772
rect 111736 40828 111800 40832
rect 111736 40772 111740 40828
rect 111740 40772 111796 40828
rect 111796 40772 111800 40828
rect 111736 40768 111800 40772
rect 111816 40828 111880 40832
rect 111816 40772 111820 40828
rect 111820 40772 111876 40828
rect 111876 40772 111880 40828
rect 111816 40768 111880 40772
rect 111896 40828 111960 40832
rect 111896 40772 111900 40828
rect 111900 40772 111956 40828
rect 111956 40772 111960 40828
rect 111896 40768 111960 40772
rect 111976 40828 112040 40832
rect 111976 40772 111980 40828
rect 111980 40772 112036 40828
rect 112036 40772 112040 40828
rect 111976 40768 112040 40772
rect 142456 40828 142520 40832
rect 142456 40772 142460 40828
rect 142460 40772 142516 40828
rect 142516 40772 142520 40828
rect 142456 40768 142520 40772
rect 142536 40828 142600 40832
rect 142536 40772 142540 40828
rect 142540 40772 142596 40828
rect 142596 40772 142600 40828
rect 142536 40768 142600 40772
rect 142616 40828 142680 40832
rect 142616 40772 142620 40828
rect 142620 40772 142676 40828
rect 142676 40772 142680 40828
rect 142616 40768 142680 40772
rect 142696 40828 142760 40832
rect 142696 40772 142700 40828
rect 142700 40772 142756 40828
rect 142756 40772 142760 40828
rect 142696 40768 142760 40772
rect 173176 40828 173240 40832
rect 173176 40772 173180 40828
rect 173180 40772 173236 40828
rect 173236 40772 173240 40828
rect 173176 40768 173240 40772
rect 173256 40828 173320 40832
rect 173256 40772 173260 40828
rect 173260 40772 173316 40828
rect 173316 40772 173320 40828
rect 173256 40768 173320 40772
rect 173336 40828 173400 40832
rect 173336 40772 173340 40828
rect 173340 40772 173396 40828
rect 173396 40772 173400 40828
rect 173336 40768 173400 40772
rect 173416 40828 173480 40832
rect 173416 40772 173420 40828
rect 173420 40772 173476 40828
rect 173476 40772 173480 40828
rect 173416 40768 173480 40772
rect 4216 40284 4280 40288
rect 4216 40228 4220 40284
rect 4220 40228 4276 40284
rect 4276 40228 4280 40284
rect 4216 40224 4280 40228
rect 4296 40284 4360 40288
rect 4296 40228 4300 40284
rect 4300 40228 4356 40284
rect 4356 40228 4360 40284
rect 4296 40224 4360 40228
rect 4376 40284 4440 40288
rect 4376 40228 4380 40284
rect 4380 40228 4436 40284
rect 4436 40228 4440 40284
rect 4376 40224 4440 40228
rect 4456 40284 4520 40288
rect 4456 40228 4460 40284
rect 4460 40228 4516 40284
rect 4516 40228 4520 40284
rect 4456 40224 4520 40228
rect 34936 40284 35000 40288
rect 34936 40228 34940 40284
rect 34940 40228 34996 40284
rect 34996 40228 35000 40284
rect 34936 40224 35000 40228
rect 35016 40284 35080 40288
rect 35016 40228 35020 40284
rect 35020 40228 35076 40284
rect 35076 40228 35080 40284
rect 35016 40224 35080 40228
rect 35096 40284 35160 40288
rect 35096 40228 35100 40284
rect 35100 40228 35156 40284
rect 35156 40228 35160 40284
rect 35096 40224 35160 40228
rect 35176 40284 35240 40288
rect 35176 40228 35180 40284
rect 35180 40228 35236 40284
rect 35236 40228 35240 40284
rect 35176 40224 35240 40228
rect 65656 40284 65720 40288
rect 65656 40228 65660 40284
rect 65660 40228 65716 40284
rect 65716 40228 65720 40284
rect 65656 40224 65720 40228
rect 65736 40284 65800 40288
rect 65736 40228 65740 40284
rect 65740 40228 65796 40284
rect 65796 40228 65800 40284
rect 65736 40224 65800 40228
rect 65816 40284 65880 40288
rect 65816 40228 65820 40284
rect 65820 40228 65876 40284
rect 65876 40228 65880 40284
rect 65816 40224 65880 40228
rect 65896 40284 65960 40288
rect 65896 40228 65900 40284
rect 65900 40228 65956 40284
rect 65956 40228 65960 40284
rect 65896 40224 65960 40228
rect 96376 40284 96440 40288
rect 96376 40228 96380 40284
rect 96380 40228 96436 40284
rect 96436 40228 96440 40284
rect 96376 40224 96440 40228
rect 96456 40284 96520 40288
rect 96456 40228 96460 40284
rect 96460 40228 96516 40284
rect 96516 40228 96520 40284
rect 96456 40224 96520 40228
rect 96536 40284 96600 40288
rect 96536 40228 96540 40284
rect 96540 40228 96596 40284
rect 96596 40228 96600 40284
rect 96536 40224 96600 40228
rect 96616 40284 96680 40288
rect 96616 40228 96620 40284
rect 96620 40228 96676 40284
rect 96676 40228 96680 40284
rect 96616 40224 96680 40228
rect 127096 40284 127160 40288
rect 127096 40228 127100 40284
rect 127100 40228 127156 40284
rect 127156 40228 127160 40284
rect 127096 40224 127160 40228
rect 127176 40284 127240 40288
rect 127176 40228 127180 40284
rect 127180 40228 127236 40284
rect 127236 40228 127240 40284
rect 127176 40224 127240 40228
rect 127256 40284 127320 40288
rect 127256 40228 127260 40284
rect 127260 40228 127316 40284
rect 127316 40228 127320 40284
rect 127256 40224 127320 40228
rect 127336 40284 127400 40288
rect 127336 40228 127340 40284
rect 127340 40228 127396 40284
rect 127396 40228 127400 40284
rect 127336 40224 127400 40228
rect 157816 40284 157880 40288
rect 157816 40228 157820 40284
rect 157820 40228 157876 40284
rect 157876 40228 157880 40284
rect 157816 40224 157880 40228
rect 157896 40284 157960 40288
rect 157896 40228 157900 40284
rect 157900 40228 157956 40284
rect 157956 40228 157960 40284
rect 157896 40224 157960 40228
rect 157976 40284 158040 40288
rect 157976 40228 157980 40284
rect 157980 40228 158036 40284
rect 158036 40228 158040 40284
rect 157976 40224 158040 40228
rect 158056 40284 158120 40288
rect 158056 40228 158060 40284
rect 158060 40228 158116 40284
rect 158116 40228 158120 40284
rect 158056 40224 158120 40228
rect 19576 39740 19640 39744
rect 19576 39684 19580 39740
rect 19580 39684 19636 39740
rect 19636 39684 19640 39740
rect 19576 39680 19640 39684
rect 19656 39740 19720 39744
rect 19656 39684 19660 39740
rect 19660 39684 19716 39740
rect 19716 39684 19720 39740
rect 19656 39680 19720 39684
rect 19736 39740 19800 39744
rect 19736 39684 19740 39740
rect 19740 39684 19796 39740
rect 19796 39684 19800 39740
rect 19736 39680 19800 39684
rect 19816 39740 19880 39744
rect 19816 39684 19820 39740
rect 19820 39684 19876 39740
rect 19876 39684 19880 39740
rect 19816 39680 19880 39684
rect 50296 39740 50360 39744
rect 50296 39684 50300 39740
rect 50300 39684 50356 39740
rect 50356 39684 50360 39740
rect 50296 39680 50360 39684
rect 50376 39740 50440 39744
rect 50376 39684 50380 39740
rect 50380 39684 50436 39740
rect 50436 39684 50440 39740
rect 50376 39680 50440 39684
rect 50456 39740 50520 39744
rect 50456 39684 50460 39740
rect 50460 39684 50516 39740
rect 50516 39684 50520 39740
rect 50456 39680 50520 39684
rect 50536 39740 50600 39744
rect 50536 39684 50540 39740
rect 50540 39684 50596 39740
rect 50596 39684 50600 39740
rect 50536 39680 50600 39684
rect 81016 39740 81080 39744
rect 81016 39684 81020 39740
rect 81020 39684 81076 39740
rect 81076 39684 81080 39740
rect 81016 39680 81080 39684
rect 81096 39740 81160 39744
rect 81096 39684 81100 39740
rect 81100 39684 81156 39740
rect 81156 39684 81160 39740
rect 81096 39680 81160 39684
rect 81176 39740 81240 39744
rect 81176 39684 81180 39740
rect 81180 39684 81236 39740
rect 81236 39684 81240 39740
rect 81176 39680 81240 39684
rect 81256 39740 81320 39744
rect 81256 39684 81260 39740
rect 81260 39684 81316 39740
rect 81316 39684 81320 39740
rect 81256 39680 81320 39684
rect 111736 39740 111800 39744
rect 111736 39684 111740 39740
rect 111740 39684 111796 39740
rect 111796 39684 111800 39740
rect 111736 39680 111800 39684
rect 111816 39740 111880 39744
rect 111816 39684 111820 39740
rect 111820 39684 111876 39740
rect 111876 39684 111880 39740
rect 111816 39680 111880 39684
rect 111896 39740 111960 39744
rect 111896 39684 111900 39740
rect 111900 39684 111956 39740
rect 111956 39684 111960 39740
rect 111896 39680 111960 39684
rect 111976 39740 112040 39744
rect 111976 39684 111980 39740
rect 111980 39684 112036 39740
rect 112036 39684 112040 39740
rect 111976 39680 112040 39684
rect 142456 39740 142520 39744
rect 142456 39684 142460 39740
rect 142460 39684 142516 39740
rect 142516 39684 142520 39740
rect 142456 39680 142520 39684
rect 142536 39740 142600 39744
rect 142536 39684 142540 39740
rect 142540 39684 142596 39740
rect 142596 39684 142600 39740
rect 142536 39680 142600 39684
rect 142616 39740 142680 39744
rect 142616 39684 142620 39740
rect 142620 39684 142676 39740
rect 142676 39684 142680 39740
rect 142616 39680 142680 39684
rect 142696 39740 142760 39744
rect 142696 39684 142700 39740
rect 142700 39684 142756 39740
rect 142756 39684 142760 39740
rect 142696 39680 142760 39684
rect 173176 39740 173240 39744
rect 173176 39684 173180 39740
rect 173180 39684 173236 39740
rect 173236 39684 173240 39740
rect 173176 39680 173240 39684
rect 173256 39740 173320 39744
rect 173256 39684 173260 39740
rect 173260 39684 173316 39740
rect 173316 39684 173320 39740
rect 173256 39680 173320 39684
rect 173336 39740 173400 39744
rect 173336 39684 173340 39740
rect 173340 39684 173396 39740
rect 173396 39684 173400 39740
rect 173336 39680 173400 39684
rect 173416 39740 173480 39744
rect 173416 39684 173420 39740
rect 173420 39684 173476 39740
rect 173476 39684 173480 39740
rect 173416 39680 173480 39684
rect 4216 39196 4280 39200
rect 4216 39140 4220 39196
rect 4220 39140 4276 39196
rect 4276 39140 4280 39196
rect 4216 39136 4280 39140
rect 4296 39196 4360 39200
rect 4296 39140 4300 39196
rect 4300 39140 4356 39196
rect 4356 39140 4360 39196
rect 4296 39136 4360 39140
rect 4376 39196 4440 39200
rect 4376 39140 4380 39196
rect 4380 39140 4436 39196
rect 4436 39140 4440 39196
rect 4376 39136 4440 39140
rect 4456 39196 4520 39200
rect 4456 39140 4460 39196
rect 4460 39140 4516 39196
rect 4516 39140 4520 39196
rect 4456 39136 4520 39140
rect 34936 39196 35000 39200
rect 34936 39140 34940 39196
rect 34940 39140 34996 39196
rect 34996 39140 35000 39196
rect 34936 39136 35000 39140
rect 35016 39196 35080 39200
rect 35016 39140 35020 39196
rect 35020 39140 35076 39196
rect 35076 39140 35080 39196
rect 35016 39136 35080 39140
rect 35096 39196 35160 39200
rect 35096 39140 35100 39196
rect 35100 39140 35156 39196
rect 35156 39140 35160 39196
rect 35096 39136 35160 39140
rect 35176 39196 35240 39200
rect 35176 39140 35180 39196
rect 35180 39140 35236 39196
rect 35236 39140 35240 39196
rect 35176 39136 35240 39140
rect 65656 39196 65720 39200
rect 65656 39140 65660 39196
rect 65660 39140 65716 39196
rect 65716 39140 65720 39196
rect 65656 39136 65720 39140
rect 65736 39196 65800 39200
rect 65736 39140 65740 39196
rect 65740 39140 65796 39196
rect 65796 39140 65800 39196
rect 65736 39136 65800 39140
rect 65816 39196 65880 39200
rect 65816 39140 65820 39196
rect 65820 39140 65876 39196
rect 65876 39140 65880 39196
rect 65816 39136 65880 39140
rect 65896 39196 65960 39200
rect 65896 39140 65900 39196
rect 65900 39140 65956 39196
rect 65956 39140 65960 39196
rect 65896 39136 65960 39140
rect 96376 39196 96440 39200
rect 96376 39140 96380 39196
rect 96380 39140 96436 39196
rect 96436 39140 96440 39196
rect 96376 39136 96440 39140
rect 96456 39196 96520 39200
rect 96456 39140 96460 39196
rect 96460 39140 96516 39196
rect 96516 39140 96520 39196
rect 96456 39136 96520 39140
rect 96536 39196 96600 39200
rect 96536 39140 96540 39196
rect 96540 39140 96596 39196
rect 96596 39140 96600 39196
rect 96536 39136 96600 39140
rect 96616 39196 96680 39200
rect 96616 39140 96620 39196
rect 96620 39140 96676 39196
rect 96676 39140 96680 39196
rect 96616 39136 96680 39140
rect 127096 39196 127160 39200
rect 127096 39140 127100 39196
rect 127100 39140 127156 39196
rect 127156 39140 127160 39196
rect 127096 39136 127160 39140
rect 127176 39196 127240 39200
rect 127176 39140 127180 39196
rect 127180 39140 127236 39196
rect 127236 39140 127240 39196
rect 127176 39136 127240 39140
rect 127256 39196 127320 39200
rect 127256 39140 127260 39196
rect 127260 39140 127316 39196
rect 127316 39140 127320 39196
rect 127256 39136 127320 39140
rect 127336 39196 127400 39200
rect 127336 39140 127340 39196
rect 127340 39140 127396 39196
rect 127396 39140 127400 39196
rect 127336 39136 127400 39140
rect 157816 39196 157880 39200
rect 157816 39140 157820 39196
rect 157820 39140 157876 39196
rect 157876 39140 157880 39196
rect 157816 39136 157880 39140
rect 157896 39196 157960 39200
rect 157896 39140 157900 39196
rect 157900 39140 157956 39196
rect 157956 39140 157960 39196
rect 157896 39136 157960 39140
rect 157976 39196 158040 39200
rect 157976 39140 157980 39196
rect 157980 39140 158036 39196
rect 158036 39140 158040 39196
rect 157976 39136 158040 39140
rect 158056 39196 158120 39200
rect 158056 39140 158060 39196
rect 158060 39140 158116 39196
rect 158116 39140 158120 39196
rect 158056 39136 158120 39140
rect 19576 38652 19640 38656
rect 19576 38596 19580 38652
rect 19580 38596 19636 38652
rect 19636 38596 19640 38652
rect 19576 38592 19640 38596
rect 19656 38652 19720 38656
rect 19656 38596 19660 38652
rect 19660 38596 19716 38652
rect 19716 38596 19720 38652
rect 19656 38592 19720 38596
rect 19736 38652 19800 38656
rect 19736 38596 19740 38652
rect 19740 38596 19796 38652
rect 19796 38596 19800 38652
rect 19736 38592 19800 38596
rect 19816 38652 19880 38656
rect 19816 38596 19820 38652
rect 19820 38596 19876 38652
rect 19876 38596 19880 38652
rect 19816 38592 19880 38596
rect 50296 38652 50360 38656
rect 50296 38596 50300 38652
rect 50300 38596 50356 38652
rect 50356 38596 50360 38652
rect 50296 38592 50360 38596
rect 50376 38652 50440 38656
rect 50376 38596 50380 38652
rect 50380 38596 50436 38652
rect 50436 38596 50440 38652
rect 50376 38592 50440 38596
rect 50456 38652 50520 38656
rect 50456 38596 50460 38652
rect 50460 38596 50516 38652
rect 50516 38596 50520 38652
rect 50456 38592 50520 38596
rect 50536 38652 50600 38656
rect 50536 38596 50540 38652
rect 50540 38596 50596 38652
rect 50596 38596 50600 38652
rect 50536 38592 50600 38596
rect 81016 38652 81080 38656
rect 81016 38596 81020 38652
rect 81020 38596 81076 38652
rect 81076 38596 81080 38652
rect 81016 38592 81080 38596
rect 81096 38652 81160 38656
rect 81096 38596 81100 38652
rect 81100 38596 81156 38652
rect 81156 38596 81160 38652
rect 81096 38592 81160 38596
rect 81176 38652 81240 38656
rect 81176 38596 81180 38652
rect 81180 38596 81236 38652
rect 81236 38596 81240 38652
rect 81176 38592 81240 38596
rect 81256 38652 81320 38656
rect 81256 38596 81260 38652
rect 81260 38596 81316 38652
rect 81316 38596 81320 38652
rect 81256 38592 81320 38596
rect 111736 38652 111800 38656
rect 111736 38596 111740 38652
rect 111740 38596 111796 38652
rect 111796 38596 111800 38652
rect 111736 38592 111800 38596
rect 111816 38652 111880 38656
rect 111816 38596 111820 38652
rect 111820 38596 111876 38652
rect 111876 38596 111880 38652
rect 111816 38592 111880 38596
rect 111896 38652 111960 38656
rect 111896 38596 111900 38652
rect 111900 38596 111956 38652
rect 111956 38596 111960 38652
rect 111896 38592 111960 38596
rect 111976 38652 112040 38656
rect 111976 38596 111980 38652
rect 111980 38596 112036 38652
rect 112036 38596 112040 38652
rect 111976 38592 112040 38596
rect 142456 38652 142520 38656
rect 142456 38596 142460 38652
rect 142460 38596 142516 38652
rect 142516 38596 142520 38652
rect 142456 38592 142520 38596
rect 142536 38652 142600 38656
rect 142536 38596 142540 38652
rect 142540 38596 142596 38652
rect 142596 38596 142600 38652
rect 142536 38592 142600 38596
rect 142616 38652 142680 38656
rect 142616 38596 142620 38652
rect 142620 38596 142676 38652
rect 142676 38596 142680 38652
rect 142616 38592 142680 38596
rect 142696 38652 142760 38656
rect 142696 38596 142700 38652
rect 142700 38596 142756 38652
rect 142756 38596 142760 38652
rect 142696 38592 142760 38596
rect 173176 38652 173240 38656
rect 173176 38596 173180 38652
rect 173180 38596 173236 38652
rect 173236 38596 173240 38652
rect 173176 38592 173240 38596
rect 173256 38652 173320 38656
rect 173256 38596 173260 38652
rect 173260 38596 173316 38652
rect 173316 38596 173320 38652
rect 173256 38592 173320 38596
rect 173336 38652 173400 38656
rect 173336 38596 173340 38652
rect 173340 38596 173396 38652
rect 173396 38596 173400 38652
rect 173336 38592 173400 38596
rect 173416 38652 173480 38656
rect 173416 38596 173420 38652
rect 173420 38596 173476 38652
rect 173476 38596 173480 38652
rect 173416 38592 173480 38596
rect 4216 38108 4280 38112
rect 4216 38052 4220 38108
rect 4220 38052 4276 38108
rect 4276 38052 4280 38108
rect 4216 38048 4280 38052
rect 4296 38108 4360 38112
rect 4296 38052 4300 38108
rect 4300 38052 4356 38108
rect 4356 38052 4360 38108
rect 4296 38048 4360 38052
rect 4376 38108 4440 38112
rect 4376 38052 4380 38108
rect 4380 38052 4436 38108
rect 4436 38052 4440 38108
rect 4376 38048 4440 38052
rect 4456 38108 4520 38112
rect 4456 38052 4460 38108
rect 4460 38052 4516 38108
rect 4516 38052 4520 38108
rect 4456 38048 4520 38052
rect 34936 38108 35000 38112
rect 34936 38052 34940 38108
rect 34940 38052 34996 38108
rect 34996 38052 35000 38108
rect 34936 38048 35000 38052
rect 35016 38108 35080 38112
rect 35016 38052 35020 38108
rect 35020 38052 35076 38108
rect 35076 38052 35080 38108
rect 35016 38048 35080 38052
rect 35096 38108 35160 38112
rect 35096 38052 35100 38108
rect 35100 38052 35156 38108
rect 35156 38052 35160 38108
rect 35096 38048 35160 38052
rect 35176 38108 35240 38112
rect 35176 38052 35180 38108
rect 35180 38052 35236 38108
rect 35236 38052 35240 38108
rect 35176 38048 35240 38052
rect 65656 38108 65720 38112
rect 65656 38052 65660 38108
rect 65660 38052 65716 38108
rect 65716 38052 65720 38108
rect 65656 38048 65720 38052
rect 65736 38108 65800 38112
rect 65736 38052 65740 38108
rect 65740 38052 65796 38108
rect 65796 38052 65800 38108
rect 65736 38048 65800 38052
rect 65816 38108 65880 38112
rect 65816 38052 65820 38108
rect 65820 38052 65876 38108
rect 65876 38052 65880 38108
rect 65816 38048 65880 38052
rect 65896 38108 65960 38112
rect 65896 38052 65900 38108
rect 65900 38052 65956 38108
rect 65956 38052 65960 38108
rect 65896 38048 65960 38052
rect 96376 38108 96440 38112
rect 96376 38052 96380 38108
rect 96380 38052 96436 38108
rect 96436 38052 96440 38108
rect 96376 38048 96440 38052
rect 96456 38108 96520 38112
rect 96456 38052 96460 38108
rect 96460 38052 96516 38108
rect 96516 38052 96520 38108
rect 96456 38048 96520 38052
rect 96536 38108 96600 38112
rect 96536 38052 96540 38108
rect 96540 38052 96596 38108
rect 96596 38052 96600 38108
rect 96536 38048 96600 38052
rect 96616 38108 96680 38112
rect 96616 38052 96620 38108
rect 96620 38052 96676 38108
rect 96676 38052 96680 38108
rect 96616 38048 96680 38052
rect 127096 38108 127160 38112
rect 127096 38052 127100 38108
rect 127100 38052 127156 38108
rect 127156 38052 127160 38108
rect 127096 38048 127160 38052
rect 127176 38108 127240 38112
rect 127176 38052 127180 38108
rect 127180 38052 127236 38108
rect 127236 38052 127240 38108
rect 127176 38048 127240 38052
rect 127256 38108 127320 38112
rect 127256 38052 127260 38108
rect 127260 38052 127316 38108
rect 127316 38052 127320 38108
rect 127256 38048 127320 38052
rect 127336 38108 127400 38112
rect 127336 38052 127340 38108
rect 127340 38052 127396 38108
rect 127396 38052 127400 38108
rect 127336 38048 127400 38052
rect 157816 38108 157880 38112
rect 157816 38052 157820 38108
rect 157820 38052 157876 38108
rect 157876 38052 157880 38108
rect 157816 38048 157880 38052
rect 157896 38108 157960 38112
rect 157896 38052 157900 38108
rect 157900 38052 157956 38108
rect 157956 38052 157960 38108
rect 157896 38048 157960 38052
rect 157976 38108 158040 38112
rect 157976 38052 157980 38108
rect 157980 38052 158036 38108
rect 158036 38052 158040 38108
rect 157976 38048 158040 38052
rect 158056 38108 158120 38112
rect 158056 38052 158060 38108
rect 158060 38052 158116 38108
rect 158116 38052 158120 38108
rect 158056 38048 158120 38052
rect 19576 37564 19640 37568
rect 19576 37508 19580 37564
rect 19580 37508 19636 37564
rect 19636 37508 19640 37564
rect 19576 37504 19640 37508
rect 19656 37564 19720 37568
rect 19656 37508 19660 37564
rect 19660 37508 19716 37564
rect 19716 37508 19720 37564
rect 19656 37504 19720 37508
rect 19736 37564 19800 37568
rect 19736 37508 19740 37564
rect 19740 37508 19796 37564
rect 19796 37508 19800 37564
rect 19736 37504 19800 37508
rect 19816 37564 19880 37568
rect 19816 37508 19820 37564
rect 19820 37508 19876 37564
rect 19876 37508 19880 37564
rect 19816 37504 19880 37508
rect 50296 37564 50360 37568
rect 50296 37508 50300 37564
rect 50300 37508 50356 37564
rect 50356 37508 50360 37564
rect 50296 37504 50360 37508
rect 50376 37564 50440 37568
rect 50376 37508 50380 37564
rect 50380 37508 50436 37564
rect 50436 37508 50440 37564
rect 50376 37504 50440 37508
rect 50456 37564 50520 37568
rect 50456 37508 50460 37564
rect 50460 37508 50516 37564
rect 50516 37508 50520 37564
rect 50456 37504 50520 37508
rect 50536 37564 50600 37568
rect 50536 37508 50540 37564
rect 50540 37508 50596 37564
rect 50596 37508 50600 37564
rect 50536 37504 50600 37508
rect 81016 37564 81080 37568
rect 81016 37508 81020 37564
rect 81020 37508 81076 37564
rect 81076 37508 81080 37564
rect 81016 37504 81080 37508
rect 81096 37564 81160 37568
rect 81096 37508 81100 37564
rect 81100 37508 81156 37564
rect 81156 37508 81160 37564
rect 81096 37504 81160 37508
rect 81176 37564 81240 37568
rect 81176 37508 81180 37564
rect 81180 37508 81236 37564
rect 81236 37508 81240 37564
rect 81176 37504 81240 37508
rect 81256 37564 81320 37568
rect 81256 37508 81260 37564
rect 81260 37508 81316 37564
rect 81316 37508 81320 37564
rect 81256 37504 81320 37508
rect 111736 37564 111800 37568
rect 111736 37508 111740 37564
rect 111740 37508 111796 37564
rect 111796 37508 111800 37564
rect 111736 37504 111800 37508
rect 111816 37564 111880 37568
rect 111816 37508 111820 37564
rect 111820 37508 111876 37564
rect 111876 37508 111880 37564
rect 111816 37504 111880 37508
rect 111896 37564 111960 37568
rect 111896 37508 111900 37564
rect 111900 37508 111956 37564
rect 111956 37508 111960 37564
rect 111896 37504 111960 37508
rect 111976 37564 112040 37568
rect 111976 37508 111980 37564
rect 111980 37508 112036 37564
rect 112036 37508 112040 37564
rect 111976 37504 112040 37508
rect 142456 37564 142520 37568
rect 142456 37508 142460 37564
rect 142460 37508 142516 37564
rect 142516 37508 142520 37564
rect 142456 37504 142520 37508
rect 142536 37564 142600 37568
rect 142536 37508 142540 37564
rect 142540 37508 142596 37564
rect 142596 37508 142600 37564
rect 142536 37504 142600 37508
rect 142616 37564 142680 37568
rect 142616 37508 142620 37564
rect 142620 37508 142676 37564
rect 142676 37508 142680 37564
rect 142616 37504 142680 37508
rect 142696 37564 142760 37568
rect 142696 37508 142700 37564
rect 142700 37508 142756 37564
rect 142756 37508 142760 37564
rect 142696 37504 142760 37508
rect 173176 37564 173240 37568
rect 173176 37508 173180 37564
rect 173180 37508 173236 37564
rect 173236 37508 173240 37564
rect 173176 37504 173240 37508
rect 173256 37564 173320 37568
rect 173256 37508 173260 37564
rect 173260 37508 173316 37564
rect 173316 37508 173320 37564
rect 173256 37504 173320 37508
rect 173336 37564 173400 37568
rect 173336 37508 173340 37564
rect 173340 37508 173396 37564
rect 173396 37508 173400 37564
rect 173336 37504 173400 37508
rect 173416 37564 173480 37568
rect 173416 37508 173420 37564
rect 173420 37508 173476 37564
rect 173476 37508 173480 37564
rect 173416 37504 173480 37508
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 34936 37020 35000 37024
rect 34936 36964 34940 37020
rect 34940 36964 34996 37020
rect 34996 36964 35000 37020
rect 34936 36960 35000 36964
rect 35016 37020 35080 37024
rect 35016 36964 35020 37020
rect 35020 36964 35076 37020
rect 35076 36964 35080 37020
rect 35016 36960 35080 36964
rect 35096 37020 35160 37024
rect 35096 36964 35100 37020
rect 35100 36964 35156 37020
rect 35156 36964 35160 37020
rect 35096 36960 35160 36964
rect 35176 37020 35240 37024
rect 35176 36964 35180 37020
rect 35180 36964 35236 37020
rect 35236 36964 35240 37020
rect 35176 36960 35240 36964
rect 65656 37020 65720 37024
rect 65656 36964 65660 37020
rect 65660 36964 65716 37020
rect 65716 36964 65720 37020
rect 65656 36960 65720 36964
rect 65736 37020 65800 37024
rect 65736 36964 65740 37020
rect 65740 36964 65796 37020
rect 65796 36964 65800 37020
rect 65736 36960 65800 36964
rect 65816 37020 65880 37024
rect 65816 36964 65820 37020
rect 65820 36964 65876 37020
rect 65876 36964 65880 37020
rect 65816 36960 65880 36964
rect 65896 37020 65960 37024
rect 65896 36964 65900 37020
rect 65900 36964 65956 37020
rect 65956 36964 65960 37020
rect 65896 36960 65960 36964
rect 96376 37020 96440 37024
rect 96376 36964 96380 37020
rect 96380 36964 96436 37020
rect 96436 36964 96440 37020
rect 96376 36960 96440 36964
rect 96456 37020 96520 37024
rect 96456 36964 96460 37020
rect 96460 36964 96516 37020
rect 96516 36964 96520 37020
rect 96456 36960 96520 36964
rect 96536 37020 96600 37024
rect 96536 36964 96540 37020
rect 96540 36964 96596 37020
rect 96596 36964 96600 37020
rect 96536 36960 96600 36964
rect 96616 37020 96680 37024
rect 96616 36964 96620 37020
rect 96620 36964 96676 37020
rect 96676 36964 96680 37020
rect 96616 36960 96680 36964
rect 127096 37020 127160 37024
rect 127096 36964 127100 37020
rect 127100 36964 127156 37020
rect 127156 36964 127160 37020
rect 127096 36960 127160 36964
rect 127176 37020 127240 37024
rect 127176 36964 127180 37020
rect 127180 36964 127236 37020
rect 127236 36964 127240 37020
rect 127176 36960 127240 36964
rect 127256 37020 127320 37024
rect 127256 36964 127260 37020
rect 127260 36964 127316 37020
rect 127316 36964 127320 37020
rect 127256 36960 127320 36964
rect 127336 37020 127400 37024
rect 127336 36964 127340 37020
rect 127340 36964 127396 37020
rect 127396 36964 127400 37020
rect 127336 36960 127400 36964
rect 157816 37020 157880 37024
rect 157816 36964 157820 37020
rect 157820 36964 157876 37020
rect 157876 36964 157880 37020
rect 157816 36960 157880 36964
rect 157896 37020 157960 37024
rect 157896 36964 157900 37020
rect 157900 36964 157956 37020
rect 157956 36964 157960 37020
rect 157896 36960 157960 36964
rect 157976 37020 158040 37024
rect 157976 36964 157980 37020
rect 157980 36964 158036 37020
rect 158036 36964 158040 37020
rect 157976 36960 158040 36964
rect 158056 37020 158120 37024
rect 158056 36964 158060 37020
rect 158060 36964 158116 37020
rect 158116 36964 158120 37020
rect 158056 36960 158120 36964
rect 19576 36476 19640 36480
rect 19576 36420 19580 36476
rect 19580 36420 19636 36476
rect 19636 36420 19640 36476
rect 19576 36416 19640 36420
rect 19656 36476 19720 36480
rect 19656 36420 19660 36476
rect 19660 36420 19716 36476
rect 19716 36420 19720 36476
rect 19656 36416 19720 36420
rect 19736 36476 19800 36480
rect 19736 36420 19740 36476
rect 19740 36420 19796 36476
rect 19796 36420 19800 36476
rect 19736 36416 19800 36420
rect 19816 36476 19880 36480
rect 19816 36420 19820 36476
rect 19820 36420 19876 36476
rect 19876 36420 19880 36476
rect 19816 36416 19880 36420
rect 50296 36476 50360 36480
rect 50296 36420 50300 36476
rect 50300 36420 50356 36476
rect 50356 36420 50360 36476
rect 50296 36416 50360 36420
rect 50376 36476 50440 36480
rect 50376 36420 50380 36476
rect 50380 36420 50436 36476
rect 50436 36420 50440 36476
rect 50376 36416 50440 36420
rect 50456 36476 50520 36480
rect 50456 36420 50460 36476
rect 50460 36420 50516 36476
rect 50516 36420 50520 36476
rect 50456 36416 50520 36420
rect 50536 36476 50600 36480
rect 50536 36420 50540 36476
rect 50540 36420 50596 36476
rect 50596 36420 50600 36476
rect 50536 36416 50600 36420
rect 81016 36476 81080 36480
rect 81016 36420 81020 36476
rect 81020 36420 81076 36476
rect 81076 36420 81080 36476
rect 81016 36416 81080 36420
rect 81096 36476 81160 36480
rect 81096 36420 81100 36476
rect 81100 36420 81156 36476
rect 81156 36420 81160 36476
rect 81096 36416 81160 36420
rect 81176 36476 81240 36480
rect 81176 36420 81180 36476
rect 81180 36420 81236 36476
rect 81236 36420 81240 36476
rect 81176 36416 81240 36420
rect 81256 36476 81320 36480
rect 81256 36420 81260 36476
rect 81260 36420 81316 36476
rect 81316 36420 81320 36476
rect 81256 36416 81320 36420
rect 111736 36476 111800 36480
rect 111736 36420 111740 36476
rect 111740 36420 111796 36476
rect 111796 36420 111800 36476
rect 111736 36416 111800 36420
rect 111816 36476 111880 36480
rect 111816 36420 111820 36476
rect 111820 36420 111876 36476
rect 111876 36420 111880 36476
rect 111816 36416 111880 36420
rect 111896 36476 111960 36480
rect 111896 36420 111900 36476
rect 111900 36420 111956 36476
rect 111956 36420 111960 36476
rect 111896 36416 111960 36420
rect 111976 36476 112040 36480
rect 111976 36420 111980 36476
rect 111980 36420 112036 36476
rect 112036 36420 112040 36476
rect 111976 36416 112040 36420
rect 142456 36476 142520 36480
rect 142456 36420 142460 36476
rect 142460 36420 142516 36476
rect 142516 36420 142520 36476
rect 142456 36416 142520 36420
rect 142536 36476 142600 36480
rect 142536 36420 142540 36476
rect 142540 36420 142596 36476
rect 142596 36420 142600 36476
rect 142536 36416 142600 36420
rect 142616 36476 142680 36480
rect 142616 36420 142620 36476
rect 142620 36420 142676 36476
rect 142676 36420 142680 36476
rect 142616 36416 142680 36420
rect 142696 36476 142760 36480
rect 142696 36420 142700 36476
rect 142700 36420 142756 36476
rect 142756 36420 142760 36476
rect 142696 36416 142760 36420
rect 173176 36476 173240 36480
rect 173176 36420 173180 36476
rect 173180 36420 173236 36476
rect 173236 36420 173240 36476
rect 173176 36416 173240 36420
rect 173256 36476 173320 36480
rect 173256 36420 173260 36476
rect 173260 36420 173316 36476
rect 173316 36420 173320 36476
rect 173256 36416 173320 36420
rect 173336 36476 173400 36480
rect 173336 36420 173340 36476
rect 173340 36420 173396 36476
rect 173396 36420 173400 36476
rect 173336 36416 173400 36420
rect 173416 36476 173480 36480
rect 173416 36420 173420 36476
rect 173420 36420 173476 36476
rect 173476 36420 173480 36476
rect 173416 36416 173480 36420
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 34936 35932 35000 35936
rect 34936 35876 34940 35932
rect 34940 35876 34996 35932
rect 34996 35876 35000 35932
rect 34936 35872 35000 35876
rect 35016 35932 35080 35936
rect 35016 35876 35020 35932
rect 35020 35876 35076 35932
rect 35076 35876 35080 35932
rect 35016 35872 35080 35876
rect 35096 35932 35160 35936
rect 35096 35876 35100 35932
rect 35100 35876 35156 35932
rect 35156 35876 35160 35932
rect 35096 35872 35160 35876
rect 35176 35932 35240 35936
rect 35176 35876 35180 35932
rect 35180 35876 35236 35932
rect 35236 35876 35240 35932
rect 35176 35872 35240 35876
rect 65656 35932 65720 35936
rect 65656 35876 65660 35932
rect 65660 35876 65716 35932
rect 65716 35876 65720 35932
rect 65656 35872 65720 35876
rect 65736 35932 65800 35936
rect 65736 35876 65740 35932
rect 65740 35876 65796 35932
rect 65796 35876 65800 35932
rect 65736 35872 65800 35876
rect 65816 35932 65880 35936
rect 65816 35876 65820 35932
rect 65820 35876 65876 35932
rect 65876 35876 65880 35932
rect 65816 35872 65880 35876
rect 65896 35932 65960 35936
rect 65896 35876 65900 35932
rect 65900 35876 65956 35932
rect 65956 35876 65960 35932
rect 65896 35872 65960 35876
rect 96376 35932 96440 35936
rect 96376 35876 96380 35932
rect 96380 35876 96436 35932
rect 96436 35876 96440 35932
rect 96376 35872 96440 35876
rect 96456 35932 96520 35936
rect 96456 35876 96460 35932
rect 96460 35876 96516 35932
rect 96516 35876 96520 35932
rect 96456 35872 96520 35876
rect 96536 35932 96600 35936
rect 96536 35876 96540 35932
rect 96540 35876 96596 35932
rect 96596 35876 96600 35932
rect 96536 35872 96600 35876
rect 96616 35932 96680 35936
rect 96616 35876 96620 35932
rect 96620 35876 96676 35932
rect 96676 35876 96680 35932
rect 96616 35872 96680 35876
rect 127096 35932 127160 35936
rect 127096 35876 127100 35932
rect 127100 35876 127156 35932
rect 127156 35876 127160 35932
rect 127096 35872 127160 35876
rect 127176 35932 127240 35936
rect 127176 35876 127180 35932
rect 127180 35876 127236 35932
rect 127236 35876 127240 35932
rect 127176 35872 127240 35876
rect 127256 35932 127320 35936
rect 127256 35876 127260 35932
rect 127260 35876 127316 35932
rect 127316 35876 127320 35932
rect 127256 35872 127320 35876
rect 127336 35932 127400 35936
rect 127336 35876 127340 35932
rect 127340 35876 127396 35932
rect 127396 35876 127400 35932
rect 127336 35872 127400 35876
rect 157816 35932 157880 35936
rect 157816 35876 157820 35932
rect 157820 35876 157876 35932
rect 157876 35876 157880 35932
rect 157816 35872 157880 35876
rect 157896 35932 157960 35936
rect 157896 35876 157900 35932
rect 157900 35876 157956 35932
rect 157956 35876 157960 35932
rect 157896 35872 157960 35876
rect 157976 35932 158040 35936
rect 157976 35876 157980 35932
rect 157980 35876 158036 35932
rect 158036 35876 158040 35932
rect 157976 35872 158040 35876
rect 158056 35932 158120 35936
rect 158056 35876 158060 35932
rect 158060 35876 158116 35932
rect 158116 35876 158120 35932
rect 158056 35872 158120 35876
rect 19576 35388 19640 35392
rect 19576 35332 19580 35388
rect 19580 35332 19636 35388
rect 19636 35332 19640 35388
rect 19576 35328 19640 35332
rect 19656 35388 19720 35392
rect 19656 35332 19660 35388
rect 19660 35332 19716 35388
rect 19716 35332 19720 35388
rect 19656 35328 19720 35332
rect 19736 35388 19800 35392
rect 19736 35332 19740 35388
rect 19740 35332 19796 35388
rect 19796 35332 19800 35388
rect 19736 35328 19800 35332
rect 19816 35388 19880 35392
rect 19816 35332 19820 35388
rect 19820 35332 19876 35388
rect 19876 35332 19880 35388
rect 19816 35328 19880 35332
rect 50296 35388 50360 35392
rect 50296 35332 50300 35388
rect 50300 35332 50356 35388
rect 50356 35332 50360 35388
rect 50296 35328 50360 35332
rect 50376 35388 50440 35392
rect 50376 35332 50380 35388
rect 50380 35332 50436 35388
rect 50436 35332 50440 35388
rect 50376 35328 50440 35332
rect 50456 35388 50520 35392
rect 50456 35332 50460 35388
rect 50460 35332 50516 35388
rect 50516 35332 50520 35388
rect 50456 35328 50520 35332
rect 50536 35388 50600 35392
rect 50536 35332 50540 35388
rect 50540 35332 50596 35388
rect 50596 35332 50600 35388
rect 50536 35328 50600 35332
rect 81016 35388 81080 35392
rect 81016 35332 81020 35388
rect 81020 35332 81076 35388
rect 81076 35332 81080 35388
rect 81016 35328 81080 35332
rect 81096 35388 81160 35392
rect 81096 35332 81100 35388
rect 81100 35332 81156 35388
rect 81156 35332 81160 35388
rect 81096 35328 81160 35332
rect 81176 35388 81240 35392
rect 81176 35332 81180 35388
rect 81180 35332 81236 35388
rect 81236 35332 81240 35388
rect 81176 35328 81240 35332
rect 81256 35388 81320 35392
rect 81256 35332 81260 35388
rect 81260 35332 81316 35388
rect 81316 35332 81320 35388
rect 81256 35328 81320 35332
rect 111736 35388 111800 35392
rect 111736 35332 111740 35388
rect 111740 35332 111796 35388
rect 111796 35332 111800 35388
rect 111736 35328 111800 35332
rect 111816 35388 111880 35392
rect 111816 35332 111820 35388
rect 111820 35332 111876 35388
rect 111876 35332 111880 35388
rect 111816 35328 111880 35332
rect 111896 35388 111960 35392
rect 111896 35332 111900 35388
rect 111900 35332 111956 35388
rect 111956 35332 111960 35388
rect 111896 35328 111960 35332
rect 111976 35388 112040 35392
rect 111976 35332 111980 35388
rect 111980 35332 112036 35388
rect 112036 35332 112040 35388
rect 111976 35328 112040 35332
rect 142456 35388 142520 35392
rect 142456 35332 142460 35388
rect 142460 35332 142516 35388
rect 142516 35332 142520 35388
rect 142456 35328 142520 35332
rect 142536 35388 142600 35392
rect 142536 35332 142540 35388
rect 142540 35332 142596 35388
rect 142596 35332 142600 35388
rect 142536 35328 142600 35332
rect 142616 35388 142680 35392
rect 142616 35332 142620 35388
rect 142620 35332 142676 35388
rect 142676 35332 142680 35388
rect 142616 35328 142680 35332
rect 142696 35388 142760 35392
rect 142696 35332 142700 35388
rect 142700 35332 142756 35388
rect 142756 35332 142760 35388
rect 142696 35328 142760 35332
rect 173176 35388 173240 35392
rect 173176 35332 173180 35388
rect 173180 35332 173236 35388
rect 173236 35332 173240 35388
rect 173176 35328 173240 35332
rect 173256 35388 173320 35392
rect 173256 35332 173260 35388
rect 173260 35332 173316 35388
rect 173316 35332 173320 35388
rect 173256 35328 173320 35332
rect 173336 35388 173400 35392
rect 173336 35332 173340 35388
rect 173340 35332 173396 35388
rect 173396 35332 173400 35388
rect 173336 35328 173400 35332
rect 173416 35388 173480 35392
rect 173416 35332 173420 35388
rect 173420 35332 173476 35388
rect 173476 35332 173480 35388
rect 173416 35328 173480 35332
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 34936 34844 35000 34848
rect 34936 34788 34940 34844
rect 34940 34788 34996 34844
rect 34996 34788 35000 34844
rect 34936 34784 35000 34788
rect 35016 34844 35080 34848
rect 35016 34788 35020 34844
rect 35020 34788 35076 34844
rect 35076 34788 35080 34844
rect 35016 34784 35080 34788
rect 35096 34844 35160 34848
rect 35096 34788 35100 34844
rect 35100 34788 35156 34844
rect 35156 34788 35160 34844
rect 35096 34784 35160 34788
rect 35176 34844 35240 34848
rect 35176 34788 35180 34844
rect 35180 34788 35236 34844
rect 35236 34788 35240 34844
rect 35176 34784 35240 34788
rect 65656 34844 65720 34848
rect 65656 34788 65660 34844
rect 65660 34788 65716 34844
rect 65716 34788 65720 34844
rect 65656 34784 65720 34788
rect 65736 34844 65800 34848
rect 65736 34788 65740 34844
rect 65740 34788 65796 34844
rect 65796 34788 65800 34844
rect 65736 34784 65800 34788
rect 65816 34844 65880 34848
rect 65816 34788 65820 34844
rect 65820 34788 65876 34844
rect 65876 34788 65880 34844
rect 65816 34784 65880 34788
rect 65896 34844 65960 34848
rect 65896 34788 65900 34844
rect 65900 34788 65956 34844
rect 65956 34788 65960 34844
rect 65896 34784 65960 34788
rect 96376 34844 96440 34848
rect 96376 34788 96380 34844
rect 96380 34788 96436 34844
rect 96436 34788 96440 34844
rect 96376 34784 96440 34788
rect 96456 34844 96520 34848
rect 96456 34788 96460 34844
rect 96460 34788 96516 34844
rect 96516 34788 96520 34844
rect 96456 34784 96520 34788
rect 96536 34844 96600 34848
rect 96536 34788 96540 34844
rect 96540 34788 96596 34844
rect 96596 34788 96600 34844
rect 96536 34784 96600 34788
rect 96616 34844 96680 34848
rect 96616 34788 96620 34844
rect 96620 34788 96676 34844
rect 96676 34788 96680 34844
rect 96616 34784 96680 34788
rect 127096 34844 127160 34848
rect 127096 34788 127100 34844
rect 127100 34788 127156 34844
rect 127156 34788 127160 34844
rect 127096 34784 127160 34788
rect 127176 34844 127240 34848
rect 127176 34788 127180 34844
rect 127180 34788 127236 34844
rect 127236 34788 127240 34844
rect 127176 34784 127240 34788
rect 127256 34844 127320 34848
rect 127256 34788 127260 34844
rect 127260 34788 127316 34844
rect 127316 34788 127320 34844
rect 127256 34784 127320 34788
rect 127336 34844 127400 34848
rect 127336 34788 127340 34844
rect 127340 34788 127396 34844
rect 127396 34788 127400 34844
rect 127336 34784 127400 34788
rect 157816 34844 157880 34848
rect 157816 34788 157820 34844
rect 157820 34788 157876 34844
rect 157876 34788 157880 34844
rect 157816 34784 157880 34788
rect 157896 34844 157960 34848
rect 157896 34788 157900 34844
rect 157900 34788 157956 34844
rect 157956 34788 157960 34844
rect 157896 34784 157960 34788
rect 157976 34844 158040 34848
rect 157976 34788 157980 34844
rect 157980 34788 158036 34844
rect 158036 34788 158040 34844
rect 157976 34784 158040 34788
rect 158056 34844 158120 34848
rect 158056 34788 158060 34844
rect 158060 34788 158116 34844
rect 158116 34788 158120 34844
rect 158056 34784 158120 34788
rect 19576 34300 19640 34304
rect 19576 34244 19580 34300
rect 19580 34244 19636 34300
rect 19636 34244 19640 34300
rect 19576 34240 19640 34244
rect 19656 34300 19720 34304
rect 19656 34244 19660 34300
rect 19660 34244 19716 34300
rect 19716 34244 19720 34300
rect 19656 34240 19720 34244
rect 19736 34300 19800 34304
rect 19736 34244 19740 34300
rect 19740 34244 19796 34300
rect 19796 34244 19800 34300
rect 19736 34240 19800 34244
rect 19816 34300 19880 34304
rect 19816 34244 19820 34300
rect 19820 34244 19876 34300
rect 19876 34244 19880 34300
rect 19816 34240 19880 34244
rect 50296 34300 50360 34304
rect 50296 34244 50300 34300
rect 50300 34244 50356 34300
rect 50356 34244 50360 34300
rect 50296 34240 50360 34244
rect 50376 34300 50440 34304
rect 50376 34244 50380 34300
rect 50380 34244 50436 34300
rect 50436 34244 50440 34300
rect 50376 34240 50440 34244
rect 50456 34300 50520 34304
rect 50456 34244 50460 34300
rect 50460 34244 50516 34300
rect 50516 34244 50520 34300
rect 50456 34240 50520 34244
rect 50536 34300 50600 34304
rect 50536 34244 50540 34300
rect 50540 34244 50596 34300
rect 50596 34244 50600 34300
rect 50536 34240 50600 34244
rect 81016 34300 81080 34304
rect 81016 34244 81020 34300
rect 81020 34244 81076 34300
rect 81076 34244 81080 34300
rect 81016 34240 81080 34244
rect 81096 34300 81160 34304
rect 81096 34244 81100 34300
rect 81100 34244 81156 34300
rect 81156 34244 81160 34300
rect 81096 34240 81160 34244
rect 81176 34300 81240 34304
rect 81176 34244 81180 34300
rect 81180 34244 81236 34300
rect 81236 34244 81240 34300
rect 81176 34240 81240 34244
rect 81256 34300 81320 34304
rect 81256 34244 81260 34300
rect 81260 34244 81316 34300
rect 81316 34244 81320 34300
rect 81256 34240 81320 34244
rect 111736 34300 111800 34304
rect 111736 34244 111740 34300
rect 111740 34244 111796 34300
rect 111796 34244 111800 34300
rect 111736 34240 111800 34244
rect 111816 34300 111880 34304
rect 111816 34244 111820 34300
rect 111820 34244 111876 34300
rect 111876 34244 111880 34300
rect 111816 34240 111880 34244
rect 111896 34300 111960 34304
rect 111896 34244 111900 34300
rect 111900 34244 111956 34300
rect 111956 34244 111960 34300
rect 111896 34240 111960 34244
rect 111976 34300 112040 34304
rect 111976 34244 111980 34300
rect 111980 34244 112036 34300
rect 112036 34244 112040 34300
rect 111976 34240 112040 34244
rect 142456 34300 142520 34304
rect 142456 34244 142460 34300
rect 142460 34244 142516 34300
rect 142516 34244 142520 34300
rect 142456 34240 142520 34244
rect 142536 34300 142600 34304
rect 142536 34244 142540 34300
rect 142540 34244 142596 34300
rect 142596 34244 142600 34300
rect 142536 34240 142600 34244
rect 142616 34300 142680 34304
rect 142616 34244 142620 34300
rect 142620 34244 142676 34300
rect 142676 34244 142680 34300
rect 142616 34240 142680 34244
rect 142696 34300 142760 34304
rect 142696 34244 142700 34300
rect 142700 34244 142756 34300
rect 142756 34244 142760 34300
rect 142696 34240 142760 34244
rect 173176 34300 173240 34304
rect 173176 34244 173180 34300
rect 173180 34244 173236 34300
rect 173236 34244 173240 34300
rect 173176 34240 173240 34244
rect 173256 34300 173320 34304
rect 173256 34244 173260 34300
rect 173260 34244 173316 34300
rect 173316 34244 173320 34300
rect 173256 34240 173320 34244
rect 173336 34300 173400 34304
rect 173336 34244 173340 34300
rect 173340 34244 173396 34300
rect 173396 34244 173400 34300
rect 173336 34240 173400 34244
rect 173416 34300 173480 34304
rect 173416 34244 173420 34300
rect 173420 34244 173476 34300
rect 173476 34244 173480 34300
rect 173416 34240 173480 34244
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 34936 33756 35000 33760
rect 34936 33700 34940 33756
rect 34940 33700 34996 33756
rect 34996 33700 35000 33756
rect 34936 33696 35000 33700
rect 35016 33756 35080 33760
rect 35016 33700 35020 33756
rect 35020 33700 35076 33756
rect 35076 33700 35080 33756
rect 35016 33696 35080 33700
rect 35096 33756 35160 33760
rect 35096 33700 35100 33756
rect 35100 33700 35156 33756
rect 35156 33700 35160 33756
rect 35096 33696 35160 33700
rect 35176 33756 35240 33760
rect 35176 33700 35180 33756
rect 35180 33700 35236 33756
rect 35236 33700 35240 33756
rect 35176 33696 35240 33700
rect 65656 33756 65720 33760
rect 65656 33700 65660 33756
rect 65660 33700 65716 33756
rect 65716 33700 65720 33756
rect 65656 33696 65720 33700
rect 65736 33756 65800 33760
rect 65736 33700 65740 33756
rect 65740 33700 65796 33756
rect 65796 33700 65800 33756
rect 65736 33696 65800 33700
rect 65816 33756 65880 33760
rect 65816 33700 65820 33756
rect 65820 33700 65876 33756
rect 65876 33700 65880 33756
rect 65816 33696 65880 33700
rect 65896 33756 65960 33760
rect 65896 33700 65900 33756
rect 65900 33700 65956 33756
rect 65956 33700 65960 33756
rect 65896 33696 65960 33700
rect 96376 33756 96440 33760
rect 96376 33700 96380 33756
rect 96380 33700 96436 33756
rect 96436 33700 96440 33756
rect 96376 33696 96440 33700
rect 96456 33756 96520 33760
rect 96456 33700 96460 33756
rect 96460 33700 96516 33756
rect 96516 33700 96520 33756
rect 96456 33696 96520 33700
rect 96536 33756 96600 33760
rect 96536 33700 96540 33756
rect 96540 33700 96596 33756
rect 96596 33700 96600 33756
rect 96536 33696 96600 33700
rect 96616 33756 96680 33760
rect 96616 33700 96620 33756
rect 96620 33700 96676 33756
rect 96676 33700 96680 33756
rect 96616 33696 96680 33700
rect 127096 33756 127160 33760
rect 127096 33700 127100 33756
rect 127100 33700 127156 33756
rect 127156 33700 127160 33756
rect 127096 33696 127160 33700
rect 127176 33756 127240 33760
rect 127176 33700 127180 33756
rect 127180 33700 127236 33756
rect 127236 33700 127240 33756
rect 127176 33696 127240 33700
rect 127256 33756 127320 33760
rect 127256 33700 127260 33756
rect 127260 33700 127316 33756
rect 127316 33700 127320 33756
rect 127256 33696 127320 33700
rect 127336 33756 127400 33760
rect 127336 33700 127340 33756
rect 127340 33700 127396 33756
rect 127396 33700 127400 33756
rect 127336 33696 127400 33700
rect 157816 33756 157880 33760
rect 157816 33700 157820 33756
rect 157820 33700 157876 33756
rect 157876 33700 157880 33756
rect 157816 33696 157880 33700
rect 157896 33756 157960 33760
rect 157896 33700 157900 33756
rect 157900 33700 157956 33756
rect 157956 33700 157960 33756
rect 157896 33696 157960 33700
rect 157976 33756 158040 33760
rect 157976 33700 157980 33756
rect 157980 33700 158036 33756
rect 158036 33700 158040 33756
rect 157976 33696 158040 33700
rect 158056 33756 158120 33760
rect 158056 33700 158060 33756
rect 158060 33700 158116 33756
rect 158116 33700 158120 33756
rect 158056 33696 158120 33700
rect 19576 33212 19640 33216
rect 19576 33156 19580 33212
rect 19580 33156 19636 33212
rect 19636 33156 19640 33212
rect 19576 33152 19640 33156
rect 19656 33212 19720 33216
rect 19656 33156 19660 33212
rect 19660 33156 19716 33212
rect 19716 33156 19720 33212
rect 19656 33152 19720 33156
rect 19736 33212 19800 33216
rect 19736 33156 19740 33212
rect 19740 33156 19796 33212
rect 19796 33156 19800 33212
rect 19736 33152 19800 33156
rect 19816 33212 19880 33216
rect 19816 33156 19820 33212
rect 19820 33156 19876 33212
rect 19876 33156 19880 33212
rect 19816 33152 19880 33156
rect 50296 33212 50360 33216
rect 50296 33156 50300 33212
rect 50300 33156 50356 33212
rect 50356 33156 50360 33212
rect 50296 33152 50360 33156
rect 50376 33212 50440 33216
rect 50376 33156 50380 33212
rect 50380 33156 50436 33212
rect 50436 33156 50440 33212
rect 50376 33152 50440 33156
rect 50456 33212 50520 33216
rect 50456 33156 50460 33212
rect 50460 33156 50516 33212
rect 50516 33156 50520 33212
rect 50456 33152 50520 33156
rect 50536 33212 50600 33216
rect 50536 33156 50540 33212
rect 50540 33156 50596 33212
rect 50596 33156 50600 33212
rect 50536 33152 50600 33156
rect 81016 33212 81080 33216
rect 81016 33156 81020 33212
rect 81020 33156 81076 33212
rect 81076 33156 81080 33212
rect 81016 33152 81080 33156
rect 81096 33212 81160 33216
rect 81096 33156 81100 33212
rect 81100 33156 81156 33212
rect 81156 33156 81160 33212
rect 81096 33152 81160 33156
rect 81176 33212 81240 33216
rect 81176 33156 81180 33212
rect 81180 33156 81236 33212
rect 81236 33156 81240 33212
rect 81176 33152 81240 33156
rect 81256 33212 81320 33216
rect 81256 33156 81260 33212
rect 81260 33156 81316 33212
rect 81316 33156 81320 33212
rect 81256 33152 81320 33156
rect 111736 33212 111800 33216
rect 111736 33156 111740 33212
rect 111740 33156 111796 33212
rect 111796 33156 111800 33212
rect 111736 33152 111800 33156
rect 111816 33212 111880 33216
rect 111816 33156 111820 33212
rect 111820 33156 111876 33212
rect 111876 33156 111880 33212
rect 111816 33152 111880 33156
rect 111896 33212 111960 33216
rect 111896 33156 111900 33212
rect 111900 33156 111956 33212
rect 111956 33156 111960 33212
rect 111896 33152 111960 33156
rect 111976 33212 112040 33216
rect 111976 33156 111980 33212
rect 111980 33156 112036 33212
rect 112036 33156 112040 33212
rect 111976 33152 112040 33156
rect 142456 33212 142520 33216
rect 142456 33156 142460 33212
rect 142460 33156 142516 33212
rect 142516 33156 142520 33212
rect 142456 33152 142520 33156
rect 142536 33212 142600 33216
rect 142536 33156 142540 33212
rect 142540 33156 142596 33212
rect 142596 33156 142600 33212
rect 142536 33152 142600 33156
rect 142616 33212 142680 33216
rect 142616 33156 142620 33212
rect 142620 33156 142676 33212
rect 142676 33156 142680 33212
rect 142616 33152 142680 33156
rect 142696 33212 142760 33216
rect 142696 33156 142700 33212
rect 142700 33156 142756 33212
rect 142756 33156 142760 33212
rect 142696 33152 142760 33156
rect 173176 33212 173240 33216
rect 173176 33156 173180 33212
rect 173180 33156 173236 33212
rect 173236 33156 173240 33212
rect 173176 33152 173240 33156
rect 173256 33212 173320 33216
rect 173256 33156 173260 33212
rect 173260 33156 173316 33212
rect 173316 33156 173320 33212
rect 173256 33152 173320 33156
rect 173336 33212 173400 33216
rect 173336 33156 173340 33212
rect 173340 33156 173396 33212
rect 173396 33156 173400 33212
rect 173336 33152 173400 33156
rect 173416 33212 173480 33216
rect 173416 33156 173420 33212
rect 173420 33156 173476 33212
rect 173476 33156 173480 33212
rect 173416 33152 173480 33156
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 34936 32668 35000 32672
rect 34936 32612 34940 32668
rect 34940 32612 34996 32668
rect 34996 32612 35000 32668
rect 34936 32608 35000 32612
rect 35016 32668 35080 32672
rect 35016 32612 35020 32668
rect 35020 32612 35076 32668
rect 35076 32612 35080 32668
rect 35016 32608 35080 32612
rect 35096 32668 35160 32672
rect 35096 32612 35100 32668
rect 35100 32612 35156 32668
rect 35156 32612 35160 32668
rect 35096 32608 35160 32612
rect 35176 32668 35240 32672
rect 35176 32612 35180 32668
rect 35180 32612 35236 32668
rect 35236 32612 35240 32668
rect 35176 32608 35240 32612
rect 65656 32668 65720 32672
rect 65656 32612 65660 32668
rect 65660 32612 65716 32668
rect 65716 32612 65720 32668
rect 65656 32608 65720 32612
rect 65736 32668 65800 32672
rect 65736 32612 65740 32668
rect 65740 32612 65796 32668
rect 65796 32612 65800 32668
rect 65736 32608 65800 32612
rect 65816 32668 65880 32672
rect 65816 32612 65820 32668
rect 65820 32612 65876 32668
rect 65876 32612 65880 32668
rect 65816 32608 65880 32612
rect 65896 32668 65960 32672
rect 65896 32612 65900 32668
rect 65900 32612 65956 32668
rect 65956 32612 65960 32668
rect 65896 32608 65960 32612
rect 96376 32668 96440 32672
rect 96376 32612 96380 32668
rect 96380 32612 96436 32668
rect 96436 32612 96440 32668
rect 96376 32608 96440 32612
rect 96456 32668 96520 32672
rect 96456 32612 96460 32668
rect 96460 32612 96516 32668
rect 96516 32612 96520 32668
rect 96456 32608 96520 32612
rect 96536 32668 96600 32672
rect 96536 32612 96540 32668
rect 96540 32612 96596 32668
rect 96596 32612 96600 32668
rect 96536 32608 96600 32612
rect 96616 32668 96680 32672
rect 96616 32612 96620 32668
rect 96620 32612 96676 32668
rect 96676 32612 96680 32668
rect 96616 32608 96680 32612
rect 127096 32668 127160 32672
rect 127096 32612 127100 32668
rect 127100 32612 127156 32668
rect 127156 32612 127160 32668
rect 127096 32608 127160 32612
rect 127176 32668 127240 32672
rect 127176 32612 127180 32668
rect 127180 32612 127236 32668
rect 127236 32612 127240 32668
rect 127176 32608 127240 32612
rect 127256 32668 127320 32672
rect 127256 32612 127260 32668
rect 127260 32612 127316 32668
rect 127316 32612 127320 32668
rect 127256 32608 127320 32612
rect 127336 32668 127400 32672
rect 127336 32612 127340 32668
rect 127340 32612 127396 32668
rect 127396 32612 127400 32668
rect 127336 32608 127400 32612
rect 157816 32668 157880 32672
rect 157816 32612 157820 32668
rect 157820 32612 157876 32668
rect 157876 32612 157880 32668
rect 157816 32608 157880 32612
rect 157896 32668 157960 32672
rect 157896 32612 157900 32668
rect 157900 32612 157956 32668
rect 157956 32612 157960 32668
rect 157896 32608 157960 32612
rect 157976 32668 158040 32672
rect 157976 32612 157980 32668
rect 157980 32612 158036 32668
rect 158036 32612 158040 32668
rect 157976 32608 158040 32612
rect 158056 32668 158120 32672
rect 158056 32612 158060 32668
rect 158060 32612 158116 32668
rect 158116 32612 158120 32668
rect 158056 32608 158120 32612
rect 19576 32124 19640 32128
rect 19576 32068 19580 32124
rect 19580 32068 19636 32124
rect 19636 32068 19640 32124
rect 19576 32064 19640 32068
rect 19656 32124 19720 32128
rect 19656 32068 19660 32124
rect 19660 32068 19716 32124
rect 19716 32068 19720 32124
rect 19656 32064 19720 32068
rect 19736 32124 19800 32128
rect 19736 32068 19740 32124
rect 19740 32068 19796 32124
rect 19796 32068 19800 32124
rect 19736 32064 19800 32068
rect 19816 32124 19880 32128
rect 19816 32068 19820 32124
rect 19820 32068 19876 32124
rect 19876 32068 19880 32124
rect 19816 32064 19880 32068
rect 50296 32124 50360 32128
rect 50296 32068 50300 32124
rect 50300 32068 50356 32124
rect 50356 32068 50360 32124
rect 50296 32064 50360 32068
rect 50376 32124 50440 32128
rect 50376 32068 50380 32124
rect 50380 32068 50436 32124
rect 50436 32068 50440 32124
rect 50376 32064 50440 32068
rect 50456 32124 50520 32128
rect 50456 32068 50460 32124
rect 50460 32068 50516 32124
rect 50516 32068 50520 32124
rect 50456 32064 50520 32068
rect 50536 32124 50600 32128
rect 50536 32068 50540 32124
rect 50540 32068 50596 32124
rect 50596 32068 50600 32124
rect 50536 32064 50600 32068
rect 81016 32124 81080 32128
rect 81016 32068 81020 32124
rect 81020 32068 81076 32124
rect 81076 32068 81080 32124
rect 81016 32064 81080 32068
rect 81096 32124 81160 32128
rect 81096 32068 81100 32124
rect 81100 32068 81156 32124
rect 81156 32068 81160 32124
rect 81096 32064 81160 32068
rect 81176 32124 81240 32128
rect 81176 32068 81180 32124
rect 81180 32068 81236 32124
rect 81236 32068 81240 32124
rect 81176 32064 81240 32068
rect 81256 32124 81320 32128
rect 81256 32068 81260 32124
rect 81260 32068 81316 32124
rect 81316 32068 81320 32124
rect 81256 32064 81320 32068
rect 111736 32124 111800 32128
rect 111736 32068 111740 32124
rect 111740 32068 111796 32124
rect 111796 32068 111800 32124
rect 111736 32064 111800 32068
rect 111816 32124 111880 32128
rect 111816 32068 111820 32124
rect 111820 32068 111876 32124
rect 111876 32068 111880 32124
rect 111816 32064 111880 32068
rect 111896 32124 111960 32128
rect 111896 32068 111900 32124
rect 111900 32068 111956 32124
rect 111956 32068 111960 32124
rect 111896 32064 111960 32068
rect 111976 32124 112040 32128
rect 111976 32068 111980 32124
rect 111980 32068 112036 32124
rect 112036 32068 112040 32124
rect 111976 32064 112040 32068
rect 142456 32124 142520 32128
rect 142456 32068 142460 32124
rect 142460 32068 142516 32124
rect 142516 32068 142520 32124
rect 142456 32064 142520 32068
rect 142536 32124 142600 32128
rect 142536 32068 142540 32124
rect 142540 32068 142596 32124
rect 142596 32068 142600 32124
rect 142536 32064 142600 32068
rect 142616 32124 142680 32128
rect 142616 32068 142620 32124
rect 142620 32068 142676 32124
rect 142676 32068 142680 32124
rect 142616 32064 142680 32068
rect 142696 32124 142760 32128
rect 142696 32068 142700 32124
rect 142700 32068 142756 32124
rect 142756 32068 142760 32124
rect 142696 32064 142760 32068
rect 173176 32124 173240 32128
rect 173176 32068 173180 32124
rect 173180 32068 173236 32124
rect 173236 32068 173240 32124
rect 173176 32064 173240 32068
rect 173256 32124 173320 32128
rect 173256 32068 173260 32124
rect 173260 32068 173316 32124
rect 173316 32068 173320 32124
rect 173256 32064 173320 32068
rect 173336 32124 173400 32128
rect 173336 32068 173340 32124
rect 173340 32068 173396 32124
rect 173396 32068 173400 32124
rect 173336 32064 173400 32068
rect 173416 32124 173480 32128
rect 173416 32068 173420 32124
rect 173420 32068 173476 32124
rect 173476 32068 173480 32124
rect 173416 32064 173480 32068
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 34936 31580 35000 31584
rect 34936 31524 34940 31580
rect 34940 31524 34996 31580
rect 34996 31524 35000 31580
rect 34936 31520 35000 31524
rect 35016 31580 35080 31584
rect 35016 31524 35020 31580
rect 35020 31524 35076 31580
rect 35076 31524 35080 31580
rect 35016 31520 35080 31524
rect 35096 31580 35160 31584
rect 35096 31524 35100 31580
rect 35100 31524 35156 31580
rect 35156 31524 35160 31580
rect 35096 31520 35160 31524
rect 35176 31580 35240 31584
rect 35176 31524 35180 31580
rect 35180 31524 35236 31580
rect 35236 31524 35240 31580
rect 35176 31520 35240 31524
rect 65656 31580 65720 31584
rect 65656 31524 65660 31580
rect 65660 31524 65716 31580
rect 65716 31524 65720 31580
rect 65656 31520 65720 31524
rect 65736 31580 65800 31584
rect 65736 31524 65740 31580
rect 65740 31524 65796 31580
rect 65796 31524 65800 31580
rect 65736 31520 65800 31524
rect 65816 31580 65880 31584
rect 65816 31524 65820 31580
rect 65820 31524 65876 31580
rect 65876 31524 65880 31580
rect 65816 31520 65880 31524
rect 65896 31580 65960 31584
rect 65896 31524 65900 31580
rect 65900 31524 65956 31580
rect 65956 31524 65960 31580
rect 65896 31520 65960 31524
rect 96376 31580 96440 31584
rect 96376 31524 96380 31580
rect 96380 31524 96436 31580
rect 96436 31524 96440 31580
rect 96376 31520 96440 31524
rect 96456 31580 96520 31584
rect 96456 31524 96460 31580
rect 96460 31524 96516 31580
rect 96516 31524 96520 31580
rect 96456 31520 96520 31524
rect 96536 31580 96600 31584
rect 96536 31524 96540 31580
rect 96540 31524 96596 31580
rect 96596 31524 96600 31580
rect 96536 31520 96600 31524
rect 96616 31580 96680 31584
rect 96616 31524 96620 31580
rect 96620 31524 96676 31580
rect 96676 31524 96680 31580
rect 96616 31520 96680 31524
rect 127096 31580 127160 31584
rect 127096 31524 127100 31580
rect 127100 31524 127156 31580
rect 127156 31524 127160 31580
rect 127096 31520 127160 31524
rect 127176 31580 127240 31584
rect 127176 31524 127180 31580
rect 127180 31524 127236 31580
rect 127236 31524 127240 31580
rect 127176 31520 127240 31524
rect 127256 31580 127320 31584
rect 127256 31524 127260 31580
rect 127260 31524 127316 31580
rect 127316 31524 127320 31580
rect 127256 31520 127320 31524
rect 127336 31580 127400 31584
rect 127336 31524 127340 31580
rect 127340 31524 127396 31580
rect 127396 31524 127400 31580
rect 127336 31520 127400 31524
rect 157816 31580 157880 31584
rect 157816 31524 157820 31580
rect 157820 31524 157876 31580
rect 157876 31524 157880 31580
rect 157816 31520 157880 31524
rect 157896 31580 157960 31584
rect 157896 31524 157900 31580
rect 157900 31524 157956 31580
rect 157956 31524 157960 31580
rect 157896 31520 157960 31524
rect 157976 31580 158040 31584
rect 157976 31524 157980 31580
rect 157980 31524 158036 31580
rect 158036 31524 158040 31580
rect 157976 31520 158040 31524
rect 158056 31580 158120 31584
rect 158056 31524 158060 31580
rect 158060 31524 158116 31580
rect 158116 31524 158120 31580
rect 158056 31520 158120 31524
rect 19576 31036 19640 31040
rect 19576 30980 19580 31036
rect 19580 30980 19636 31036
rect 19636 30980 19640 31036
rect 19576 30976 19640 30980
rect 19656 31036 19720 31040
rect 19656 30980 19660 31036
rect 19660 30980 19716 31036
rect 19716 30980 19720 31036
rect 19656 30976 19720 30980
rect 19736 31036 19800 31040
rect 19736 30980 19740 31036
rect 19740 30980 19796 31036
rect 19796 30980 19800 31036
rect 19736 30976 19800 30980
rect 19816 31036 19880 31040
rect 19816 30980 19820 31036
rect 19820 30980 19876 31036
rect 19876 30980 19880 31036
rect 19816 30976 19880 30980
rect 50296 31036 50360 31040
rect 50296 30980 50300 31036
rect 50300 30980 50356 31036
rect 50356 30980 50360 31036
rect 50296 30976 50360 30980
rect 50376 31036 50440 31040
rect 50376 30980 50380 31036
rect 50380 30980 50436 31036
rect 50436 30980 50440 31036
rect 50376 30976 50440 30980
rect 50456 31036 50520 31040
rect 50456 30980 50460 31036
rect 50460 30980 50516 31036
rect 50516 30980 50520 31036
rect 50456 30976 50520 30980
rect 50536 31036 50600 31040
rect 50536 30980 50540 31036
rect 50540 30980 50596 31036
rect 50596 30980 50600 31036
rect 50536 30976 50600 30980
rect 81016 31036 81080 31040
rect 81016 30980 81020 31036
rect 81020 30980 81076 31036
rect 81076 30980 81080 31036
rect 81016 30976 81080 30980
rect 81096 31036 81160 31040
rect 81096 30980 81100 31036
rect 81100 30980 81156 31036
rect 81156 30980 81160 31036
rect 81096 30976 81160 30980
rect 81176 31036 81240 31040
rect 81176 30980 81180 31036
rect 81180 30980 81236 31036
rect 81236 30980 81240 31036
rect 81176 30976 81240 30980
rect 81256 31036 81320 31040
rect 81256 30980 81260 31036
rect 81260 30980 81316 31036
rect 81316 30980 81320 31036
rect 81256 30976 81320 30980
rect 111736 31036 111800 31040
rect 111736 30980 111740 31036
rect 111740 30980 111796 31036
rect 111796 30980 111800 31036
rect 111736 30976 111800 30980
rect 111816 31036 111880 31040
rect 111816 30980 111820 31036
rect 111820 30980 111876 31036
rect 111876 30980 111880 31036
rect 111816 30976 111880 30980
rect 111896 31036 111960 31040
rect 111896 30980 111900 31036
rect 111900 30980 111956 31036
rect 111956 30980 111960 31036
rect 111896 30976 111960 30980
rect 111976 31036 112040 31040
rect 111976 30980 111980 31036
rect 111980 30980 112036 31036
rect 112036 30980 112040 31036
rect 111976 30976 112040 30980
rect 142456 31036 142520 31040
rect 142456 30980 142460 31036
rect 142460 30980 142516 31036
rect 142516 30980 142520 31036
rect 142456 30976 142520 30980
rect 142536 31036 142600 31040
rect 142536 30980 142540 31036
rect 142540 30980 142596 31036
rect 142596 30980 142600 31036
rect 142536 30976 142600 30980
rect 142616 31036 142680 31040
rect 142616 30980 142620 31036
rect 142620 30980 142676 31036
rect 142676 30980 142680 31036
rect 142616 30976 142680 30980
rect 142696 31036 142760 31040
rect 142696 30980 142700 31036
rect 142700 30980 142756 31036
rect 142756 30980 142760 31036
rect 142696 30976 142760 30980
rect 173176 31036 173240 31040
rect 173176 30980 173180 31036
rect 173180 30980 173236 31036
rect 173236 30980 173240 31036
rect 173176 30976 173240 30980
rect 173256 31036 173320 31040
rect 173256 30980 173260 31036
rect 173260 30980 173316 31036
rect 173316 30980 173320 31036
rect 173256 30976 173320 30980
rect 173336 31036 173400 31040
rect 173336 30980 173340 31036
rect 173340 30980 173396 31036
rect 173396 30980 173400 31036
rect 173336 30976 173400 30980
rect 173416 31036 173480 31040
rect 173416 30980 173420 31036
rect 173420 30980 173476 31036
rect 173476 30980 173480 31036
rect 173416 30976 173480 30980
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 34936 30492 35000 30496
rect 34936 30436 34940 30492
rect 34940 30436 34996 30492
rect 34996 30436 35000 30492
rect 34936 30432 35000 30436
rect 35016 30492 35080 30496
rect 35016 30436 35020 30492
rect 35020 30436 35076 30492
rect 35076 30436 35080 30492
rect 35016 30432 35080 30436
rect 35096 30492 35160 30496
rect 35096 30436 35100 30492
rect 35100 30436 35156 30492
rect 35156 30436 35160 30492
rect 35096 30432 35160 30436
rect 35176 30492 35240 30496
rect 35176 30436 35180 30492
rect 35180 30436 35236 30492
rect 35236 30436 35240 30492
rect 35176 30432 35240 30436
rect 65656 30492 65720 30496
rect 65656 30436 65660 30492
rect 65660 30436 65716 30492
rect 65716 30436 65720 30492
rect 65656 30432 65720 30436
rect 65736 30492 65800 30496
rect 65736 30436 65740 30492
rect 65740 30436 65796 30492
rect 65796 30436 65800 30492
rect 65736 30432 65800 30436
rect 65816 30492 65880 30496
rect 65816 30436 65820 30492
rect 65820 30436 65876 30492
rect 65876 30436 65880 30492
rect 65816 30432 65880 30436
rect 65896 30492 65960 30496
rect 65896 30436 65900 30492
rect 65900 30436 65956 30492
rect 65956 30436 65960 30492
rect 65896 30432 65960 30436
rect 96376 30492 96440 30496
rect 96376 30436 96380 30492
rect 96380 30436 96436 30492
rect 96436 30436 96440 30492
rect 96376 30432 96440 30436
rect 96456 30492 96520 30496
rect 96456 30436 96460 30492
rect 96460 30436 96516 30492
rect 96516 30436 96520 30492
rect 96456 30432 96520 30436
rect 96536 30492 96600 30496
rect 96536 30436 96540 30492
rect 96540 30436 96596 30492
rect 96596 30436 96600 30492
rect 96536 30432 96600 30436
rect 96616 30492 96680 30496
rect 96616 30436 96620 30492
rect 96620 30436 96676 30492
rect 96676 30436 96680 30492
rect 96616 30432 96680 30436
rect 127096 30492 127160 30496
rect 127096 30436 127100 30492
rect 127100 30436 127156 30492
rect 127156 30436 127160 30492
rect 127096 30432 127160 30436
rect 127176 30492 127240 30496
rect 127176 30436 127180 30492
rect 127180 30436 127236 30492
rect 127236 30436 127240 30492
rect 127176 30432 127240 30436
rect 127256 30492 127320 30496
rect 127256 30436 127260 30492
rect 127260 30436 127316 30492
rect 127316 30436 127320 30492
rect 127256 30432 127320 30436
rect 127336 30492 127400 30496
rect 127336 30436 127340 30492
rect 127340 30436 127396 30492
rect 127396 30436 127400 30492
rect 127336 30432 127400 30436
rect 157816 30492 157880 30496
rect 157816 30436 157820 30492
rect 157820 30436 157876 30492
rect 157876 30436 157880 30492
rect 157816 30432 157880 30436
rect 157896 30492 157960 30496
rect 157896 30436 157900 30492
rect 157900 30436 157956 30492
rect 157956 30436 157960 30492
rect 157896 30432 157960 30436
rect 157976 30492 158040 30496
rect 157976 30436 157980 30492
rect 157980 30436 158036 30492
rect 158036 30436 158040 30492
rect 157976 30432 158040 30436
rect 158056 30492 158120 30496
rect 158056 30436 158060 30492
rect 158060 30436 158116 30492
rect 158116 30436 158120 30492
rect 158056 30432 158120 30436
rect 19576 29948 19640 29952
rect 19576 29892 19580 29948
rect 19580 29892 19636 29948
rect 19636 29892 19640 29948
rect 19576 29888 19640 29892
rect 19656 29948 19720 29952
rect 19656 29892 19660 29948
rect 19660 29892 19716 29948
rect 19716 29892 19720 29948
rect 19656 29888 19720 29892
rect 19736 29948 19800 29952
rect 19736 29892 19740 29948
rect 19740 29892 19796 29948
rect 19796 29892 19800 29948
rect 19736 29888 19800 29892
rect 19816 29948 19880 29952
rect 19816 29892 19820 29948
rect 19820 29892 19876 29948
rect 19876 29892 19880 29948
rect 19816 29888 19880 29892
rect 50296 29948 50360 29952
rect 50296 29892 50300 29948
rect 50300 29892 50356 29948
rect 50356 29892 50360 29948
rect 50296 29888 50360 29892
rect 50376 29948 50440 29952
rect 50376 29892 50380 29948
rect 50380 29892 50436 29948
rect 50436 29892 50440 29948
rect 50376 29888 50440 29892
rect 50456 29948 50520 29952
rect 50456 29892 50460 29948
rect 50460 29892 50516 29948
rect 50516 29892 50520 29948
rect 50456 29888 50520 29892
rect 50536 29948 50600 29952
rect 50536 29892 50540 29948
rect 50540 29892 50596 29948
rect 50596 29892 50600 29948
rect 50536 29888 50600 29892
rect 81016 29948 81080 29952
rect 81016 29892 81020 29948
rect 81020 29892 81076 29948
rect 81076 29892 81080 29948
rect 81016 29888 81080 29892
rect 81096 29948 81160 29952
rect 81096 29892 81100 29948
rect 81100 29892 81156 29948
rect 81156 29892 81160 29948
rect 81096 29888 81160 29892
rect 81176 29948 81240 29952
rect 81176 29892 81180 29948
rect 81180 29892 81236 29948
rect 81236 29892 81240 29948
rect 81176 29888 81240 29892
rect 81256 29948 81320 29952
rect 81256 29892 81260 29948
rect 81260 29892 81316 29948
rect 81316 29892 81320 29948
rect 81256 29888 81320 29892
rect 111736 29948 111800 29952
rect 111736 29892 111740 29948
rect 111740 29892 111796 29948
rect 111796 29892 111800 29948
rect 111736 29888 111800 29892
rect 111816 29948 111880 29952
rect 111816 29892 111820 29948
rect 111820 29892 111876 29948
rect 111876 29892 111880 29948
rect 111816 29888 111880 29892
rect 111896 29948 111960 29952
rect 111896 29892 111900 29948
rect 111900 29892 111956 29948
rect 111956 29892 111960 29948
rect 111896 29888 111960 29892
rect 111976 29948 112040 29952
rect 111976 29892 111980 29948
rect 111980 29892 112036 29948
rect 112036 29892 112040 29948
rect 111976 29888 112040 29892
rect 142456 29948 142520 29952
rect 142456 29892 142460 29948
rect 142460 29892 142516 29948
rect 142516 29892 142520 29948
rect 142456 29888 142520 29892
rect 142536 29948 142600 29952
rect 142536 29892 142540 29948
rect 142540 29892 142596 29948
rect 142596 29892 142600 29948
rect 142536 29888 142600 29892
rect 142616 29948 142680 29952
rect 142616 29892 142620 29948
rect 142620 29892 142676 29948
rect 142676 29892 142680 29948
rect 142616 29888 142680 29892
rect 142696 29948 142760 29952
rect 142696 29892 142700 29948
rect 142700 29892 142756 29948
rect 142756 29892 142760 29948
rect 142696 29888 142760 29892
rect 173176 29948 173240 29952
rect 173176 29892 173180 29948
rect 173180 29892 173236 29948
rect 173236 29892 173240 29948
rect 173176 29888 173240 29892
rect 173256 29948 173320 29952
rect 173256 29892 173260 29948
rect 173260 29892 173316 29948
rect 173316 29892 173320 29948
rect 173256 29888 173320 29892
rect 173336 29948 173400 29952
rect 173336 29892 173340 29948
rect 173340 29892 173396 29948
rect 173396 29892 173400 29948
rect 173336 29888 173400 29892
rect 173416 29948 173480 29952
rect 173416 29892 173420 29948
rect 173420 29892 173476 29948
rect 173476 29892 173480 29948
rect 173416 29888 173480 29892
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 34936 29404 35000 29408
rect 34936 29348 34940 29404
rect 34940 29348 34996 29404
rect 34996 29348 35000 29404
rect 34936 29344 35000 29348
rect 35016 29404 35080 29408
rect 35016 29348 35020 29404
rect 35020 29348 35076 29404
rect 35076 29348 35080 29404
rect 35016 29344 35080 29348
rect 35096 29404 35160 29408
rect 35096 29348 35100 29404
rect 35100 29348 35156 29404
rect 35156 29348 35160 29404
rect 35096 29344 35160 29348
rect 35176 29404 35240 29408
rect 35176 29348 35180 29404
rect 35180 29348 35236 29404
rect 35236 29348 35240 29404
rect 35176 29344 35240 29348
rect 65656 29404 65720 29408
rect 65656 29348 65660 29404
rect 65660 29348 65716 29404
rect 65716 29348 65720 29404
rect 65656 29344 65720 29348
rect 65736 29404 65800 29408
rect 65736 29348 65740 29404
rect 65740 29348 65796 29404
rect 65796 29348 65800 29404
rect 65736 29344 65800 29348
rect 65816 29404 65880 29408
rect 65816 29348 65820 29404
rect 65820 29348 65876 29404
rect 65876 29348 65880 29404
rect 65816 29344 65880 29348
rect 65896 29404 65960 29408
rect 65896 29348 65900 29404
rect 65900 29348 65956 29404
rect 65956 29348 65960 29404
rect 65896 29344 65960 29348
rect 96376 29404 96440 29408
rect 96376 29348 96380 29404
rect 96380 29348 96436 29404
rect 96436 29348 96440 29404
rect 96376 29344 96440 29348
rect 96456 29404 96520 29408
rect 96456 29348 96460 29404
rect 96460 29348 96516 29404
rect 96516 29348 96520 29404
rect 96456 29344 96520 29348
rect 96536 29404 96600 29408
rect 96536 29348 96540 29404
rect 96540 29348 96596 29404
rect 96596 29348 96600 29404
rect 96536 29344 96600 29348
rect 96616 29404 96680 29408
rect 96616 29348 96620 29404
rect 96620 29348 96676 29404
rect 96676 29348 96680 29404
rect 96616 29344 96680 29348
rect 127096 29404 127160 29408
rect 127096 29348 127100 29404
rect 127100 29348 127156 29404
rect 127156 29348 127160 29404
rect 127096 29344 127160 29348
rect 127176 29404 127240 29408
rect 127176 29348 127180 29404
rect 127180 29348 127236 29404
rect 127236 29348 127240 29404
rect 127176 29344 127240 29348
rect 127256 29404 127320 29408
rect 127256 29348 127260 29404
rect 127260 29348 127316 29404
rect 127316 29348 127320 29404
rect 127256 29344 127320 29348
rect 127336 29404 127400 29408
rect 127336 29348 127340 29404
rect 127340 29348 127396 29404
rect 127396 29348 127400 29404
rect 127336 29344 127400 29348
rect 157816 29404 157880 29408
rect 157816 29348 157820 29404
rect 157820 29348 157876 29404
rect 157876 29348 157880 29404
rect 157816 29344 157880 29348
rect 157896 29404 157960 29408
rect 157896 29348 157900 29404
rect 157900 29348 157956 29404
rect 157956 29348 157960 29404
rect 157896 29344 157960 29348
rect 157976 29404 158040 29408
rect 157976 29348 157980 29404
rect 157980 29348 158036 29404
rect 158036 29348 158040 29404
rect 157976 29344 158040 29348
rect 158056 29404 158120 29408
rect 158056 29348 158060 29404
rect 158060 29348 158116 29404
rect 158116 29348 158120 29404
rect 158056 29344 158120 29348
rect 19576 28860 19640 28864
rect 19576 28804 19580 28860
rect 19580 28804 19636 28860
rect 19636 28804 19640 28860
rect 19576 28800 19640 28804
rect 19656 28860 19720 28864
rect 19656 28804 19660 28860
rect 19660 28804 19716 28860
rect 19716 28804 19720 28860
rect 19656 28800 19720 28804
rect 19736 28860 19800 28864
rect 19736 28804 19740 28860
rect 19740 28804 19796 28860
rect 19796 28804 19800 28860
rect 19736 28800 19800 28804
rect 19816 28860 19880 28864
rect 19816 28804 19820 28860
rect 19820 28804 19876 28860
rect 19876 28804 19880 28860
rect 19816 28800 19880 28804
rect 50296 28860 50360 28864
rect 50296 28804 50300 28860
rect 50300 28804 50356 28860
rect 50356 28804 50360 28860
rect 50296 28800 50360 28804
rect 50376 28860 50440 28864
rect 50376 28804 50380 28860
rect 50380 28804 50436 28860
rect 50436 28804 50440 28860
rect 50376 28800 50440 28804
rect 50456 28860 50520 28864
rect 50456 28804 50460 28860
rect 50460 28804 50516 28860
rect 50516 28804 50520 28860
rect 50456 28800 50520 28804
rect 50536 28860 50600 28864
rect 50536 28804 50540 28860
rect 50540 28804 50596 28860
rect 50596 28804 50600 28860
rect 50536 28800 50600 28804
rect 81016 28860 81080 28864
rect 81016 28804 81020 28860
rect 81020 28804 81076 28860
rect 81076 28804 81080 28860
rect 81016 28800 81080 28804
rect 81096 28860 81160 28864
rect 81096 28804 81100 28860
rect 81100 28804 81156 28860
rect 81156 28804 81160 28860
rect 81096 28800 81160 28804
rect 81176 28860 81240 28864
rect 81176 28804 81180 28860
rect 81180 28804 81236 28860
rect 81236 28804 81240 28860
rect 81176 28800 81240 28804
rect 81256 28860 81320 28864
rect 81256 28804 81260 28860
rect 81260 28804 81316 28860
rect 81316 28804 81320 28860
rect 81256 28800 81320 28804
rect 111736 28860 111800 28864
rect 111736 28804 111740 28860
rect 111740 28804 111796 28860
rect 111796 28804 111800 28860
rect 111736 28800 111800 28804
rect 111816 28860 111880 28864
rect 111816 28804 111820 28860
rect 111820 28804 111876 28860
rect 111876 28804 111880 28860
rect 111816 28800 111880 28804
rect 111896 28860 111960 28864
rect 111896 28804 111900 28860
rect 111900 28804 111956 28860
rect 111956 28804 111960 28860
rect 111896 28800 111960 28804
rect 111976 28860 112040 28864
rect 111976 28804 111980 28860
rect 111980 28804 112036 28860
rect 112036 28804 112040 28860
rect 111976 28800 112040 28804
rect 142456 28860 142520 28864
rect 142456 28804 142460 28860
rect 142460 28804 142516 28860
rect 142516 28804 142520 28860
rect 142456 28800 142520 28804
rect 142536 28860 142600 28864
rect 142536 28804 142540 28860
rect 142540 28804 142596 28860
rect 142596 28804 142600 28860
rect 142536 28800 142600 28804
rect 142616 28860 142680 28864
rect 142616 28804 142620 28860
rect 142620 28804 142676 28860
rect 142676 28804 142680 28860
rect 142616 28800 142680 28804
rect 142696 28860 142760 28864
rect 142696 28804 142700 28860
rect 142700 28804 142756 28860
rect 142756 28804 142760 28860
rect 142696 28800 142760 28804
rect 173176 28860 173240 28864
rect 173176 28804 173180 28860
rect 173180 28804 173236 28860
rect 173236 28804 173240 28860
rect 173176 28800 173240 28804
rect 173256 28860 173320 28864
rect 173256 28804 173260 28860
rect 173260 28804 173316 28860
rect 173316 28804 173320 28860
rect 173256 28800 173320 28804
rect 173336 28860 173400 28864
rect 173336 28804 173340 28860
rect 173340 28804 173396 28860
rect 173396 28804 173400 28860
rect 173336 28800 173400 28804
rect 173416 28860 173480 28864
rect 173416 28804 173420 28860
rect 173420 28804 173476 28860
rect 173476 28804 173480 28860
rect 173416 28800 173480 28804
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 34936 28316 35000 28320
rect 34936 28260 34940 28316
rect 34940 28260 34996 28316
rect 34996 28260 35000 28316
rect 34936 28256 35000 28260
rect 35016 28316 35080 28320
rect 35016 28260 35020 28316
rect 35020 28260 35076 28316
rect 35076 28260 35080 28316
rect 35016 28256 35080 28260
rect 35096 28316 35160 28320
rect 35096 28260 35100 28316
rect 35100 28260 35156 28316
rect 35156 28260 35160 28316
rect 35096 28256 35160 28260
rect 35176 28316 35240 28320
rect 35176 28260 35180 28316
rect 35180 28260 35236 28316
rect 35236 28260 35240 28316
rect 35176 28256 35240 28260
rect 65656 28316 65720 28320
rect 65656 28260 65660 28316
rect 65660 28260 65716 28316
rect 65716 28260 65720 28316
rect 65656 28256 65720 28260
rect 65736 28316 65800 28320
rect 65736 28260 65740 28316
rect 65740 28260 65796 28316
rect 65796 28260 65800 28316
rect 65736 28256 65800 28260
rect 65816 28316 65880 28320
rect 65816 28260 65820 28316
rect 65820 28260 65876 28316
rect 65876 28260 65880 28316
rect 65816 28256 65880 28260
rect 65896 28316 65960 28320
rect 65896 28260 65900 28316
rect 65900 28260 65956 28316
rect 65956 28260 65960 28316
rect 65896 28256 65960 28260
rect 96376 28316 96440 28320
rect 96376 28260 96380 28316
rect 96380 28260 96436 28316
rect 96436 28260 96440 28316
rect 96376 28256 96440 28260
rect 96456 28316 96520 28320
rect 96456 28260 96460 28316
rect 96460 28260 96516 28316
rect 96516 28260 96520 28316
rect 96456 28256 96520 28260
rect 96536 28316 96600 28320
rect 96536 28260 96540 28316
rect 96540 28260 96596 28316
rect 96596 28260 96600 28316
rect 96536 28256 96600 28260
rect 96616 28316 96680 28320
rect 96616 28260 96620 28316
rect 96620 28260 96676 28316
rect 96676 28260 96680 28316
rect 96616 28256 96680 28260
rect 127096 28316 127160 28320
rect 127096 28260 127100 28316
rect 127100 28260 127156 28316
rect 127156 28260 127160 28316
rect 127096 28256 127160 28260
rect 127176 28316 127240 28320
rect 127176 28260 127180 28316
rect 127180 28260 127236 28316
rect 127236 28260 127240 28316
rect 127176 28256 127240 28260
rect 127256 28316 127320 28320
rect 127256 28260 127260 28316
rect 127260 28260 127316 28316
rect 127316 28260 127320 28316
rect 127256 28256 127320 28260
rect 127336 28316 127400 28320
rect 127336 28260 127340 28316
rect 127340 28260 127396 28316
rect 127396 28260 127400 28316
rect 127336 28256 127400 28260
rect 157816 28316 157880 28320
rect 157816 28260 157820 28316
rect 157820 28260 157876 28316
rect 157876 28260 157880 28316
rect 157816 28256 157880 28260
rect 157896 28316 157960 28320
rect 157896 28260 157900 28316
rect 157900 28260 157956 28316
rect 157956 28260 157960 28316
rect 157896 28256 157960 28260
rect 157976 28316 158040 28320
rect 157976 28260 157980 28316
rect 157980 28260 158036 28316
rect 158036 28260 158040 28316
rect 157976 28256 158040 28260
rect 158056 28316 158120 28320
rect 158056 28260 158060 28316
rect 158060 28260 158116 28316
rect 158116 28260 158120 28316
rect 158056 28256 158120 28260
rect 19576 27772 19640 27776
rect 19576 27716 19580 27772
rect 19580 27716 19636 27772
rect 19636 27716 19640 27772
rect 19576 27712 19640 27716
rect 19656 27772 19720 27776
rect 19656 27716 19660 27772
rect 19660 27716 19716 27772
rect 19716 27716 19720 27772
rect 19656 27712 19720 27716
rect 19736 27772 19800 27776
rect 19736 27716 19740 27772
rect 19740 27716 19796 27772
rect 19796 27716 19800 27772
rect 19736 27712 19800 27716
rect 19816 27772 19880 27776
rect 19816 27716 19820 27772
rect 19820 27716 19876 27772
rect 19876 27716 19880 27772
rect 19816 27712 19880 27716
rect 50296 27772 50360 27776
rect 50296 27716 50300 27772
rect 50300 27716 50356 27772
rect 50356 27716 50360 27772
rect 50296 27712 50360 27716
rect 50376 27772 50440 27776
rect 50376 27716 50380 27772
rect 50380 27716 50436 27772
rect 50436 27716 50440 27772
rect 50376 27712 50440 27716
rect 50456 27772 50520 27776
rect 50456 27716 50460 27772
rect 50460 27716 50516 27772
rect 50516 27716 50520 27772
rect 50456 27712 50520 27716
rect 50536 27772 50600 27776
rect 50536 27716 50540 27772
rect 50540 27716 50596 27772
rect 50596 27716 50600 27772
rect 50536 27712 50600 27716
rect 81016 27772 81080 27776
rect 81016 27716 81020 27772
rect 81020 27716 81076 27772
rect 81076 27716 81080 27772
rect 81016 27712 81080 27716
rect 81096 27772 81160 27776
rect 81096 27716 81100 27772
rect 81100 27716 81156 27772
rect 81156 27716 81160 27772
rect 81096 27712 81160 27716
rect 81176 27772 81240 27776
rect 81176 27716 81180 27772
rect 81180 27716 81236 27772
rect 81236 27716 81240 27772
rect 81176 27712 81240 27716
rect 81256 27772 81320 27776
rect 81256 27716 81260 27772
rect 81260 27716 81316 27772
rect 81316 27716 81320 27772
rect 81256 27712 81320 27716
rect 111736 27772 111800 27776
rect 111736 27716 111740 27772
rect 111740 27716 111796 27772
rect 111796 27716 111800 27772
rect 111736 27712 111800 27716
rect 111816 27772 111880 27776
rect 111816 27716 111820 27772
rect 111820 27716 111876 27772
rect 111876 27716 111880 27772
rect 111816 27712 111880 27716
rect 111896 27772 111960 27776
rect 111896 27716 111900 27772
rect 111900 27716 111956 27772
rect 111956 27716 111960 27772
rect 111896 27712 111960 27716
rect 111976 27772 112040 27776
rect 111976 27716 111980 27772
rect 111980 27716 112036 27772
rect 112036 27716 112040 27772
rect 111976 27712 112040 27716
rect 142456 27772 142520 27776
rect 142456 27716 142460 27772
rect 142460 27716 142516 27772
rect 142516 27716 142520 27772
rect 142456 27712 142520 27716
rect 142536 27772 142600 27776
rect 142536 27716 142540 27772
rect 142540 27716 142596 27772
rect 142596 27716 142600 27772
rect 142536 27712 142600 27716
rect 142616 27772 142680 27776
rect 142616 27716 142620 27772
rect 142620 27716 142676 27772
rect 142676 27716 142680 27772
rect 142616 27712 142680 27716
rect 142696 27772 142760 27776
rect 142696 27716 142700 27772
rect 142700 27716 142756 27772
rect 142756 27716 142760 27772
rect 142696 27712 142760 27716
rect 173176 27772 173240 27776
rect 173176 27716 173180 27772
rect 173180 27716 173236 27772
rect 173236 27716 173240 27772
rect 173176 27712 173240 27716
rect 173256 27772 173320 27776
rect 173256 27716 173260 27772
rect 173260 27716 173316 27772
rect 173316 27716 173320 27772
rect 173256 27712 173320 27716
rect 173336 27772 173400 27776
rect 173336 27716 173340 27772
rect 173340 27716 173396 27772
rect 173396 27716 173400 27772
rect 173336 27712 173400 27716
rect 173416 27772 173480 27776
rect 173416 27716 173420 27772
rect 173420 27716 173476 27772
rect 173476 27716 173480 27772
rect 173416 27712 173480 27716
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 34936 27228 35000 27232
rect 34936 27172 34940 27228
rect 34940 27172 34996 27228
rect 34996 27172 35000 27228
rect 34936 27168 35000 27172
rect 35016 27228 35080 27232
rect 35016 27172 35020 27228
rect 35020 27172 35076 27228
rect 35076 27172 35080 27228
rect 35016 27168 35080 27172
rect 35096 27228 35160 27232
rect 35096 27172 35100 27228
rect 35100 27172 35156 27228
rect 35156 27172 35160 27228
rect 35096 27168 35160 27172
rect 35176 27228 35240 27232
rect 35176 27172 35180 27228
rect 35180 27172 35236 27228
rect 35236 27172 35240 27228
rect 35176 27168 35240 27172
rect 65656 27228 65720 27232
rect 65656 27172 65660 27228
rect 65660 27172 65716 27228
rect 65716 27172 65720 27228
rect 65656 27168 65720 27172
rect 65736 27228 65800 27232
rect 65736 27172 65740 27228
rect 65740 27172 65796 27228
rect 65796 27172 65800 27228
rect 65736 27168 65800 27172
rect 65816 27228 65880 27232
rect 65816 27172 65820 27228
rect 65820 27172 65876 27228
rect 65876 27172 65880 27228
rect 65816 27168 65880 27172
rect 65896 27228 65960 27232
rect 65896 27172 65900 27228
rect 65900 27172 65956 27228
rect 65956 27172 65960 27228
rect 65896 27168 65960 27172
rect 96376 27228 96440 27232
rect 96376 27172 96380 27228
rect 96380 27172 96436 27228
rect 96436 27172 96440 27228
rect 96376 27168 96440 27172
rect 96456 27228 96520 27232
rect 96456 27172 96460 27228
rect 96460 27172 96516 27228
rect 96516 27172 96520 27228
rect 96456 27168 96520 27172
rect 96536 27228 96600 27232
rect 96536 27172 96540 27228
rect 96540 27172 96596 27228
rect 96596 27172 96600 27228
rect 96536 27168 96600 27172
rect 96616 27228 96680 27232
rect 96616 27172 96620 27228
rect 96620 27172 96676 27228
rect 96676 27172 96680 27228
rect 96616 27168 96680 27172
rect 127096 27228 127160 27232
rect 127096 27172 127100 27228
rect 127100 27172 127156 27228
rect 127156 27172 127160 27228
rect 127096 27168 127160 27172
rect 127176 27228 127240 27232
rect 127176 27172 127180 27228
rect 127180 27172 127236 27228
rect 127236 27172 127240 27228
rect 127176 27168 127240 27172
rect 127256 27228 127320 27232
rect 127256 27172 127260 27228
rect 127260 27172 127316 27228
rect 127316 27172 127320 27228
rect 127256 27168 127320 27172
rect 127336 27228 127400 27232
rect 127336 27172 127340 27228
rect 127340 27172 127396 27228
rect 127396 27172 127400 27228
rect 127336 27168 127400 27172
rect 157816 27228 157880 27232
rect 157816 27172 157820 27228
rect 157820 27172 157876 27228
rect 157876 27172 157880 27228
rect 157816 27168 157880 27172
rect 157896 27228 157960 27232
rect 157896 27172 157900 27228
rect 157900 27172 157956 27228
rect 157956 27172 157960 27228
rect 157896 27168 157960 27172
rect 157976 27228 158040 27232
rect 157976 27172 157980 27228
rect 157980 27172 158036 27228
rect 158036 27172 158040 27228
rect 157976 27168 158040 27172
rect 158056 27228 158120 27232
rect 158056 27172 158060 27228
rect 158060 27172 158116 27228
rect 158116 27172 158120 27228
rect 158056 27168 158120 27172
rect 19576 26684 19640 26688
rect 19576 26628 19580 26684
rect 19580 26628 19636 26684
rect 19636 26628 19640 26684
rect 19576 26624 19640 26628
rect 19656 26684 19720 26688
rect 19656 26628 19660 26684
rect 19660 26628 19716 26684
rect 19716 26628 19720 26684
rect 19656 26624 19720 26628
rect 19736 26684 19800 26688
rect 19736 26628 19740 26684
rect 19740 26628 19796 26684
rect 19796 26628 19800 26684
rect 19736 26624 19800 26628
rect 19816 26684 19880 26688
rect 19816 26628 19820 26684
rect 19820 26628 19876 26684
rect 19876 26628 19880 26684
rect 19816 26624 19880 26628
rect 50296 26684 50360 26688
rect 50296 26628 50300 26684
rect 50300 26628 50356 26684
rect 50356 26628 50360 26684
rect 50296 26624 50360 26628
rect 50376 26684 50440 26688
rect 50376 26628 50380 26684
rect 50380 26628 50436 26684
rect 50436 26628 50440 26684
rect 50376 26624 50440 26628
rect 50456 26684 50520 26688
rect 50456 26628 50460 26684
rect 50460 26628 50516 26684
rect 50516 26628 50520 26684
rect 50456 26624 50520 26628
rect 50536 26684 50600 26688
rect 50536 26628 50540 26684
rect 50540 26628 50596 26684
rect 50596 26628 50600 26684
rect 50536 26624 50600 26628
rect 81016 26684 81080 26688
rect 81016 26628 81020 26684
rect 81020 26628 81076 26684
rect 81076 26628 81080 26684
rect 81016 26624 81080 26628
rect 81096 26684 81160 26688
rect 81096 26628 81100 26684
rect 81100 26628 81156 26684
rect 81156 26628 81160 26684
rect 81096 26624 81160 26628
rect 81176 26684 81240 26688
rect 81176 26628 81180 26684
rect 81180 26628 81236 26684
rect 81236 26628 81240 26684
rect 81176 26624 81240 26628
rect 81256 26684 81320 26688
rect 81256 26628 81260 26684
rect 81260 26628 81316 26684
rect 81316 26628 81320 26684
rect 81256 26624 81320 26628
rect 111736 26684 111800 26688
rect 111736 26628 111740 26684
rect 111740 26628 111796 26684
rect 111796 26628 111800 26684
rect 111736 26624 111800 26628
rect 111816 26684 111880 26688
rect 111816 26628 111820 26684
rect 111820 26628 111876 26684
rect 111876 26628 111880 26684
rect 111816 26624 111880 26628
rect 111896 26684 111960 26688
rect 111896 26628 111900 26684
rect 111900 26628 111956 26684
rect 111956 26628 111960 26684
rect 111896 26624 111960 26628
rect 111976 26684 112040 26688
rect 111976 26628 111980 26684
rect 111980 26628 112036 26684
rect 112036 26628 112040 26684
rect 111976 26624 112040 26628
rect 142456 26684 142520 26688
rect 142456 26628 142460 26684
rect 142460 26628 142516 26684
rect 142516 26628 142520 26684
rect 142456 26624 142520 26628
rect 142536 26684 142600 26688
rect 142536 26628 142540 26684
rect 142540 26628 142596 26684
rect 142596 26628 142600 26684
rect 142536 26624 142600 26628
rect 142616 26684 142680 26688
rect 142616 26628 142620 26684
rect 142620 26628 142676 26684
rect 142676 26628 142680 26684
rect 142616 26624 142680 26628
rect 142696 26684 142760 26688
rect 142696 26628 142700 26684
rect 142700 26628 142756 26684
rect 142756 26628 142760 26684
rect 142696 26624 142760 26628
rect 173176 26684 173240 26688
rect 173176 26628 173180 26684
rect 173180 26628 173236 26684
rect 173236 26628 173240 26684
rect 173176 26624 173240 26628
rect 173256 26684 173320 26688
rect 173256 26628 173260 26684
rect 173260 26628 173316 26684
rect 173316 26628 173320 26684
rect 173256 26624 173320 26628
rect 173336 26684 173400 26688
rect 173336 26628 173340 26684
rect 173340 26628 173396 26684
rect 173396 26628 173400 26684
rect 173336 26624 173400 26628
rect 173416 26684 173480 26688
rect 173416 26628 173420 26684
rect 173420 26628 173476 26684
rect 173476 26628 173480 26684
rect 173416 26624 173480 26628
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 34936 26140 35000 26144
rect 34936 26084 34940 26140
rect 34940 26084 34996 26140
rect 34996 26084 35000 26140
rect 34936 26080 35000 26084
rect 35016 26140 35080 26144
rect 35016 26084 35020 26140
rect 35020 26084 35076 26140
rect 35076 26084 35080 26140
rect 35016 26080 35080 26084
rect 35096 26140 35160 26144
rect 35096 26084 35100 26140
rect 35100 26084 35156 26140
rect 35156 26084 35160 26140
rect 35096 26080 35160 26084
rect 35176 26140 35240 26144
rect 35176 26084 35180 26140
rect 35180 26084 35236 26140
rect 35236 26084 35240 26140
rect 35176 26080 35240 26084
rect 65656 26140 65720 26144
rect 65656 26084 65660 26140
rect 65660 26084 65716 26140
rect 65716 26084 65720 26140
rect 65656 26080 65720 26084
rect 65736 26140 65800 26144
rect 65736 26084 65740 26140
rect 65740 26084 65796 26140
rect 65796 26084 65800 26140
rect 65736 26080 65800 26084
rect 65816 26140 65880 26144
rect 65816 26084 65820 26140
rect 65820 26084 65876 26140
rect 65876 26084 65880 26140
rect 65816 26080 65880 26084
rect 65896 26140 65960 26144
rect 65896 26084 65900 26140
rect 65900 26084 65956 26140
rect 65956 26084 65960 26140
rect 65896 26080 65960 26084
rect 96376 26140 96440 26144
rect 96376 26084 96380 26140
rect 96380 26084 96436 26140
rect 96436 26084 96440 26140
rect 96376 26080 96440 26084
rect 96456 26140 96520 26144
rect 96456 26084 96460 26140
rect 96460 26084 96516 26140
rect 96516 26084 96520 26140
rect 96456 26080 96520 26084
rect 96536 26140 96600 26144
rect 96536 26084 96540 26140
rect 96540 26084 96596 26140
rect 96596 26084 96600 26140
rect 96536 26080 96600 26084
rect 96616 26140 96680 26144
rect 96616 26084 96620 26140
rect 96620 26084 96676 26140
rect 96676 26084 96680 26140
rect 96616 26080 96680 26084
rect 127096 26140 127160 26144
rect 127096 26084 127100 26140
rect 127100 26084 127156 26140
rect 127156 26084 127160 26140
rect 127096 26080 127160 26084
rect 127176 26140 127240 26144
rect 127176 26084 127180 26140
rect 127180 26084 127236 26140
rect 127236 26084 127240 26140
rect 127176 26080 127240 26084
rect 127256 26140 127320 26144
rect 127256 26084 127260 26140
rect 127260 26084 127316 26140
rect 127316 26084 127320 26140
rect 127256 26080 127320 26084
rect 127336 26140 127400 26144
rect 127336 26084 127340 26140
rect 127340 26084 127396 26140
rect 127396 26084 127400 26140
rect 127336 26080 127400 26084
rect 157816 26140 157880 26144
rect 157816 26084 157820 26140
rect 157820 26084 157876 26140
rect 157876 26084 157880 26140
rect 157816 26080 157880 26084
rect 157896 26140 157960 26144
rect 157896 26084 157900 26140
rect 157900 26084 157956 26140
rect 157956 26084 157960 26140
rect 157896 26080 157960 26084
rect 157976 26140 158040 26144
rect 157976 26084 157980 26140
rect 157980 26084 158036 26140
rect 158036 26084 158040 26140
rect 157976 26080 158040 26084
rect 158056 26140 158120 26144
rect 158056 26084 158060 26140
rect 158060 26084 158116 26140
rect 158116 26084 158120 26140
rect 158056 26080 158120 26084
rect 19576 25596 19640 25600
rect 19576 25540 19580 25596
rect 19580 25540 19636 25596
rect 19636 25540 19640 25596
rect 19576 25536 19640 25540
rect 19656 25596 19720 25600
rect 19656 25540 19660 25596
rect 19660 25540 19716 25596
rect 19716 25540 19720 25596
rect 19656 25536 19720 25540
rect 19736 25596 19800 25600
rect 19736 25540 19740 25596
rect 19740 25540 19796 25596
rect 19796 25540 19800 25596
rect 19736 25536 19800 25540
rect 19816 25596 19880 25600
rect 19816 25540 19820 25596
rect 19820 25540 19876 25596
rect 19876 25540 19880 25596
rect 19816 25536 19880 25540
rect 50296 25596 50360 25600
rect 50296 25540 50300 25596
rect 50300 25540 50356 25596
rect 50356 25540 50360 25596
rect 50296 25536 50360 25540
rect 50376 25596 50440 25600
rect 50376 25540 50380 25596
rect 50380 25540 50436 25596
rect 50436 25540 50440 25596
rect 50376 25536 50440 25540
rect 50456 25596 50520 25600
rect 50456 25540 50460 25596
rect 50460 25540 50516 25596
rect 50516 25540 50520 25596
rect 50456 25536 50520 25540
rect 50536 25596 50600 25600
rect 50536 25540 50540 25596
rect 50540 25540 50596 25596
rect 50596 25540 50600 25596
rect 50536 25536 50600 25540
rect 81016 25596 81080 25600
rect 81016 25540 81020 25596
rect 81020 25540 81076 25596
rect 81076 25540 81080 25596
rect 81016 25536 81080 25540
rect 81096 25596 81160 25600
rect 81096 25540 81100 25596
rect 81100 25540 81156 25596
rect 81156 25540 81160 25596
rect 81096 25536 81160 25540
rect 81176 25596 81240 25600
rect 81176 25540 81180 25596
rect 81180 25540 81236 25596
rect 81236 25540 81240 25596
rect 81176 25536 81240 25540
rect 81256 25596 81320 25600
rect 81256 25540 81260 25596
rect 81260 25540 81316 25596
rect 81316 25540 81320 25596
rect 81256 25536 81320 25540
rect 111736 25596 111800 25600
rect 111736 25540 111740 25596
rect 111740 25540 111796 25596
rect 111796 25540 111800 25596
rect 111736 25536 111800 25540
rect 111816 25596 111880 25600
rect 111816 25540 111820 25596
rect 111820 25540 111876 25596
rect 111876 25540 111880 25596
rect 111816 25536 111880 25540
rect 111896 25596 111960 25600
rect 111896 25540 111900 25596
rect 111900 25540 111956 25596
rect 111956 25540 111960 25596
rect 111896 25536 111960 25540
rect 111976 25596 112040 25600
rect 111976 25540 111980 25596
rect 111980 25540 112036 25596
rect 112036 25540 112040 25596
rect 111976 25536 112040 25540
rect 142456 25596 142520 25600
rect 142456 25540 142460 25596
rect 142460 25540 142516 25596
rect 142516 25540 142520 25596
rect 142456 25536 142520 25540
rect 142536 25596 142600 25600
rect 142536 25540 142540 25596
rect 142540 25540 142596 25596
rect 142596 25540 142600 25596
rect 142536 25536 142600 25540
rect 142616 25596 142680 25600
rect 142616 25540 142620 25596
rect 142620 25540 142676 25596
rect 142676 25540 142680 25596
rect 142616 25536 142680 25540
rect 142696 25596 142760 25600
rect 142696 25540 142700 25596
rect 142700 25540 142756 25596
rect 142756 25540 142760 25596
rect 142696 25536 142760 25540
rect 173176 25596 173240 25600
rect 173176 25540 173180 25596
rect 173180 25540 173236 25596
rect 173236 25540 173240 25596
rect 173176 25536 173240 25540
rect 173256 25596 173320 25600
rect 173256 25540 173260 25596
rect 173260 25540 173316 25596
rect 173316 25540 173320 25596
rect 173256 25536 173320 25540
rect 173336 25596 173400 25600
rect 173336 25540 173340 25596
rect 173340 25540 173396 25596
rect 173396 25540 173400 25596
rect 173336 25536 173400 25540
rect 173416 25596 173480 25600
rect 173416 25540 173420 25596
rect 173420 25540 173476 25596
rect 173476 25540 173480 25596
rect 173416 25536 173480 25540
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 34936 25052 35000 25056
rect 34936 24996 34940 25052
rect 34940 24996 34996 25052
rect 34996 24996 35000 25052
rect 34936 24992 35000 24996
rect 35016 25052 35080 25056
rect 35016 24996 35020 25052
rect 35020 24996 35076 25052
rect 35076 24996 35080 25052
rect 35016 24992 35080 24996
rect 35096 25052 35160 25056
rect 35096 24996 35100 25052
rect 35100 24996 35156 25052
rect 35156 24996 35160 25052
rect 35096 24992 35160 24996
rect 35176 25052 35240 25056
rect 35176 24996 35180 25052
rect 35180 24996 35236 25052
rect 35236 24996 35240 25052
rect 35176 24992 35240 24996
rect 65656 25052 65720 25056
rect 65656 24996 65660 25052
rect 65660 24996 65716 25052
rect 65716 24996 65720 25052
rect 65656 24992 65720 24996
rect 65736 25052 65800 25056
rect 65736 24996 65740 25052
rect 65740 24996 65796 25052
rect 65796 24996 65800 25052
rect 65736 24992 65800 24996
rect 65816 25052 65880 25056
rect 65816 24996 65820 25052
rect 65820 24996 65876 25052
rect 65876 24996 65880 25052
rect 65816 24992 65880 24996
rect 65896 25052 65960 25056
rect 65896 24996 65900 25052
rect 65900 24996 65956 25052
rect 65956 24996 65960 25052
rect 65896 24992 65960 24996
rect 96376 25052 96440 25056
rect 96376 24996 96380 25052
rect 96380 24996 96436 25052
rect 96436 24996 96440 25052
rect 96376 24992 96440 24996
rect 96456 25052 96520 25056
rect 96456 24996 96460 25052
rect 96460 24996 96516 25052
rect 96516 24996 96520 25052
rect 96456 24992 96520 24996
rect 96536 25052 96600 25056
rect 96536 24996 96540 25052
rect 96540 24996 96596 25052
rect 96596 24996 96600 25052
rect 96536 24992 96600 24996
rect 96616 25052 96680 25056
rect 96616 24996 96620 25052
rect 96620 24996 96676 25052
rect 96676 24996 96680 25052
rect 96616 24992 96680 24996
rect 127096 25052 127160 25056
rect 127096 24996 127100 25052
rect 127100 24996 127156 25052
rect 127156 24996 127160 25052
rect 127096 24992 127160 24996
rect 127176 25052 127240 25056
rect 127176 24996 127180 25052
rect 127180 24996 127236 25052
rect 127236 24996 127240 25052
rect 127176 24992 127240 24996
rect 127256 25052 127320 25056
rect 127256 24996 127260 25052
rect 127260 24996 127316 25052
rect 127316 24996 127320 25052
rect 127256 24992 127320 24996
rect 127336 25052 127400 25056
rect 127336 24996 127340 25052
rect 127340 24996 127396 25052
rect 127396 24996 127400 25052
rect 127336 24992 127400 24996
rect 157816 25052 157880 25056
rect 157816 24996 157820 25052
rect 157820 24996 157876 25052
rect 157876 24996 157880 25052
rect 157816 24992 157880 24996
rect 157896 25052 157960 25056
rect 157896 24996 157900 25052
rect 157900 24996 157956 25052
rect 157956 24996 157960 25052
rect 157896 24992 157960 24996
rect 157976 25052 158040 25056
rect 157976 24996 157980 25052
rect 157980 24996 158036 25052
rect 158036 24996 158040 25052
rect 157976 24992 158040 24996
rect 158056 25052 158120 25056
rect 158056 24996 158060 25052
rect 158060 24996 158116 25052
rect 158116 24996 158120 25052
rect 158056 24992 158120 24996
rect 19576 24508 19640 24512
rect 19576 24452 19580 24508
rect 19580 24452 19636 24508
rect 19636 24452 19640 24508
rect 19576 24448 19640 24452
rect 19656 24508 19720 24512
rect 19656 24452 19660 24508
rect 19660 24452 19716 24508
rect 19716 24452 19720 24508
rect 19656 24448 19720 24452
rect 19736 24508 19800 24512
rect 19736 24452 19740 24508
rect 19740 24452 19796 24508
rect 19796 24452 19800 24508
rect 19736 24448 19800 24452
rect 19816 24508 19880 24512
rect 19816 24452 19820 24508
rect 19820 24452 19876 24508
rect 19876 24452 19880 24508
rect 19816 24448 19880 24452
rect 50296 24508 50360 24512
rect 50296 24452 50300 24508
rect 50300 24452 50356 24508
rect 50356 24452 50360 24508
rect 50296 24448 50360 24452
rect 50376 24508 50440 24512
rect 50376 24452 50380 24508
rect 50380 24452 50436 24508
rect 50436 24452 50440 24508
rect 50376 24448 50440 24452
rect 50456 24508 50520 24512
rect 50456 24452 50460 24508
rect 50460 24452 50516 24508
rect 50516 24452 50520 24508
rect 50456 24448 50520 24452
rect 50536 24508 50600 24512
rect 50536 24452 50540 24508
rect 50540 24452 50596 24508
rect 50596 24452 50600 24508
rect 50536 24448 50600 24452
rect 81016 24508 81080 24512
rect 81016 24452 81020 24508
rect 81020 24452 81076 24508
rect 81076 24452 81080 24508
rect 81016 24448 81080 24452
rect 81096 24508 81160 24512
rect 81096 24452 81100 24508
rect 81100 24452 81156 24508
rect 81156 24452 81160 24508
rect 81096 24448 81160 24452
rect 81176 24508 81240 24512
rect 81176 24452 81180 24508
rect 81180 24452 81236 24508
rect 81236 24452 81240 24508
rect 81176 24448 81240 24452
rect 81256 24508 81320 24512
rect 81256 24452 81260 24508
rect 81260 24452 81316 24508
rect 81316 24452 81320 24508
rect 81256 24448 81320 24452
rect 111736 24508 111800 24512
rect 111736 24452 111740 24508
rect 111740 24452 111796 24508
rect 111796 24452 111800 24508
rect 111736 24448 111800 24452
rect 111816 24508 111880 24512
rect 111816 24452 111820 24508
rect 111820 24452 111876 24508
rect 111876 24452 111880 24508
rect 111816 24448 111880 24452
rect 111896 24508 111960 24512
rect 111896 24452 111900 24508
rect 111900 24452 111956 24508
rect 111956 24452 111960 24508
rect 111896 24448 111960 24452
rect 111976 24508 112040 24512
rect 111976 24452 111980 24508
rect 111980 24452 112036 24508
rect 112036 24452 112040 24508
rect 111976 24448 112040 24452
rect 142456 24508 142520 24512
rect 142456 24452 142460 24508
rect 142460 24452 142516 24508
rect 142516 24452 142520 24508
rect 142456 24448 142520 24452
rect 142536 24508 142600 24512
rect 142536 24452 142540 24508
rect 142540 24452 142596 24508
rect 142596 24452 142600 24508
rect 142536 24448 142600 24452
rect 142616 24508 142680 24512
rect 142616 24452 142620 24508
rect 142620 24452 142676 24508
rect 142676 24452 142680 24508
rect 142616 24448 142680 24452
rect 142696 24508 142760 24512
rect 142696 24452 142700 24508
rect 142700 24452 142756 24508
rect 142756 24452 142760 24508
rect 142696 24448 142760 24452
rect 173176 24508 173240 24512
rect 173176 24452 173180 24508
rect 173180 24452 173236 24508
rect 173236 24452 173240 24508
rect 173176 24448 173240 24452
rect 173256 24508 173320 24512
rect 173256 24452 173260 24508
rect 173260 24452 173316 24508
rect 173316 24452 173320 24508
rect 173256 24448 173320 24452
rect 173336 24508 173400 24512
rect 173336 24452 173340 24508
rect 173340 24452 173396 24508
rect 173396 24452 173400 24508
rect 173336 24448 173400 24452
rect 173416 24508 173480 24512
rect 173416 24452 173420 24508
rect 173420 24452 173476 24508
rect 173476 24452 173480 24508
rect 173416 24448 173480 24452
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 34936 23964 35000 23968
rect 34936 23908 34940 23964
rect 34940 23908 34996 23964
rect 34996 23908 35000 23964
rect 34936 23904 35000 23908
rect 35016 23964 35080 23968
rect 35016 23908 35020 23964
rect 35020 23908 35076 23964
rect 35076 23908 35080 23964
rect 35016 23904 35080 23908
rect 35096 23964 35160 23968
rect 35096 23908 35100 23964
rect 35100 23908 35156 23964
rect 35156 23908 35160 23964
rect 35096 23904 35160 23908
rect 35176 23964 35240 23968
rect 35176 23908 35180 23964
rect 35180 23908 35236 23964
rect 35236 23908 35240 23964
rect 35176 23904 35240 23908
rect 65656 23964 65720 23968
rect 65656 23908 65660 23964
rect 65660 23908 65716 23964
rect 65716 23908 65720 23964
rect 65656 23904 65720 23908
rect 65736 23964 65800 23968
rect 65736 23908 65740 23964
rect 65740 23908 65796 23964
rect 65796 23908 65800 23964
rect 65736 23904 65800 23908
rect 65816 23964 65880 23968
rect 65816 23908 65820 23964
rect 65820 23908 65876 23964
rect 65876 23908 65880 23964
rect 65816 23904 65880 23908
rect 65896 23964 65960 23968
rect 65896 23908 65900 23964
rect 65900 23908 65956 23964
rect 65956 23908 65960 23964
rect 65896 23904 65960 23908
rect 96376 23964 96440 23968
rect 96376 23908 96380 23964
rect 96380 23908 96436 23964
rect 96436 23908 96440 23964
rect 96376 23904 96440 23908
rect 96456 23964 96520 23968
rect 96456 23908 96460 23964
rect 96460 23908 96516 23964
rect 96516 23908 96520 23964
rect 96456 23904 96520 23908
rect 96536 23964 96600 23968
rect 96536 23908 96540 23964
rect 96540 23908 96596 23964
rect 96596 23908 96600 23964
rect 96536 23904 96600 23908
rect 96616 23964 96680 23968
rect 96616 23908 96620 23964
rect 96620 23908 96676 23964
rect 96676 23908 96680 23964
rect 96616 23904 96680 23908
rect 127096 23964 127160 23968
rect 127096 23908 127100 23964
rect 127100 23908 127156 23964
rect 127156 23908 127160 23964
rect 127096 23904 127160 23908
rect 127176 23964 127240 23968
rect 127176 23908 127180 23964
rect 127180 23908 127236 23964
rect 127236 23908 127240 23964
rect 127176 23904 127240 23908
rect 127256 23964 127320 23968
rect 127256 23908 127260 23964
rect 127260 23908 127316 23964
rect 127316 23908 127320 23964
rect 127256 23904 127320 23908
rect 127336 23964 127400 23968
rect 127336 23908 127340 23964
rect 127340 23908 127396 23964
rect 127396 23908 127400 23964
rect 127336 23904 127400 23908
rect 157816 23964 157880 23968
rect 157816 23908 157820 23964
rect 157820 23908 157876 23964
rect 157876 23908 157880 23964
rect 157816 23904 157880 23908
rect 157896 23964 157960 23968
rect 157896 23908 157900 23964
rect 157900 23908 157956 23964
rect 157956 23908 157960 23964
rect 157896 23904 157960 23908
rect 157976 23964 158040 23968
rect 157976 23908 157980 23964
rect 157980 23908 158036 23964
rect 158036 23908 158040 23964
rect 157976 23904 158040 23908
rect 158056 23964 158120 23968
rect 158056 23908 158060 23964
rect 158060 23908 158116 23964
rect 158116 23908 158120 23964
rect 158056 23904 158120 23908
rect 19576 23420 19640 23424
rect 19576 23364 19580 23420
rect 19580 23364 19636 23420
rect 19636 23364 19640 23420
rect 19576 23360 19640 23364
rect 19656 23420 19720 23424
rect 19656 23364 19660 23420
rect 19660 23364 19716 23420
rect 19716 23364 19720 23420
rect 19656 23360 19720 23364
rect 19736 23420 19800 23424
rect 19736 23364 19740 23420
rect 19740 23364 19796 23420
rect 19796 23364 19800 23420
rect 19736 23360 19800 23364
rect 19816 23420 19880 23424
rect 19816 23364 19820 23420
rect 19820 23364 19876 23420
rect 19876 23364 19880 23420
rect 19816 23360 19880 23364
rect 50296 23420 50360 23424
rect 50296 23364 50300 23420
rect 50300 23364 50356 23420
rect 50356 23364 50360 23420
rect 50296 23360 50360 23364
rect 50376 23420 50440 23424
rect 50376 23364 50380 23420
rect 50380 23364 50436 23420
rect 50436 23364 50440 23420
rect 50376 23360 50440 23364
rect 50456 23420 50520 23424
rect 50456 23364 50460 23420
rect 50460 23364 50516 23420
rect 50516 23364 50520 23420
rect 50456 23360 50520 23364
rect 50536 23420 50600 23424
rect 50536 23364 50540 23420
rect 50540 23364 50596 23420
rect 50596 23364 50600 23420
rect 50536 23360 50600 23364
rect 81016 23420 81080 23424
rect 81016 23364 81020 23420
rect 81020 23364 81076 23420
rect 81076 23364 81080 23420
rect 81016 23360 81080 23364
rect 81096 23420 81160 23424
rect 81096 23364 81100 23420
rect 81100 23364 81156 23420
rect 81156 23364 81160 23420
rect 81096 23360 81160 23364
rect 81176 23420 81240 23424
rect 81176 23364 81180 23420
rect 81180 23364 81236 23420
rect 81236 23364 81240 23420
rect 81176 23360 81240 23364
rect 81256 23420 81320 23424
rect 81256 23364 81260 23420
rect 81260 23364 81316 23420
rect 81316 23364 81320 23420
rect 81256 23360 81320 23364
rect 111736 23420 111800 23424
rect 111736 23364 111740 23420
rect 111740 23364 111796 23420
rect 111796 23364 111800 23420
rect 111736 23360 111800 23364
rect 111816 23420 111880 23424
rect 111816 23364 111820 23420
rect 111820 23364 111876 23420
rect 111876 23364 111880 23420
rect 111816 23360 111880 23364
rect 111896 23420 111960 23424
rect 111896 23364 111900 23420
rect 111900 23364 111956 23420
rect 111956 23364 111960 23420
rect 111896 23360 111960 23364
rect 111976 23420 112040 23424
rect 111976 23364 111980 23420
rect 111980 23364 112036 23420
rect 112036 23364 112040 23420
rect 111976 23360 112040 23364
rect 142456 23420 142520 23424
rect 142456 23364 142460 23420
rect 142460 23364 142516 23420
rect 142516 23364 142520 23420
rect 142456 23360 142520 23364
rect 142536 23420 142600 23424
rect 142536 23364 142540 23420
rect 142540 23364 142596 23420
rect 142596 23364 142600 23420
rect 142536 23360 142600 23364
rect 142616 23420 142680 23424
rect 142616 23364 142620 23420
rect 142620 23364 142676 23420
rect 142676 23364 142680 23420
rect 142616 23360 142680 23364
rect 142696 23420 142760 23424
rect 142696 23364 142700 23420
rect 142700 23364 142756 23420
rect 142756 23364 142760 23420
rect 142696 23360 142760 23364
rect 173176 23420 173240 23424
rect 173176 23364 173180 23420
rect 173180 23364 173236 23420
rect 173236 23364 173240 23420
rect 173176 23360 173240 23364
rect 173256 23420 173320 23424
rect 173256 23364 173260 23420
rect 173260 23364 173316 23420
rect 173316 23364 173320 23420
rect 173256 23360 173320 23364
rect 173336 23420 173400 23424
rect 173336 23364 173340 23420
rect 173340 23364 173396 23420
rect 173396 23364 173400 23420
rect 173336 23360 173400 23364
rect 173416 23420 173480 23424
rect 173416 23364 173420 23420
rect 173420 23364 173476 23420
rect 173476 23364 173480 23420
rect 173416 23360 173480 23364
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 34936 22876 35000 22880
rect 34936 22820 34940 22876
rect 34940 22820 34996 22876
rect 34996 22820 35000 22876
rect 34936 22816 35000 22820
rect 35016 22876 35080 22880
rect 35016 22820 35020 22876
rect 35020 22820 35076 22876
rect 35076 22820 35080 22876
rect 35016 22816 35080 22820
rect 35096 22876 35160 22880
rect 35096 22820 35100 22876
rect 35100 22820 35156 22876
rect 35156 22820 35160 22876
rect 35096 22816 35160 22820
rect 35176 22876 35240 22880
rect 35176 22820 35180 22876
rect 35180 22820 35236 22876
rect 35236 22820 35240 22876
rect 35176 22816 35240 22820
rect 65656 22876 65720 22880
rect 65656 22820 65660 22876
rect 65660 22820 65716 22876
rect 65716 22820 65720 22876
rect 65656 22816 65720 22820
rect 65736 22876 65800 22880
rect 65736 22820 65740 22876
rect 65740 22820 65796 22876
rect 65796 22820 65800 22876
rect 65736 22816 65800 22820
rect 65816 22876 65880 22880
rect 65816 22820 65820 22876
rect 65820 22820 65876 22876
rect 65876 22820 65880 22876
rect 65816 22816 65880 22820
rect 65896 22876 65960 22880
rect 65896 22820 65900 22876
rect 65900 22820 65956 22876
rect 65956 22820 65960 22876
rect 65896 22816 65960 22820
rect 96376 22876 96440 22880
rect 96376 22820 96380 22876
rect 96380 22820 96436 22876
rect 96436 22820 96440 22876
rect 96376 22816 96440 22820
rect 96456 22876 96520 22880
rect 96456 22820 96460 22876
rect 96460 22820 96516 22876
rect 96516 22820 96520 22876
rect 96456 22816 96520 22820
rect 96536 22876 96600 22880
rect 96536 22820 96540 22876
rect 96540 22820 96596 22876
rect 96596 22820 96600 22876
rect 96536 22816 96600 22820
rect 96616 22876 96680 22880
rect 96616 22820 96620 22876
rect 96620 22820 96676 22876
rect 96676 22820 96680 22876
rect 96616 22816 96680 22820
rect 127096 22876 127160 22880
rect 127096 22820 127100 22876
rect 127100 22820 127156 22876
rect 127156 22820 127160 22876
rect 127096 22816 127160 22820
rect 127176 22876 127240 22880
rect 127176 22820 127180 22876
rect 127180 22820 127236 22876
rect 127236 22820 127240 22876
rect 127176 22816 127240 22820
rect 127256 22876 127320 22880
rect 127256 22820 127260 22876
rect 127260 22820 127316 22876
rect 127316 22820 127320 22876
rect 127256 22816 127320 22820
rect 127336 22876 127400 22880
rect 127336 22820 127340 22876
rect 127340 22820 127396 22876
rect 127396 22820 127400 22876
rect 127336 22816 127400 22820
rect 157816 22876 157880 22880
rect 157816 22820 157820 22876
rect 157820 22820 157876 22876
rect 157876 22820 157880 22876
rect 157816 22816 157880 22820
rect 157896 22876 157960 22880
rect 157896 22820 157900 22876
rect 157900 22820 157956 22876
rect 157956 22820 157960 22876
rect 157896 22816 157960 22820
rect 157976 22876 158040 22880
rect 157976 22820 157980 22876
rect 157980 22820 158036 22876
rect 158036 22820 158040 22876
rect 157976 22816 158040 22820
rect 158056 22876 158120 22880
rect 158056 22820 158060 22876
rect 158060 22820 158116 22876
rect 158116 22820 158120 22876
rect 158056 22816 158120 22820
rect 19576 22332 19640 22336
rect 19576 22276 19580 22332
rect 19580 22276 19636 22332
rect 19636 22276 19640 22332
rect 19576 22272 19640 22276
rect 19656 22332 19720 22336
rect 19656 22276 19660 22332
rect 19660 22276 19716 22332
rect 19716 22276 19720 22332
rect 19656 22272 19720 22276
rect 19736 22332 19800 22336
rect 19736 22276 19740 22332
rect 19740 22276 19796 22332
rect 19796 22276 19800 22332
rect 19736 22272 19800 22276
rect 19816 22332 19880 22336
rect 19816 22276 19820 22332
rect 19820 22276 19876 22332
rect 19876 22276 19880 22332
rect 19816 22272 19880 22276
rect 50296 22332 50360 22336
rect 50296 22276 50300 22332
rect 50300 22276 50356 22332
rect 50356 22276 50360 22332
rect 50296 22272 50360 22276
rect 50376 22332 50440 22336
rect 50376 22276 50380 22332
rect 50380 22276 50436 22332
rect 50436 22276 50440 22332
rect 50376 22272 50440 22276
rect 50456 22332 50520 22336
rect 50456 22276 50460 22332
rect 50460 22276 50516 22332
rect 50516 22276 50520 22332
rect 50456 22272 50520 22276
rect 50536 22332 50600 22336
rect 50536 22276 50540 22332
rect 50540 22276 50596 22332
rect 50596 22276 50600 22332
rect 50536 22272 50600 22276
rect 81016 22332 81080 22336
rect 81016 22276 81020 22332
rect 81020 22276 81076 22332
rect 81076 22276 81080 22332
rect 81016 22272 81080 22276
rect 81096 22332 81160 22336
rect 81096 22276 81100 22332
rect 81100 22276 81156 22332
rect 81156 22276 81160 22332
rect 81096 22272 81160 22276
rect 81176 22332 81240 22336
rect 81176 22276 81180 22332
rect 81180 22276 81236 22332
rect 81236 22276 81240 22332
rect 81176 22272 81240 22276
rect 81256 22332 81320 22336
rect 81256 22276 81260 22332
rect 81260 22276 81316 22332
rect 81316 22276 81320 22332
rect 81256 22272 81320 22276
rect 111736 22332 111800 22336
rect 111736 22276 111740 22332
rect 111740 22276 111796 22332
rect 111796 22276 111800 22332
rect 111736 22272 111800 22276
rect 111816 22332 111880 22336
rect 111816 22276 111820 22332
rect 111820 22276 111876 22332
rect 111876 22276 111880 22332
rect 111816 22272 111880 22276
rect 111896 22332 111960 22336
rect 111896 22276 111900 22332
rect 111900 22276 111956 22332
rect 111956 22276 111960 22332
rect 111896 22272 111960 22276
rect 111976 22332 112040 22336
rect 111976 22276 111980 22332
rect 111980 22276 112036 22332
rect 112036 22276 112040 22332
rect 111976 22272 112040 22276
rect 142456 22332 142520 22336
rect 142456 22276 142460 22332
rect 142460 22276 142516 22332
rect 142516 22276 142520 22332
rect 142456 22272 142520 22276
rect 142536 22332 142600 22336
rect 142536 22276 142540 22332
rect 142540 22276 142596 22332
rect 142596 22276 142600 22332
rect 142536 22272 142600 22276
rect 142616 22332 142680 22336
rect 142616 22276 142620 22332
rect 142620 22276 142676 22332
rect 142676 22276 142680 22332
rect 142616 22272 142680 22276
rect 142696 22332 142760 22336
rect 142696 22276 142700 22332
rect 142700 22276 142756 22332
rect 142756 22276 142760 22332
rect 142696 22272 142760 22276
rect 173176 22332 173240 22336
rect 173176 22276 173180 22332
rect 173180 22276 173236 22332
rect 173236 22276 173240 22332
rect 173176 22272 173240 22276
rect 173256 22332 173320 22336
rect 173256 22276 173260 22332
rect 173260 22276 173316 22332
rect 173316 22276 173320 22332
rect 173256 22272 173320 22276
rect 173336 22332 173400 22336
rect 173336 22276 173340 22332
rect 173340 22276 173396 22332
rect 173396 22276 173400 22332
rect 173336 22272 173400 22276
rect 173416 22332 173480 22336
rect 173416 22276 173420 22332
rect 173420 22276 173476 22332
rect 173476 22276 173480 22332
rect 173416 22272 173480 22276
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 34936 21788 35000 21792
rect 34936 21732 34940 21788
rect 34940 21732 34996 21788
rect 34996 21732 35000 21788
rect 34936 21728 35000 21732
rect 35016 21788 35080 21792
rect 35016 21732 35020 21788
rect 35020 21732 35076 21788
rect 35076 21732 35080 21788
rect 35016 21728 35080 21732
rect 35096 21788 35160 21792
rect 35096 21732 35100 21788
rect 35100 21732 35156 21788
rect 35156 21732 35160 21788
rect 35096 21728 35160 21732
rect 35176 21788 35240 21792
rect 35176 21732 35180 21788
rect 35180 21732 35236 21788
rect 35236 21732 35240 21788
rect 35176 21728 35240 21732
rect 65656 21788 65720 21792
rect 65656 21732 65660 21788
rect 65660 21732 65716 21788
rect 65716 21732 65720 21788
rect 65656 21728 65720 21732
rect 65736 21788 65800 21792
rect 65736 21732 65740 21788
rect 65740 21732 65796 21788
rect 65796 21732 65800 21788
rect 65736 21728 65800 21732
rect 65816 21788 65880 21792
rect 65816 21732 65820 21788
rect 65820 21732 65876 21788
rect 65876 21732 65880 21788
rect 65816 21728 65880 21732
rect 65896 21788 65960 21792
rect 65896 21732 65900 21788
rect 65900 21732 65956 21788
rect 65956 21732 65960 21788
rect 65896 21728 65960 21732
rect 96376 21788 96440 21792
rect 96376 21732 96380 21788
rect 96380 21732 96436 21788
rect 96436 21732 96440 21788
rect 96376 21728 96440 21732
rect 96456 21788 96520 21792
rect 96456 21732 96460 21788
rect 96460 21732 96516 21788
rect 96516 21732 96520 21788
rect 96456 21728 96520 21732
rect 96536 21788 96600 21792
rect 96536 21732 96540 21788
rect 96540 21732 96596 21788
rect 96596 21732 96600 21788
rect 96536 21728 96600 21732
rect 96616 21788 96680 21792
rect 96616 21732 96620 21788
rect 96620 21732 96676 21788
rect 96676 21732 96680 21788
rect 96616 21728 96680 21732
rect 127096 21788 127160 21792
rect 127096 21732 127100 21788
rect 127100 21732 127156 21788
rect 127156 21732 127160 21788
rect 127096 21728 127160 21732
rect 127176 21788 127240 21792
rect 127176 21732 127180 21788
rect 127180 21732 127236 21788
rect 127236 21732 127240 21788
rect 127176 21728 127240 21732
rect 127256 21788 127320 21792
rect 127256 21732 127260 21788
rect 127260 21732 127316 21788
rect 127316 21732 127320 21788
rect 127256 21728 127320 21732
rect 127336 21788 127400 21792
rect 127336 21732 127340 21788
rect 127340 21732 127396 21788
rect 127396 21732 127400 21788
rect 127336 21728 127400 21732
rect 157816 21788 157880 21792
rect 157816 21732 157820 21788
rect 157820 21732 157876 21788
rect 157876 21732 157880 21788
rect 157816 21728 157880 21732
rect 157896 21788 157960 21792
rect 157896 21732 157900 21788
rect 157900 21732 157956 21788
rect 157956 21732 157960 21788
rect 157896 21728 157960 21732
rect 157976 21788 158040 21792
rect 157976 21732 157980 21788
rect 157980 21732 158036 21788
rect 158036 21732 158040 21788
rect 157976 21728 158040 21732
rect 158056 21788 158120 21792
rect 158056 21732 158060 21788
rect 158060 21732 158116 21788
rect 158116 21732 158120 21788
rect 158056 21728 158120 21732
rect 19576 21244 19640 21248
rect 19576 21188 19580 21244
rect 19580 21188 19636 21244
rect 19636 21188 19640 21244
rect 19576 21184 19640 21188
rect 19656 21244 19720 21248
rect 19656 21188 19660 21244
rect 19660 21188 19716 21244
rect 19716 21188 19720 21244
rect 19656 21184 19720 21188
rect 19736 21244 19800 21248
rect 19736 21188 19740 21244
rect 19740 21188 19796 21244
rect 19796 21188 19800 21244
rect 19736 21184 19800 21188
rect 19816 21244 19880 21248
rect 19816 21188 19820 21244
rect 19820 21188 19876 21244
rect 19876 21188 19880 21244
rect 19816 21184 19880 21188
rect 50296 21244 50360 21248
rect 50296 21188 50300 21244
rect 50300 21188 50356 21244
rect 50356 21188 50360 21244
rect 50296 21184 50360 21188
rect 50376 21244 50440 21248
rect 50376 21188 50380 21244
rect 50380 21188 50436 21244
rect 50436 21188 50440 21244
rect 50376 21184 50440 21188
rect 50456 21244 50520 21248
rect 50456 21188 50460 21244
rect 50460 21188 50516 21244
rect 50516 21188 50520 21244
rect 50456 21184 50520 21188
rect 50536 21244 50600 21248
rect 50536 21188 50540 21244
rect 50540 21188 50596 21244
rect 50596 21188 50600 21244
rect 50536 21184 50600 21188
rect 81016 21244 81080 21248
rect 81016 21188 81020 21244
rect 81020 21188 81076 21244
rect 81076 21188 81080 21244
rect 81016 21184 81080 21188
rect 81096 21244 81160 21248
rect 81096 21188 81100 21244
rect 81100 21188 81156 21244
rect 81156 21188 81160 21244
rect 81096 21184 81160 21188
rect 81176 21244 81240 21248
rect 81176 21188 81180 21244
rect 81180 21188 81236 21244
rect 81236 21188 81240 21244
rect 81176 21184 81240 21188
rect 81256 21244 81320 21248
rect 81256 21188 81260 21244
rect 81260 21188 81316 21244
rect 81316 21188 81320 21244
rect 81256 21184 81320 21188
rect 111736 21244 111800 21248
rect 111736 21188 111740 21244
rect 111740 21188 111796 21244
rect 111796 21188 111800 21244
rect 111736 21184 111800 21188
rect 111816 21244 111880 21248
rect 111816 21188 111820 21244
rect 111820 21188 111876 21244
rect 111876 21188 111880 21244
rect 111816 21184 111880 21188
rect 111896 21244 111960 21248
rect 111896 21188 111900 21244
rect 111900 21188 111956 21244
rect 111956 21188 111960 21244
rect 111896 21184 111960 21188
rect 111976 21244 112040 21248
rect 111976 21188 111980 21244
rect 111980 21188 112036 21244
rect 112036 21188 112040 21244
rect 111976 21184 112040 21188
rect 142456 21244 142520 21248
rect 142456 21188 142460 21244
rect 142460 21188 142516 21244
rect 142516 21188 142520 21244
rect 142456 21184 142520 21188
rect 142536 21244 142600 21248
rect 142536 21188 142540 21244
rect 142540 21188 142596 21244
rect 142596 21188 142600 21244
rect 142536 21184 142600 21188
rect 142616 21244 142680 21248
rect 142616 21188 142620 21244
rect 142620 21188 142676 21244
rect 142676 21188 142680 21244
rect 142616 21184 142680 21188
rect 142696 21244 142760 21248
rect 142696 21188 142700 21244
rect 142700 21188 142756 21244
rect 142756 21188 142760 21244
rect 142696 21184 142760 21188
rect 173176 21244 173240 21248
rect 173176 21188 173180 21244
rect 173180 21188 173236 21244
rect 173236 21188 173240 21244
rect 173176 21184 173240 21188
rect 173256 21244 173320 21248
rect 173256 21188 173260 21244
rect 173260 21188 173316 21244
rect 173316 21188 173320 21244
rect 173256 21184 173320 21188
rect 173336 21244 173400 21248
rect 173336 21188 173340 21244
rect 173340 21188 173396 21244
rect 173396 21188 173400 21244
rect 173336 21184 173400 21188
rect 173416 21244 173480 21248
rect 173416 21188 173420 21244
rect 173420 21188 173476 21244
rect 173476 21188 173480 21244
rect 173416 21184 173480 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 34936 20700 35000 20704
rect 34936 20644 34940 20700
rect 34940 20644 34996 20700
rect 34996 20644 35000 20700
rect 34936 20640 35000 20644
rect 35016 20700 35080 20704
rect 35016 20644 35020 20700
rect 35020 20644 35076 20700
rect 35076 20644 35080 20700
rect 35016 20640 35080 20644
rect 35096 20700 35160 20704
rect 35096 20644 35100 20700
rect 35100 20644 35156 20700
rect 35156 20644 35160 20700
rect 35096 20640 35160 20644
rect 35176 20700 35240 20704
rect 35176 20644 35180 20700
rect 35180 20644 35236 20700
rect 35236 20644 35240 20700
rect 35176 20640 35240 20644
rect 65656 20700 65720 20704
rect 65656 20644 65660 20700
rect 65660 20644 65716 20700
rect 65716 20644 65720 20700
rect 65656 20640 65720 20644
rect 65736 20700 65800 20704
rect 65736 20644 65740 20700
rect 65740 20644 65796 20700
rect 65796 20644 65800 20700
rect 65736 20640 65800 20644
rect 65816 20700 65880 20704
rect 65816 20644 65820 20700
rect 65820 20644 65876 20700
rect 65876 20644 65880 20700
rect 65816 20640 65880 20644
rect 65896 20700 65960 20704
rect 65896 20644 65900 20700
rect 65900 20644 65956 20700
rect 65956 20644 65960 20700
rect 65896 20640 65960 20644
rect 96376 20700 96440 20704
rect 96376 20644 96380 20700
rect 96380 20644 96436 20700
rect 96436 20644 96440 20700
rect 96376 20640 96440 20644
rect 96456 20700 96520 20704
rect 96456 20644 96460 20700
rect 96460 20644 96516 20700
rect 96516 20644 96520 20700
rect 96456 20640 96520 20644
rect 96536 20700 96600 20704
rect 96536 20644 96540 20700
rect 96540 20644 96596 20700
rect 96596 20644 96600 20700
rect 96536 20640 96600 20644
rect 96616 20700 96680 20704
rect 96616 20644 96620 20700
rect 96620 20644 96676 20700
rect 96676 20644 96680 20700
rect 96616 20640 96680 20644
rect 127096 20700 127160 20704
rect 127096 20644 127100 20700
rect 127100 20644 127156 20700
rect 127156 20644 127160 20700
rect 127096 20640 127160 20644
rect 127176 20700 127240 20704
rect 127176 20644 127180 20700
rect 127180 20644 127236 20700
rect 127236 20644 127240 20700
rect 127176 20640 127240 20644
rect 127256 20700 127320 20704
rect 127256 20644 127260 20700
rect 127260 20644 127316 20700
rect 127316 20644 127320 20700
rect 127256 20640 127320 20644
rect 127336 20700 127400 20704
rect 127336 20644 127340 20700
rect 127340 20644 127396 20700
rect 127396 20644 127400 20700
rect 127336 20640 127400 20644
rect 157816 20700 157880 20704
rect 157816 20644 157820 20700
rect 157820 20644 157876 20700
rect 157876 20644 157880 20700
rect 157816 20640 157880 20644
rect 157896 20700 157960 20704
rect 157896 20644 157900 20700
rect 157900 20644 157956 20700
rect 157956 20644 157960 20700
rect 157896 20640 157960 20644
rect 157976 20700 158040 20704
rect 157976 20644 157980 20700
rect 157980 20644 158036 20700
rect 158036 20644 158040 20700
rect 157976 20640 158040 20644
rect 158056 20700 158120 20704
rect 158056 20644 158060 20700
rect 158060 20644 158116 20700
rect 158116 20644 158120 20700
rect 158056 20640 158120 20644
rect 19576 20156 19640 20160
rect 19576 20100 19580 20156
rect 19580 20100 19636 20156
rect 19636 20100 19640 20156
rect 19576 20096 19640 20100
rect 19656 20156 19720 20160
rect 19656 20100 19660 20156
rect 19660 20100 19716 20156
rect 19716 20100 19720 20156
rect 19656 20096 19720 20100
rect 19736 20156 19800 20160
rect 19736 20100 19740 20156
rect 19740 20100 19796 20156
rect 19796 20100 19800 20156
rect 19736 20096 19800 20100
rect 19816 20156 19880 20160
rect 19816 20100 19820 20156
rect 19820 20100 19876 20156
rect 19876 20100 19880 20156
rect 19816 20096 19880 20100
rect 50296 20156 50360 20160
rect 50296 20100 50300 20156
rect 50300 20100 50356 20156
rect 50356 20100 50360 20156
rect 50296 20096 50360 20100
rect 50376 20156 50440 20160
rect 50376 20100 50380 20156
rect 50380 20100 50436 20156
rect 50436 20100 50440 20156
rect 50376 20096 50440 20100
rect 50456 20156 50520 20160
rect 50456 20100 50460 20156
rect 50460 20100 50516 20156
rect 50516 20100 50520 20156
rect 50456 20096 50520 20100
rect 50536 20156 50600 20160
rect 50536 20100 50540 20156
rect 50540 20100 50596 20156
rect 50596 20100 50600 20156
rect 50536 20096 50600 20100
rect 81016 20156 81080 20160
rect 81016 20100 81020 20156
rect 81020 20100 81076 20156
rect 81076 20100 81080 20156
rect 81016 20096 81080 20100
rect 81096 20156 81160 20160
rect 81096 20100 81100 20156
rect 81100 20100 81156 20156
rect 81156 20100 81160 20156
rect 81096 20096 81160 20100
rect 81176 20156 81240 20160
rect 81176 20100 81180 20156
rect 81180 20100 81236 20156
rect 81236 20100 81240 20156
rect 81176 20096 81240 20100
rect 81256 20156 81320 20160
rect 81256 20100 81260 20156
rect 81260 20100 81316 20156
rect 81316 20100 81320 20156
rect 81256 20096 81320 20100
rect 111736 20156 111800 20160
rect 111736 20100 111740 20156
rect 111740 20100 111796 20156
rect 111796 20100 111800 20156
rect 111736 20096 111800 20100
rect 111816 20156 111880 20160
rect 111816 20100 111820 20156
rect 111820 20100 111876 20156
rect 111876 20100 111880 20156
rect 111816 20096 111880 20100
rect 111896 20156 111960 20160
rect 111896 20100 111900 20156
rect 111900 20100 111956 20156
rect 111956 20100 111960 20156
rect 111896 20096 111960 20100
rect 111976 20156 112040 20160
rect 111976 20100 111980 20156
rect 111980 20100 112036 20156
rect 112036 20100 112040 20156
rect 111976 20096 112040 20100
rect 142456 20156 142520 20160
rect 142456 20100 142460 20156
rect 142460 20100 142516 20156
rect 142516 20100 142520 20156
rect 142456 20096 142520 20100
rect 142536 20156 142600 20160
rect 142536 20100 142540 20156
rect 142540 20100 142596 20156
rect 142596 20100 142600 20156
rect 142536 20096 142600 20100
rect 142616 20156 142680 20160
rect 142616 20100 142620 20156
rect 142620 20100 142676 20156
rect 142676 20100 142680 20156
rect 142616 20096 142680 20100
rect 142696 20156 142760 20160
rect 142696 20100 142700 20156
rect 142700 20100 142756 20156
rect 142756 20100 142760 20156
rect 142696 20096 142760 20100
rect 173176 20156 173240 20160
rect 173176 20100 173180 20156
rect 173180 20100 173236 20156
rect 173236 20100 173240 20156
rect 173176 20096 173240 20100
rect 173256 20156 173320 20160
rect 173256 20100 173260 20156
rect 173260 20100 173316 20156
rect 173316 20100 173320 20156
rect 173256 20096 173320 20100
rect 173336 20156 173400 20160
rect 173336 20100 173340 20156
rect 173340 20100 173396 20156
rect 173396 20100 173400 20156
rect 173336 20096 173400 20100
rect 173416 20156 173480 20160
rect 173416 20100 173420 20156
rect 173420 20100 173476 20156
rect 173476 20100 173480 20156
rect 173416 20096 173480 20100
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 34936 19612 35000 19616
rect 34936 19556 34940 19612
rect 34940 19556 34996 19612
rect 34996 19556 35000 19612
rect 34936 19552 35000 19556
rect 35016 19612 35080 19616
rect 35016 19556 35020 19612
rect 35020 19556 35076 19612
rect 35076 19556 35080 19612
rect 35016 19552 35080 19556
rect 35096 19612 35160 19616
rect 35096 19556 35100 19612
rect 35100 19556 35156 19612
rect 35156 19556 35160 19612
rect 35096 19552 35160 19556
rect 35176 19612 35240 19616
rect 35176 19556 35180 19612
rect 35180 19556 35236 19612
rect 35236 19556 35240 19612
rect 35176 19552 35240 19556
rect 65656 19612 65720 19616
rect 65656 19556 65660 19612
rect 65660 19556 65716 19612
rect 65716 19556 65720 19612
rect 65656 19552 65720 19556
rect 65736 19612 65800 19616
rect 65736 19556 65740 19612
rect 65740 19556 65796 19612
rect 65796 19556 65800 19612
rect 65736 19552 65800 19556
rect 65816 19612 65880 19616
rect 65816 19556 65820 19612
rect 65820 19556 65876 19612
rect 65876 19556 65880 19612
rect 65816 19552 65880 19556
rect 65896 19612 65960 19616
rect 65896 19556 65900 19612
rect 65900 19556 65956 19612
rect 65956 19556 65960 19612
rect 65896 19552 65960 19556
rect 96376 19612 96440 19616
rect 96376 19556 96380 19612
rect 96380 19556 96436 19612
rect 96436 19556 96440 19612
rect 96376 19552 96440 19556
rect 96456 19612 96520 19616
rect 96456 19556 96460 19612
rect 96460 19556 96516 19612
rect 96516 19556 96520 19612
rect 96456 19552 96520 19556
rect 96536 19612 96600 19616
rect 96536 19556 96540 19612
rect 96540 19556 96596 19612
rect 96596 19556 96600 19612
rect 96536 19552 96600 19556
rect 96616 19612 96680 19616
rect 96616 19556 96620 19612
rect 96620 19556 96676 19612
rect 96676 19556 96680 19612
rect 96616 19552 96680 19556
rect 127096 19612 127160 19616
rect 127096 19556 127100 19612
rect 127100 19556 127156 19612
rect 127156 19556 127160 19612
rect 127096 19552 127160 19556
rect 127176 19612 127240 19616
rect 127176 19556 127180 19612
rect 127180 19556 127236 19612
rect 127236 19556 127240 19612
rect 127176 19552 127240 19556
rect 127256 19612 127320 19616
rect 127256 19556 127260 19612
rect 127260 19556 127316 19612
rect 127316 19556 127320 19612
rect 127256 19552 127320 19556
rect 127336 19612 127400 19616
rect 127336 19556 127340 19612
rect 127340 19556 127396 19612
rect 127396 19556 127400 19612
rect 127336 19552 127400 19556
rect 157816 19612 157880 19616
rect 157816 19556 157820 19612
rect 157820 19556 157876 19612
rect 157876 19556 157880 19612
rect 157816 19552 157880 19556
rect 157896 19612 157960 19616
rect 157896 19556 157900 19612
rect 157900 19556 157956 19612
rect 157956 19556 157960 19612
rect 157896 19552 157960 19556
rect 157976 19612 158040 19616
rect 157976 19556 157980 19612
rect 157980 19556 158036 19612
rect 158036 19556 158040 19612
rect 157976 19552 158040 19556
rect 158056 19612 158120 19616
rect 158056 19556 158060 19612
rect 158060 19556 158116 19612
rect 158116 19556 158120 19612
rect 158056 19552 158120 19556
rect 19576 19068 19640 19072
rect 19576 19012 19580 19068
rect 19580 19012 19636 19068
rect 19636 19012 19640 19068
rect 19576 19008 19640 19012
rect 19656 19068 19720 19072
rect 19656 19012 19660 19068
rect 19660 19012 19716 19068
rect 19716 19012 19720 19068
rect 19656 19008 19720 19012
rect 19736 19068 19800 19072
rect 19736 19012 19740 19068
rect 19740 19012 19796 19068
rect 19796 19012 19800 19068
rect 19736 19008 19800 19012
rect 19816 19068 19880 19072
rect 19816 19012 19820 19068
rect 19820 19012 19876 19068
rect 19876 19012 19880 19068
rect 19816 19008 19880 19012
rect 50296 19068 50360 19072
rect 50296 19012 50300 19068
rect 50300 19012 50356 19068
rect 50356 19012 50360 19068
rect 50296 19008 50360 19012
rect 50376 19068 50440 19072
rect 50376 19012 50380 19068
rect 50380 19012 50436 19068
rect 50436 19012 50440 19068
rect 50376 19008 50440 19012
rect 50456 19068 50520 19072
rect 50456 19012 50460 19068
rect 50460 19012 50516 19068
rect 50516 19012 50520 19068
rect 50456 19008 50520 19012
rect 50536 19068 50600 19072
rect 50536 19012 50540 19068
rect 50540 19012 50596 19068
rect 50596 19012 50600 19068
rect 50536 19008 50600 19012
rect 81016 19068 81080 19072
rect 81016 19012 81020 19068
rect 81020 19012 81076 19068
rect 81076 19012 81080 19068
rect 81016 19008 81080 19012
rect 81096 19068 81160 19072
rect 81096 19012 81100 19068
rect 81100 19012 81156 19068
rect 81156 19012 81160 19068
rect 81096 19008 81160 19012
rect 81176 19068 81240 19072
rect 81176 19012 81180 19068
rect 81180 19012 81236 19068
rect 81236 19012 81240 19068
rect 81176 19008 81240 19012
rect 81256 19068 81320 19072
rect 81256 19012 81260 19068
rect 81260 19012 81316 19068
rect 81316 19012 81320 19068
rect 81256 19008 81320 19012
rect 111736 19068 111800 19072
rect 111736 19012 111740 19068
rect 111740 19012 111796 19068
rect 111796 19012 111800 19068
rect 111736 19008 111800 19012
rect 111816 19068 111880 19072
rect 111816 19012 111820 19068
rect 111820 19012 111876 19068
rect 111876 19012 111880 19068
rect 111816 19008 111880 19012
rect 111896 19068 111960 19072
rect 111896 19012 111900 19068
rect 111900 19012 111956 19068
rect 111956 19012 111960 19068
rect 111896 19008 111960 19012
rect 111976 19068 112040 19072
rect 111976 19012 111980 19068
rect 111980 19012 112036 19068
rect 112036 19012 112040 19068
rect 111976 19008 112040 19012
rect 142456 19068 142520 19072
rect 142456 19012 142460 19068
rect 142460 19012 142516 19068
rect 142516 19012 142520 19068
rect 142456 19008 142520 19012
rect 142536 19068 142600 19072
rect 142536 19012 142540 19068
rect 142540 19012 142596 19068
rect 142596 19012 142600 19068
rect 142536 19008 142600 19012
rect 142616 19068 142680 19072
rect 142616 19012 142620 19068
rect 142620 19012 142676 19068
rect 142676 19012 142680 19068
rect 142616 19008 142680 19012
rect 142696 19068 142760 19072
rect 142696 19012 142700 19068
rect 142700 19012 142756 19068
rect 142756 19012 142760 19068
rect 142696 19008 142760 19012
rect 173176 19068 173240 19072
rect 173176 19012 173180 19068
rect 173180 19012 173236 19068
rect 173236 19012 173240 19068
rect 173176 19008 173240 19012
rect 173256 19068 173320 19072
rect 173256 19012 173260 19068
rect 173260 19012 173316 19068
rect 173316 19012 173320 19068
rect 173256 19008 173320 19012
rect 173336 19068 173400 19072
rect 173336 19012 173340 19068
rect 173340 19012 173396 19068
rect 173396 19012 173400 19068
rect 173336 19008 173400 19012
rect 173416 19068 173480 19072
rect 173416 19012 173420 19068
rect 173420 19012 173476 19068
rect 173476 19012 173480 19068
rect 173416 19008 173480 19012
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 34936 18524 35000 18528
rect 34936 18468 34940 18524
rect 34940 18468 34996 18524
rect 34996 18468 35000 18524
rect 34936 18464 35000 18468
rect 35016 18524 35080 18528
rect 35016 18468 35020 18524
rect 35020 18468 35076 18524
rect 35076 18468 35080 18524
rect 35016 18464 35080 18468
rect 35096 18524 35160 18528
rect 35096 18468 35100 18524
rect 35100 18468 35156 18524
rect 35156 18468 35160 18524
rect 35096 18464 35160 18468
rect 35176 18524 35240 18528
rect 35176 18468 35180 18524
rect 35180 18468 35236 18524
rect 35236 18468 35240 18524
rect 35176 18464 35240 18468
rect 65656 18524 65720 18528
rect 65656 18468 65660 18524
rect 65660 18468 65716 18524
rect 65716 18468 65720 18524
rect 65656 18464 65720 18468
rect 65736 18524 65800 18528
rect 65736 18468 65740 18524
rect 65740 18468 65796 18524
rect 65796 18468 65800 18524
rect 65736 18464 65800 18468
rect 65816 18524 65880 18528
rect 65816 18468 65820 18524
rect 65820 18468 65876 18524
rect 65876 18468 65880 18524
rect 65816 18464 65880 18468
rect 65896 18524 65960 18528
rect 65896 18468 65900 18524
rect 65900 18468 65956 18524
rect 65956 18468 65960 18524
rect 65896 18464 65960 18468
rect 96376 18524 96440 18528
rect 96376 18468 96380 18524
rect 96380 18468 96436 18524
rect 96436 18468 96440 18524
rect 96376 18464 96440 18468
rect 96456 18524 96520 18528
rect 96456 18468 96460 18524
rect 96460 18468 96516 18524
rect 96516 18468 96520 18524
rect 96456 18464 96520 18468
rect 96536 18524 96600 18528
rect 96536 18468 96540 18524
rect 96540 18468 96596 18524
rect 96596 18468 96600 18524
rect 96536 18464 96600 18468
rect 96616 18524 96680 18528
rect 96616 18468 96620 18524
rect 96620 18468 96676 18524
rect 96676 18468 96680 18524
rect 96616 18464 96680 18468
rect 127096 18524 127160 18528
rect 127096 18468 127100 18524
rect 127100 18468 127156 18524
rect 127156 18468 127160 18524
rect 127096 18464 127160 18468
rect 127176 18524 127240 18528
rect 127176 18468 127180 18524
rect 127180 18468 127236 18524
rect 127236 18468 127240 18524
rect 127176 18464 127240 18468
rect 127256 18524 127320 18528
rect 127256 18468 127260 18524
rect 127260 18468 127316 18524
rect 127316 18468 127320 18524
rect 127256 18464 127320 18468
rect 127336 18524 127400 18528
rect 127336 18468 127340 18524
rect 127340 18468 127396 18524
rect 127396 18468 127400 18524
rect 127336 18464 127400 18468
rect 157816 18524 157880 18528
rect 157816 18468 157820 18524
rect 157820 18468 157876 18524
rect 157876 18468 157880 18524
rect 157816 18464 157880 18468
rect 157896 18524 157960 18528
rect 157896 18468 157900 18524
rect 157900 18468 157956 18524
rect 157956 18468 157960 18524
rect 157896 18464 157960 18468
rect 157976 18524 158040 18528
rect 157976 18468 157980 18524
rect 157980 18468 158036 18524
rect 158036 18468 158040 18524
rect 157976 18464 158040 18468
rect 158056 18524 158120 18528
rect 158056 18468 158060 18524
rect 158060 18468 158116 18524
rect 158116 18468 158120 18524
rect 158056 18464 158120 18468
rect 19576 17980 19640 17984
rect 19576 17924 19580 17980
rect 19580 17924 19636 17980
rect 19636 17924 19640 17980
rect 19576 17920 19640 17924
rect 19656 17980 19720 17984
rect 19656 17924 19660 17980
rect 19660 17924 19716 17980
rect 19716 17924 19720 17980
rect 19656 17920 19720 17924
rect 19736 17980 19800 17984
rect 19736 17924 19740 17980
rect 19740 17924 19796 17980
rect 19796 17924 19800 17980
rect 19736 17920 19800 17924
rect 19816 17980 19880 17984
rect 19816 17924 19820 17980
rect 19820 17924 19876 17980
rect 19876 17924 19880 17980
rect 19816 17920 19880 17924
rect 50296 17980 50360 17984
rect 50296 17924 50300 17980
rect 50300 17924 50356 17980
rect 50356 17924 50360 17980
rect 50296 17920 50360 17924
rect 50376 17980 50440 17984
rect 50376 17924 50380 17980
rect 50380 17924 50436 17980
rect 50436 17924 50440 17980
rect 50376 17920 50440 17924
rect 50456 17980 50520 17984
rect 50456 17924 50460 17980
rect 50460 17924 50516 17980
rect 50516 17924 50520 17980
rect 50456 17920 50520 17924
rect 50536 17980 50600 17984
rect 50536 17924 50540 17980
rect 50540 17924 50596 17980
rect 50596 17924 50600 17980
rect 50536 17920 50600 17924
rect 81016 17980 81080 17984
rect 81016 17924 81020 17980
rect 81020 17924 81076 17980
rect 81076 17924 81080 17980
rect 81016 17920 81080 17924
rect 81096 17980 81160 17984
rect 81096 17924 81100 17980
rect 81100 17924 81156 17980
rect 81156 17924 81160 17980
rect 81096 17920 81160 17924
rect 81176 17980 81240 17984
rect 81176 17924 81180 17980
rect 81180 17924 81236 17980
rect 81236 17924 81240 17980
rect 81176 17920 81240 17924
rect 81256 17980 81320 17984
rect 81256 17924 81260 17980
rect 81260 17924 81316 17980
rect 81316 17924 81320 17980
rect 81256 17920 81320 17924
rect 111736 17980 111800 17984
rect 111736 17924 111740 17980
rect 111740 17924 111796 17980
rect 111796 17924 111800 17980
rect 111736 17920 111800 17924
rect 111816 17980 111880 17984
rect 111816 17924 111820 17980
rect 111820 17924 111876 17980
rect 111876 17924 111880 17980
rect 111816 17920 111880 17924
rect 111896 17980 111960 17984
rect 111896 17924 111900 17980
rect 111900 17924 111956 17980
rect 111956 17924 111960 17980
rect 111896 17920 111960 17924
rect 111976 17980 112040 17984
rect 111976 17924 111980 17980
rect 111980 17924 112036 17980
rect 112036 17924 112040 17980
rect 111976 17920 112040 17924
rect 142456 17980 142520 17984
rect 142456 17924 142460 17980
rect 142460 17924 142516 17980
rect 142516 17924 142520 17980
rect 142456 17920 142520 17924
rect 142536 17980 142600 17984
rect 142536 17924 142540 17980
rect 142540 17924 142596 17980
rect 142596 17924 142600 17980
rect 142536 17920 142600 17924
rect 142616 17980 142680 17984
rect 142616 17924 142620 17980
rect 142620 17924 142676 17980
rect 142676 17924 142680 17980
rect 142616 17920 142680 17924
rect 142696 17980 142760 17984
rect 142696 17924 142700 17980
rect 142700 17924 142756 17980
rect 142756 17924 142760 17980
rect 142696 17920 142760 17924
rect 173176 17980 173240 17984
rect 173176 17924 173180 17980
rect 173180 17924 173236 17980
rect 173236 17924 173240 17980
rect 173176 17920 173240 17924
rect 173256 17980 173320 17984
rect 173256 17924 173260 17980
rect 173260 17924 173316 17980
rect 173316 17924 173320 17980
rect 173256 17920 173320 17924
rect 173336 17980 173400 17984
rect 173336 17924 173340 17980
rect 173340 17924 173396 17980
rect 173396 17924 173400 17980
rect 173336 17920 173400 17924
rect 173416 17980 173480 17984
rect 173416 17924 173420 17980
rect 173420 17924 173476 17980
rect 173476 17924 173480 17980
rect 173416 17920 173480 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 34936 17436 35000 17440
rect 34936 17380 34940 17436
rect 34940 17380 34996 17436
rect 34996 17380 35000 17436
rect 34936 17376 35000 17380
rect 35016 17436 35080 17440
rect 35016 17380 35020 17436
rect 35020 17380 35076 17436
rect 35076 17380 35080 17436
rect 35016 17376 35080 17380
rect 35096 17436 35160 17440
rect 35096 17380 35100 17436
rect 35100 17380 35156 17436
rect 35156 17380 35160 17436
rect 35096 17376 35160 17380
rect 35176 17436 35240 17440
rect 35176 17380 35180 17436
rect 35180 17380 35236 17436
rect 35236 17380 35240 17436
rect 35176 17376 35240 17380
rect 65656 17436 65720 17440
rect 65656 17380 65660 17436
rect 65660 17380 65716 17436
rect 65716 17380 65720 17436
rect 65656 17376 65720 17380
rect 65736 17436 65800 17440
rect 65736 17380 65740 17436
rect 65740 17380 65796 17436
rect 65796 17380 65800 17436
rect 65736 17376 65800 17380
rect 65816 17436 65880 17440
rect 65816 17380 65820 17436
rect 65820 17380 65876 17436
rect 65876 17380 65880 17436
rect 65816 17376 65880 17380
rect 65896 17436 65960 17440
rect 65896 17380 65900 17436
rect 65900 17380 65956 17436
rect 65956 17380 65960 17436
rect 65896 17376 65960 17380
rect 96376 17436 96440 17440
rect 96376 17380 96380 17436
rect 96380 17380 96436 17436
rect 96436 17380 96440 17436
rect 96376 17376 96440 17380
rect 96456 17436 96520 17440
rect 96456 17380 96460 17436
rect 96460 17380 96516 17436
rect 96516 17380 96520 17436
rect 96456 17376 96520 17380
rect 96536 17436 96600 17440
rect 96536 17380 96540 17436
rect 96540 17380 96596 17436
rect 96596 17380 96600 17436
rect 96536 17376 96600 17380
rect 96616 17436 96680 17440
rect 96616 17380 96620 17436
rect 96620 17380 96676 17436
rect 96676 17380 96680 17436
rect 96616 17376 96680 17380
rect 127096 17436 127160 17440
rect 127096 17380 127100 17436
rect 127100 17380 127156 17436
rect 127156 17380 127160 17436
rect 127096 17376 127160 17380
rect 127176 17436 127240 17440
rect 127176 17380 127180 17436
rect 127180 17380 127236 17436
rect 127236 17380 127240 17436
rect 127176 17376 127240 17380
rect 127256 17436 127320 17440
rect 127256 17380 127260 17436
rect 127260 17380 127316 17436
rect 127316 17380 127320 17436
rect 127256 17376 127320 17380
rect 127336 17436 127400 17440
rect 127336 17380 127340 17436
rect 127340 17380 127396 17436
rect 127396 17380 127400 17436
rect 127336 17376 127400 17380
rect 157816 17436 157880 17440
rect 157816 17380 157820 17436
rect 157820 17380 157876 17436
rect 157876 17380 157880 17436
rect 157816 17376 157880 17380
rect 157896 17436 157960 17440
rect 157896 17380 157900 17436
rect 157900 17380 157956 17436
rect 157956 17380 157960 17436
rect 157896 17376 157960 17380
rect 157976 17436 158040 17440
rect 157976 17380 157980 17436
rect 157980 17380 158036 17436
rect 158036 17380 158040 17436
rect 157976 17376 158040 17380
rect 158056 17436 158120 17440
rect 158056 17380 158060 17436
rect 158060 17380 158116 17436
rect 158116 17380 158120 17436
rect 158056 17376 158120 17380
rect 19576 16892 19640 16896
rect 19576 16836 19580 16892
rect 19580 16836 19636 16892
rect 19636 16836 19640 16892
rect 19576 16832 19640 16836
rect 19656 16892 19720 16896
rect 19656 16836 19660 16892
rect 19660 16836 19716 16892
rect 19716 16836 19720 16892
rect 19656 16832 19720 16836
rect 19736 16892 19800 16896
rect 19736 16836 19740 16892
rect 19740 16836 19796 16892
rect 19796 16836 19800 16892
rect 19736 16832 19800 16836
rect 19816 16892 19880 16896
rect 19816 16836 19820 16892
rect 19820 16836 19876 16892
rect 19876 16836 19880 16892
rect 19816 16832 19880 16836
rect 50296 16892 50360 16896
rect 50296 16836 50300 16892
rect 50300 16836 50356 16892
rect 50356 16836 50360 16892
rect 50296 16832 50360 16836
rect 50376 16892 50440 16896
rect 50376 16836 50380 16892
rect 50380 16836 50436 16892
rect 50436 16836 50440 16892
rect 50376 16832 50440 16836
rect 50456 16892 50520 16896
rect 50456 16836 50460 16892
rect 50460 16836 50516 16892
rect 50516 16836 50520 16892
rect 50456 16832 50520 16836
rect 50536 16892 50600 16896
rect 50536 16836 50540 16892
rect 50540 16836 50596 16892
rect 50596 16836 50600 16892
rect 50536 16832 50600 16836
rect 81016 16892 81080 16896
rect 81016 16836 81020 16892
rect 81020 16836 81076 16892
rect 81076 16836 81080 16892
rect 81016 16832 81080 16836
rect 81096 16892 81160 16896
rect 81096 16836 81100 16892
rect 81100 16836 81156 16892
rect 81156 16836 81160 16892
rect 81096 16832 81160 16836
rect 81176 16892 81240 16896
rect 81176 16836 81180 16892
rect 81180 16836 81236 16892
rect 81236 16836 81240 16892
rect 81176 16832 81240 16836
rect 81256 16892 81320 16896
rect 81256 16836 81260 16892
rect 81260 16836 81316 16892
rect 81316 16836 81320 16892
rect 81256 16832 81320 16836
rect 111736 16892 111800 16896
rect 111736 16836 111740 16892
rect 111740 16836 111796 16892
rect 111796 16836 111800 16892
rect 111736 16832 111800 16836
rect 111816 16892 111880 16896
rect 111816 16836 111820 16892
rect 111820 16836 111876 16892
rect 111876 16836 111880 16892
rect 111816 16832 111880 16836
rect 111896 16892 111960 16896
rect 111896 16836 111900 16892
rect 111900 16836 111956 16892
rect 111956 16836 111960 16892
rect 111896 16832 111960 16836
rect 111976 16892 112040 16896
rect 111976 16836 111980 16892
rect 111980 16836 112036 16892
rect 112036 16836 112040 16892
rect 111976 16832 112040 16836
rect 142456 16892 142520 16896
rect 142456 16836 142460 16892
rect 142460 16836 142516 16892
rect 142516 16836 142520 16892
rect 142456 16832 142520 16836
rect 142536 16892 142600 16896
rect 142536 16836 142540 16892
rect 142540 16836 142596 16892
rect 142596 16836 142600 16892
rect 142536 16832 142600 16836
rect 142616 16892 142680 16896
rect 142616 16836 142620 16892
rect 142620 16836 142676 16892
rect 142676 16836 142680 16892
rect 142616 16832 142680 16836
rect 142696 16892 142760 16896
rect 142696 16836 142700 16892
rect 142700 16836 142756 16892
rect 142756 16836 142760 16892
rect 142696 16832 142760 16836
rect 173176 16892 173240 16896
rect 173176 16836 173180 16892
rect 173180 16836 173236 16892
rect 173236 16836 173240 16892
rect 173176 16832 173240 16836
rect 173256 16892 173320 16896
rect 173256 16836 173260 16892
rect 173260 16836 173316 16892
rect 173316 16836 173320 16892
rect 173256 16832 173320 16836
rect 173336 16892 173400 16896
rect 173336 16836 173340 16892
rect 173340 16836 173396 16892
rect 173396 16836 173400 16892
rect 173336 16832 173400 16836
rect 173416 16892 173480 16896
rect 173416 16836 173420 16892
rect 173420 16836 173476 16892
rect 173476 16836 173480 16892
rect 173416 16832 173480 16836
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 34936 16348 35000 16352
rect 34936 16292 34940 16348
rect 34940 16292 34996 16348
rect 34996 16292 35000 16348
rect 34936 16288 35000 16292
rect 35016 16348 35080 16352
rect 35016 16292 35020 16348
rect 35020 16292 35076 16348
rect 35076 16292 35080 16348
rect 35016 16288 35080 16292
rect 35096 16348 35160 16352
rect 35096 16292 35100 16348
rect 35100 16292 35156 16348
rect 35156 16292 35160 16348
rect 35096 16288 35160 16292
rect 35176 16348 35240 16352
rect 35176 16292 35180 16348
rect 35180 16292 35236 16348
rect 35236 16292 35240 16348
rect 35176 16288 35240 16292
rect 65656 16348 65720 16352
rect 65656 16292 65660 16348
rect 65660 16292 65716 16348
rect 65716 16292 65720 16348
rect 65656 16288 65720 16292
rect 65736 16348 65800 16352
rect 65736 16292 65740 16348
rect 65740 16292 65796 16348
rect 65796 16292 65800 16348
rect 65736 16288 65800 16292
rect 65816 16348 65880 16352
rect 65816 16292 65820 16348
rect 65820 16292 65876 16348
rect 65876 16292 65880 16348
rect 65816 16288 65880 16292
rect 65896 16348 65960 16352
rect 65896 16292 65900 16348
rect 65900 16292 65956 16348
rect 65956 16292 65960 16348
rect 65896 16288 65960 16292
rect 96376 16348 96440 16352
rect 96376 16292 96380 16348
rect 96380 16292 96436 16348
rect 96436 16292 96440 16348
rect 96376 16288 96440 16292
rect 96456 16348 96520 16352
rect 96456 16292 96460 16348
rect 96460 16292 96516 16348
rect 96516 16292 96520 16348
rect 96456 16288 96520 16292
rect 96536 16348 96600 16352
rect 96536 16292 96540 16348
rect 96540 16292 96596 16348
rect 96596 16292 96600 16348
rect 96536 16288 96600 16292
rect 96616 16348 96680 16352
rect 96616 16292 96620 16348
rect 96620 16292 96676 16348
rect 96676 16292 96680 16348
rect 96616 16288 96680 16292
rect 127096 16348 127160 16352
rect 127096 16292 127100 16348
rect 127100 16292 127156 16348
rect 127156 16292 127160 16348
rect 127096 16288 127160 16292
rect 127176 16348 127240 16352
rect 127176 16292 127180 16348
rect 127180 16292 127236 16348
rect 127236 16292 127240 16348
rect 127176 16288 127240 16292
rect 127256 16348 127320 16352
rect 127256 16292 127260 16348
rect 127260 16292 127316 16348
rect 127316 16292 127320 16348
rect 127256 16288 127320 16292
rect 127336 16348 127400 16352
rect 127336 16292 127340 16348
rect 127340 16292 127396 16348
rect 127396 16292 127400 16348
rect 127336 16288 127400 16292
rect 157816 16348 157880 16352
rect 157816 16292 157820 16348
rect 157820 16292 157876 16348
rect 157876 16292 157880 16348
rect 157816 16288 157880 16292
rect 157896 16348 157960 16352
rect 157896 16292 157900 16348
rect 157900 16292 157956 16348
rect 157956 16292 157960 16348
rect 157896 16288 157960 16292
rect 157976 16348 158040 16352
rect 157976 16292 157980 16348
rect 157980 16292 158036 16348
rect 158036 16292 158040 16348
rect 157976 16288 158040 16292
rect 158056 16348 158120 16352
rect 158056 16292 158060 16348
rect 158060 16292 158116 16348
rect 158116 16292 158120 16348
rect 158056 16288 158120 16292
rect 19576 15804 19640 15808
rect 19576 15748 19580 15804
rect 19580 15748 19636 15804
rect 19636 15748 19640 15804
rect 19576 15744 19640 15748
rect 19656 15804 19720 15808
rect 19656 15748 19660 15804
rect 19660 15748 19716 15804
rect 19716 15748 19720 15804
rect 19656 15744 19720 15748
rect 19736 15804 19800 15808
rect 19736 15748 19740 15804
rect 19740 15748 19796 15804
rect 19796 15748 19800 15804
rect 19736 15744 19800 15748
rect 19816 15804 19880 15808
rect 19816 15748 19820 15804
rect 19820 15748 19876 15804
rect 19876 15748 19880 15804
rect 19816 15744 19880 15748
rect 50296 15804 50360 15808
rect 50296 15748 50300 15804
rect 50300 15748 50356 15804
rect 50356 15748 50360 15804
rect 50296 15744 50360 15748
rect 50376 15804 50440 15808
rect 50376 15748 50380 15804
rect 50380 15748 50436 15804
rect 50436 15748 50440 15804
rect 50376 15744 50440 15748
rect 50456 15804 50520 15808
rect 50456 15748 50460 15804
rect 50460 15748 50516 15804
rect 50516 15748 50520 15804
rect 50456 15744 50520 15748
rect 50536 15804 50600 15808
rect 50536 15748 50540 15804
rect 50540 15748 50596 15804
rect 50596 15748 50600 15804
rect 50536 15744 50600 15748
rect 81016 15804 81080 15808
rect 81016 15748 81020 15804
rect 81020 15748 81076 15804
rect 81076 15748 81080 15804
rect 81016 15744 81080 15748
rect 81096 15804 81160 15808
rect 81096 15748 81100 15804
rect 81100 15748 81156 15804
rect 81156 15748 81160 15804
rect 81096 15744 81160 15748
rect 81176 15804 81240 15808
rect 81176 15748 81180 15804
rect 81180 15748 81236 15804
rect 81236 15748 81240 15804
rect 81176 15744 81240 15748
rect 81256 15804 81320 15808
rect 81256 15748 81260 15804
rect 81260 15748 81316 15804
rect 81316 15748 81320 15804
rect 81256 15744 81320 15748
rect 111736 15804 111800 15808
rect 111736 15748 111740 15804
rect 111740 15748 111796 15804
rect 111796 15748 111800 15804
rect 111736 15744 111800 15748
rect 111816 15804 111880 15808
rect 111816 15748 111820 15804
rect 111820 15748 111876 15804
rect 111876 15748 111880 15804
rect 111816 15744 111880 15748
rect 111896 15804 111960 15808
rect 111896 15748 111900 15804
rect 111900 15748 111956 15804
rect 111956 15748 111960 15804
rect 111896 15744 111960 15748
rect 111976 15804 112040 15808
rect 111976 15748 111980 15804
rect 111980 15748 112036 15804
rect 112036 15748 112040 15804
rect 111976 15744 112040 15748
rect 142456 15804 142520 15808
rect 142456 15748 142460 15804
rect 142460 15748 142516 15804
rect 142516 15748 142520 15804
rect 142456 15744 142520 15748
rect 142536 15804 142600 15808
rect 142536 15748 142540 15804
rect 142540 15748 142596 15804
rect 142596 15748 142600 15804
rect 142536 15744 142600 15748
rect 142616 15804 142680 15808
rect 142616 15748 142620 15804
rect 142620 15748 142676 15804
rect 142676 15748 142680 15804
rect 142616 15744 142680 15748
rect 142696 15804 142760 15808
rect 142696 15748 142700 15804
rect 142700 15748 142756 15804
rect 142756 15748 142760 15804
rect 142696 15744 142760 15748
rect 173176 15804 173240 15808
rect 173176 15748 173180 15804
rect 173180 15748 173236 15804
rect 173236 15748 173240 15804
rect 173176 15744 173240 15748
rect 173256 15804 173320 15808
rect 173256 15748 173260 15804
rect 173260 15748 173316 15804
rect 173316 15748 173320 15804
rect 173256 15744 173320 15748
rect 173336 15804 173400 15808
rect 173336 15748 173340 15804
rect 173340 15748 173396 15804
rect 173396 15748 173400 15804
rect 173336 15744 173400 15748
rect 173416 15804 173480 15808
rect 173416 15748 173420 15804
rect 173420 15748 173476 15804
rect 173476 15748 173480 15804
rect 173416 15744 173480 15748
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 34936 15260 35000 15264
rect 34936 15204 34940 15260
rect 34940 15204 34996 15260
rect 34996 15204 35000 15260
rect 34936 15200 35000 15204
rect 35016 15260 35080 15264
rect 35016 15204 35020 15260
rect 35020 15204 35076 15260
rect 35076 15204 35080 15260
rect 35016 15200 35080 15204
rect 35096 15260 35160 15264
rect 35096 15204 35100 15260
rect 35100 15204 35156 15260
rect 35156 15204 35160 15260
rect 35096 15200 35160 15204
rect 35176 15260 35240 15264
rect 35176 15204 35180 15260
rect 35180 15204 35236 15260
rect 35236 15204 35240 15260
rect 35176 15200 35240 15204
rect 65656 15260 65720 15264
rect 65656 15204 65660 15260
rect 65660 15204 65716 15260
rect 65716 15204 65720 15260
rect 65656 15200 65720 15204
rect 65736 15260 65800 15264
rect 65736 15204 65740 15260
rect 65740 15204 65796 15260
rect 65796 15204 65800 15260
rect 65736 15200 65800 15204
rect 65816 15260 65880 15264
rect 65816 15204 65820 15260
rect 65820 15204 65876 15260
rect 65876 15204 65880 15260
rect 65816 15200 65880 15204
rect 65896 15260 65960 15264
rect 65896 15204 65900 15260
rect 65900 15204 65956 15260
rect 65956 15204 65960 15260
rect 65896 15200 65960 15204
rect 96376 15260 96440 15264
rect 96376 15204 96380 15260
rect 96380 15204 96436 15260
rect 96436 15204 96440 15260
rect 96376 15200 96440 15204
rect 96456 15260 96520 15264
rect 96456 15204 96460 15260
rect 96460 15204 96516 15260
rect 96516 15204 96520 15260
rect 96456 15200 96520 15204
rect 96536 15260 96600 15264
rect 96536 15204 96540 15260
rect 96540 15204 96596 15260
rect 96596 15204 96600 15260
rect 96536 15200 96600 15204
rect 96616 15260 96680 15264
rect 96616 15204 96620 15260
rect 96620 15204 96676 15260
rect 96676 15204 96680 15260
rect 96616 15200 96680 15204
rect 127096 15260 127160 15264
rect 127096 15204 127100 15260
rect 127100 15204 127156 15260
rect 127156 15204 127160 15260
rect 127096 15200 127160 15204
rect 127176 15260 127240 15264
rect 127176 15204 127180 15260
rect 127180 15204 127236 15260
rect 127236 15204 127240 15260
rect 127176 15200 127240 15204
rect 127256 15260 127320 15264
rect 127256 15204 127260 15260
rect 127260 15204 127316 15260
rect 127316 15204 127320 15260
rect 127256 15200 127320 15204
rect 127336 15260 127400 15264
rect 127336 15204 127340 15260
rect 127340 15204 127396 15260
rect 127396 15204 127400 15260
rect 127336 15200 127400 15204
rect 157816 15260 157880 15264
rect 157816 15204 157820 15260
rect 157820 15204 157876 15260
rect 157876 15204 157880 15260
rect 157816 15200 157880 15204
rect 157896 15260 157960 15264
rect 157896 15204 157900 15260
rect 157900 15204 157956 15260
rect 157956 15204 157960 15260
rect 157896 15200 157960 15204
rect 157976 15260 158040 15264
rect 157976 15204 157980 15260
rect 157980 15204 158036 15260
rect 158036 15204 158040 15260
rect 157976 15200 158040 15204
rect 158056 15260 158120 15264
rect 158056 15204 158060 15260
rect 158060 15204 158116 15260
rect 158116 15204 158120 15260
rect 158056 15200 158120 15204
rect 19576 14716 19640 14720
rect 19576 14660 19580 14716
rect 19580 14660 19636 14716
rect 19636 14660 19640 14716
rect 19576 14656 19640 14660
rect 19656 14716 19720 14720
rect 19656 14660 19660 14716
rect 19660 14660 19716 14716
rect 19716 14660 19720 14716
rect 19656 14656 19720 14660
rect 19736 14716 19800 14720
rect 19736 14660 19740 14716
rect 19740 14660 19796 14716
rect 19796 14660 19800 14716
rect 19736 14656 19800 14660
rect 19816 14716 19880 14720
rect 19816 14660 19820 14716
rect 19820 14660 19876 14716
rect 19876 14660 19880 14716
rect 19816 14656 19880 14660
rect 50296 14716 50360 14720
rect 50296 14660 50300 14716
rect 50300 14660 50356 14716
rect 50356 14660 50360 14716
rect 50296 14656 50360 14660
rect 50376 14716 50440 14720
rect 50376 14660 50380 14716
rect 50380 14660 50436 14716
rect 50436 14660 50440 14716
rect 50376 14656 50440 14660
rect 50456 14716 50520 14720
rect 50456 14660 50460 14716
rect 50460 14660 50516 14716
rect 50516 14660 50520 14716
rect 50456 14656 50520 14660
rect 50536 14716 50600 14720
rect 50536 14660 50540 14716
rect 50540 14660 50596 14716
rect 50596 14660 50600 14716
rect 50536 14656 50600 14660
rect 81016 14716 81080 14720
rect 81016 14660 81020 14716
rect 81020 14660 81076 14716
rect 81076 14660 81080 14716
rect 81016 14656 81080 14660
rect 81096 14716 81160 14720
rect 81096 14660 81100 14716
rect 81100 14660 81156 14716
rect 81156 14660 81160 14716
rect 81096 14656 81160 14660
rect 81176 14716 81240 14720
rect 81176 14660 81180 14716
rect 81180 14660 81236 14716
rect 81236 14660 81240 14716
rect 81176 14656 81240 14660
rect 81256 14716 81320 14720
rect 81256 14660 81260 14716
rect 81260 14660 81316 14716
rect 81316 14660 81320 14716
rect 81256 14656 81320 14660
rect 111736 14716 111800 14720
rect 111736 14660 111740 14716
rect 111740 14660 111796 14716
rect 111796 14660 111800 14716
rect 111736 14656 111800 14660
rect 111816 14716 111880 14720
rect 111816 14660 111820 14716
rect 111820 14660 111876 14716
rect 111876 14660 111880 14716
rect 111816 14656 111880 14660
rect 111896 14716 111960 14720
rect 111896 14660 111900 14716
rect 111900 14660 111956 14716
rect 111956 14660 111960 14716
rect 111896 14656 111960 14660
rect 111976 14716 112040 14720
rect 111976 14660 111980 14716
rect 111980 14660 112036 14716
rect 112036 14660 112040 14716
rect 111976 14656 112040 14660
rect 142456 14716 142520 14720
rect 142456 14660 142460 14716
rect 142460 14660 142516 14716
rect 142516 14660 142520 14716
rect 142456 14656 142520 14660
rect 142536 14716 142600 14720
rect 142536 14660 142540 14716
rect 142540 14660 142596 14716
rect 142596 14660 142600 14716
rect 142536 14656 142600 14660
rect 142616 14716 142680 14720
rect 142616 14660 142620 14716
rect 142620 14660 142676 14716
rect 142676 14660 142680 14716
rect 142616 14656 142680 14660
rect 142696 14716 142760 14720
rect 142696 14660 142700 14716
rect 142700 14660 142756 14716
rect 142756 14660 142760 14716
rect 142696 14656 142760 14660
rect 173176 14716 173240 14720
rect 173176 14660 173180 14716
rect 173180 14660 173236 14716
rect 173236 14660 173240 14716
rect 173176 14656 173240 14660
rect 173256 14716 173320 14720
rect 173256 14660 173260 14716
rect 173260 14660 173316 14716
rect 173316 14660 173320 14716
rect 173256 14656 173320 14660
rect 173336 14716 173400 14720
rect 173336 14660 173340 14716
rect 173340 14660 173396 14716
rect 173396 14660 173400 14716
rect 173336 14656 173400 14660
rect 173416 14716 173480 14720
rect 173416 14660 173420 14716
rect 173420 14660 173476 14716
rect 173476 14660 173480 14716
rect 173416 14656 173480 14660
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 34936 14172 35000 14176
rect 34936 14116 34940 14172
rect 34940 14116 34996 14172
rect 34996 14116 35000 14172
rect 34936 14112 35000 14116
rect 35016 14172 35080 14176
rect 35016 14116 35020 14172
rect 35020 14116 35076 14172
rect 35076 14116 35080 14172
rect 35016 14112 35080 14116
rect 35096 14172 35160 14176
rect 35096 14116 35100 14172
rect 35100 14116 35156 14172
rect 35156 14116 35160 14172
rect 35096 14112 35160 14116
rect 35176 14172 35240 14176
rect 35176 14116 35180 14172
rect 35180 14116 35236 14172
rect 35236 14116 35240 14172
rect 35176 14112 35240 14116
rect 65656 14172 65720 14176
rect 65656 14116 65660 14172
rect 65660 14116 65716 14172
rect 65716 14116 65720 14172
rect 65656 14112 65720 14116
rect 65736 14172 65800 14176
rect 65736 14116 65740 14172
rect 65740 14116 65796 14172
rect 65796 14116 65800 14172
rect 65736 14112 65800 14116
rect 65816 14172 65880 14176
rect 65816 14116 65820 14172
rect 65820 14116 65876 14172
rect 65876 14116 65880 14172
rect 65816 14112 65880 14116
rect 65896 14172 65960 14176
rect 65896 14116 65900 14172
rect 65900 14116 65956 14172
rect 65956 14116 65960 14172
rect 65896 14112 65960 14116
rect 96376 14172 96440 14176
rect 96376 14116 96380 14172
rect 96380 14116 96436 14172
rect 96436 14116 96440 14172
rect 96376 14112 96440 14116
rect 96456 14172 96520 14176
rect 96456 14116 96460 14172
rect 96460 14116 96516 14172
rect 96516 14116 96520 14172
rect 96456 14112 96520 14116
rect 96536 14172 96600 14176
rect 96536 14116 96540 14172
rect 96540 14116 96596 14172
rect 96596 14116 96600 14172
rect 96536 14112 96600 14116
rect 96616 14172 96680 14176
rect 96616 14116 96620 14172
rect 96620 14116 96676 14172
rect 96676 14116 96680 14172
rect 96616 14112 96680 14116
rect 127096 14172 127160 14176
rect 127096 14116 127100 14172
rect 127100 14116 127156 14172
rect 127156 14116 127160 14172
rect 127096 14112 127160 14116
rect 127176 14172 127240 14176
rect 127176 14116 127180 14172
rect 127180 14116 127236 14172
rect 127236 14116 127240 14172
rect 127176 14112 127240 14116
rect 127256 14172 127320 14176
rect 127256 14116 127260 14172
rect 127260 14116 127316 14172
rect 127316 14116 127320 14172
rect 127256 14112 127320 14116
rect 127336 14172 127400 14176
rect 127336 14116 127340 14172
rect 127340 14116 127396 14172
rect 127396 14116 127400 14172
rect 127336 14112 127400 14116
rect 157816 14172 157880 14176
rect 157816 14116 157820 14172
rect 157820 14116 157876 14172
rect 157876 14116 157880 14172
rect 157816 14112 157880 14116
rect 157896 14172 157960 14176
rect 157896 14116 157900 14172
rect 157900 14116 157956 14172
rect 157956 14116 157960 14172
rect 157896 14112 157960 14116
rect 157976 14172 158040 14176
rect 157976 14116 157980 14172
rect 157980 14116 158036 14172
rect 158036 14116 158040 14172
rect 157976 14112 158040 14116
rect 158056 14172 158120 14176
rect 158056 14116 158060 14172
rect 158060 14116 158116 14172
rect 158116 14116 158120 14172
rect 158056 14112 158120 14116
rect 19576 13628 19640 13632
rect 19576 13572 19580 13628
rect 19580 13572 19636 13628
rect 19636 13572 19640 13628
rect 19576 13568 19640 13572
rect 19656 13628 19720 13632
rect 19656 13572 19660 13628
rect 19660 13572 19716 13628
rect 19716 13572 19720 13628
rect 19656 13568 19720 13572
rect 19736 13628 19800 13632
rect 19736 13572 19740 13628
rect 19740 13572 19796 13628
rect 19796 13572 19800 13628
rect 19736 13568 19800 13572
rect 19816 13628 19880 13632
rect 19816 13572 19820 13628
rect 19820 13572 19876 13628
rect 19876 13572 19880 13628
rect 19816 13568 19880 13572
rect 50296 13628 50360 13632
rect 50296 13572 50300 13628
rect 50300 13572 50356 13628
rect 50356 13572 50360 13628
rect 50296 13568 50360 13572
rect 50376 13628 50440 13632
rect 50376 13572 50380 13628
rect 50380 13572 50436 13628
rect 50436 13572 50440 13628
rect 50376 13568 50440 13572
rect 50456 13628 50520 13632
rect 50456 13572 50460 13628
rect 50460 13572 50516 13628
rect 50516 13572 50520 13628
rect 50456 13568 50520 13572
rect 50536 13628 50600 13632
rect 50536 13572 50540 13628
rect 50540 13572 50596 13628
rect 50596 13572 50600 13628
rect 50536 13568 50600 13572
rect 81016 13628 81080 13632
rect 81016 13572 81020 13628
rect 81020 13572 81076 13628
rect 81076 13572 81080 13628
rect 81016 13568 81080 13572
rect 81096 13628 81160 13632
rect 81096 13572 81100 13628
rect 81100 13572 81156 13628
rect 81156 13572 81160 13628
rect 81096 13568 81160 13572
rect 81176 13628 81240 13632
rect 81176 13572 81180 13628
rect 81180 13572 81236 13628
rect 81236 13572 81240 13628
rect 81176 13568 81240 13572
rect 81256 13628 81320 13632
rect 81256 13572 81260 13628
rect 81260 13572 81316 13628
rect 81316 13572 81320 13628
rect 81256 13568 81320 13572
rect 111736 13628 111800 13632
rect 111736 13572 111740 13628
rect 111740 13572 111796 13628
rect 111796 13572 111800 13628
rect 111736 13568 111800 13572
rect 111816 13628 111880 13632
rect 111816 13572 111820 13628
rect 111820 13572 111876 13628
rect 111876 13572 111880 13628
rect 111816 13568 111880 13572
rect 111896 13628 111960 13632
rect 111896 13572 111900 13628
rect 111900 13572 111956 13628
rect 111956 13572 111960 13628
rect 111896 13568 111960 13572
rect 111976 13628 112040 13632
rect 111976 13572 111980 13628
rect 111980 13572 112036 13628
rect 112036 13572 112040 13628
rect 111976 13568 112040 13572
rect 142456 13628 142520 13632
rect 142456 13572 142460 13628
rect 142460 13572 142516 13628
rect 142516 13572 142520 13628
rect 142456 13568 142520 13572
rect 142536 13628 142600 13632
rect 142536 13572 142540 13628
rect 142540 13572 142596 13628
rect 142596 13572 142600 13628
rect 142536 13568 142600 13572
rect 142616 13628 142680 13632
rect 142616 13572 142620 13628
rect 142620 13572 142676 13628
rect 142676 13572 142680 13628
rect 142616 13568 142680 13572
rect 142696 13628 142760 13632
rect 142696 13572 142700 13628
rect 142700 13572 142756 13628
rect 142756 13572 142760 13628
rect 142696 13568 142760 13572
rect 173176 13628 173240 13632
rect 173176 13572 173180 13628
rect 173180 13572 173236 13628
rect 173236 13572 173240 13628
rect 173176 13568 173240 13572
rect 173256 13628 173320 13632
rect 173256 13572 173260 13628
rect 173260 13572 173316 13628
rect 173316 13572 173320 13628
rect 173256 13568 173320 13572
rect 173336 13628 173400 13632
rect 173336 13572 173340 13628
rect 173340 13572 173396 13628
rect 173396 13572 173400 13628
rect 173336 13568 173400 13572
rect 173416 13628 173480 13632
rect 173416 13572 173420 13628
rect 173420 13572 173476 13628
rect 173476 13572 173480 13628
rect 173416 13568 173480 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 34936 13084 35000 13088
rect 34936 13028 34940 13084
rect 34940 13028 34996 13084
rect 34996 13028 35000 13084
rect 34936 13024 35000 13028
rect 35016 13084 35080 13088
rect 35016 13028 35020 13084
rect 35020 13028 35076 13084
rect 35076 13028 35080 13084
rect 35016 13024 35080 13028
rect 35096 13084 35160 13088
rect 35096 13028 35100 13084
rect 35100 13028 35156 13084
rect 35156 13028 35160 13084
rect 35096 13024 35160 13028
rect 35176 13084 35240 13088
rect 35176 13028 35180 13084
rect 35180 13028 35236 13084
rect 35236 13028 35240 13084
rect 35176 13024 35240 13028
rect 65656 13084 65720 13088
rect 65656 13028 65660 13084
rect 65660 13028 65716 13084
rect 65716 13028 65720 13084
rect 65656 13024 65720 13028
rect 65736 13084 65800 13088
rect 65736 13028 65740 13084
rect 65740 13028 65796 13084
rect 65796 13028 65800 13084
rect 65736 13024 65800 13028
rect 65816 13084 65880 13088
rect 65816 13028 65820 13084
rect 65820 13028 65876 13084
rect 65876 13028 65880 13084
rect 65816 13024 65880 13028
rect 65896 13084 65960 13088
rect 65896 13028 65900 13084
rect 65900 13028 65956 13084
rect 65956 13028 65960 13084
rect 65896 13024 65960 13028
rect 96376 13084 96440 13088
rect 96376 13028 96380 13084
rect 96380 13028 96436 13084
rect 96436 13028 96440 13084
rect 96376 13024 96440 13028
rect 96456 13084 96520 13088
rect 96456 13028 96460 13084
rect 96460 13028 96516 13084
rect 96516 13028 96520 13084
rect 96456 13024 96520 13028
rect 96536 13084 96600 13088
rect 96536 13028 96540 13084
rect 96540 13028 96596 13084
rect 96596 13028 96600 13084
rect 96536 13024 96600 13028
rect 96616 13084 96680 13088
rect 96616 13028 96620 13084
rect 96620 13028 96676 13084
rect 96676 13028 96680 13084
rect 96616 13024 96680 13028
rect 127096 13084 127160 13088
rect 127096 13028 127100 13084
rect 127100 13028 127156 13084
rect 127156 13028 127160 13084
rect 127096 13024 127160 13028
rect 127176 13084 127240 13088
rect 127176 13028 127180 13084
rect 127180 13028 127236 13084
rect 127236 13028 127240 13084
rect 127176 13024 127240 13028
rect 127256 13084 127320 13088
rect 127256 13028 127260 13084
rect 127260 13028 127316 13084
rect 127316 13028 127320 13084
rect 127256 13024 127320 13028
rect 127336 13084 127400 13088
rect 127336 13028 127340 13084
rect 127340 13028 127396 13084
rect 127396 13028 127400 13084
rect 127336 13024 127400 13028
rect 157816 13084 157880 13088
rect 157816 13028 157820 13084
rect 157820 13028 157876 13084
rect 157876 13028 157880 13084
rect 157816 13024 157880 13028
rect 157896 13084 157960 13088
rect 157896 13028 157900 13084
rect 157900 13028 157956 13084
rect 157956 13028 157960 13084
rect 157896 13024 157960 13028
rect 157976 13084 158040 13088
rect 157976 13028 157980 13084
rect 157980 13028 158036 13084
rect 158036 13028 158040 13084
rect 157976 13024 158040 13028
rect 158056 13084 158120 13088
rect 158056 13028 158060 13084
rect 158060 13028 158116 13084
rect 158116 13028 158120 13084
rect 158056 13024 158120 13028
rect 19576 12540 19640 12544
rect 19576 12484 19580 12540
rect 19580 12484 19636 12540
rect 19636 12484 19640 12540
rect 19576 12480 19640 12484
rect 19656 12540 19720 12544
rect 19656 12484 19660 12540
rect 19660 12484 19716 12540
rect 19716 12484 19720 12540
rect 19656 12480 19720 12484
rect 19736 12540 19800 12544
rect 19736 12484 19740 12540
rect 19740 12484 19796 12540
rect 19796 12484 19800 12540
rect 19736 12480 19800 12484
rect 19816 12540 19880 12544
rect 19816 12484 19820 12540
rect 19820 12484 19876 12540
rect 19876 12484 19880 12540
rect 19816 12480 19880 12484
rect 50296 12540 50360 12544
rect 50296 12484 50300 12540
rect 50300 12484 50356 12540
rect 50356 12484 50360 12540
rect 50296 12480 50360 12484
rect 50376 12540 50440 12544
rect 50376 12484 50380 12540
rect 50380 12484 50436 12540
rect 50436 12484 50440 12540
rect 50376 12480 50440 12484
rect 50456 12540 50520 12544
rect 50456 12484 50460 12540
rect 50460 12484 50516 12540
rect 50516 12484 50520 12540
rect 50456 12480 50520 12484
rect 50536 12540 50600 12544
rect 50536 12484 50540 12540
rect 50540 12484 50596 12540
rect 50596 12484 50600 12540
rect 50536 12480 50600 12484
rect 81016 12540 81080 12544
rect 81016 12484 81020 12540
rect 81020 12484 81076 12540
rect 81076 12484 81080 12540
rect 81016 12480 81080 12484
rect 81096 12540 81160 12544
rect 81096 12484 81100 12540
rect 81100 12484 81156 12540
rect 81156 12484 81160 12540
rect 81096 12480 81160 12484
rect 81176 12540 81240 12544
rect 81176 12484 81180 12540
rect 81180 12484 81236 12540
rect 81236 12484 81240 12540
rect 81176 12480 81240 12484
rect 81256 12540 81320 12544
rect 81256 12484 81260 12540
rect 81260 12484 81316 12540
rect 81316 12484 81320 12540
rect 81256 12480 81320 12484
rect 111736 12540 111800 12544
rect 111736 12484 111740 12540
rect 111740 12484 111796 12540
rect 111796 12484 111800 12540
rect 111736 12480 111800 12484
rect 111816 12540 111880 12544
rect 111816 12484 111820 12540
rect 111820 12484 111876 12540
rect 111876 12484 111880 12540
rect 111816 12480 111880 12484
rect 111896 12540 111960 12544
rect 111896 12484 111900 12540
rect 111900 12484 111956 12540
rect 111956 12484 111960 12540
rect 111896 12480 111960 12484
rect 111976 12540 112040 12544
rect 111976 12484 111980 12540
rect 111980 12484 112036 12540
rect 112036 12484 112040 12540
rect 111976 12480 112040 12484
rect 142456 12540 142520 12544
rect 142456 12484 142460 12540
rect 142460 12484 142516 12540
rect 142516 12484 142520 12540
rect 142456 12480 142520 12484
rect 142536 12540 142600 12544
rect 142536 12484 142540 12540
rect 142540 12484 142596 12540
rect 142596 12484 142600 12540
rect 142536 12480 142600 12484
rect 142616 12540 142680 12544
rect 142616 12484 142620 12540
rect 142620 12484 142676 12540
rect 142676 12484 142680 12540
rect 142616 12480 142680 12484
rect 142696 12540 142760 12544
rect 142696 12484 142700 12540
rect 142700 12484 142756 12540
rect 142756 12484 142760 12540
rect 142696 12480 142760 12484
rect 173176 12540 173240 12544
rect 173176 12484 173180 12540
rect 173180 12484 173236 12540
rect 173236 12484 173240 12540
rect 173176 12480 173240 12484
rect 173256 12540 173320 12544
rect 173256 12484 173260 12540
rect 173260 12484 173316 12540
rect 173316 12484 173320 12540
rect 173256 12480 173320 12484
rect 173336 12540 173400 12544
rect 173336 12484 173340 12540
rect 173340 12484 173396 12540
rect 173396 12484 173400 12540
rect 173336 12480 173400 12484
rect 173416 12540 173480 12544
rect 173416 12484 173420 12540
rect 173420 12484 173476 12540
rect 173476 12484 173480 12540
rect 173416 12480 173480 12484
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 34936 11996 35000 12000
rect 34936 11940 34940 11996
rect 34940 11940 34996 11996
rect 34996 11940 35000 11996
rect 34936 11936 35000 11940
rect 35016 11996 35080 12000
rect 35016 11940 35020 11996
rect 35020 11940 35076 11996
rect 35076 11940 35080 11996
rect 35016 11936 35080 11940
rect 35096 11996 35160 12000
rect 35096 11940 35100 11996
rect 35100 11940 35156 11996
rect 35156 11940 35160 11996
rect 35096 11936 35160 11940
rect 35176 11996 35240 12000
rect 35176 11940 35180 11996
rect 35180 11940 35236 11996
rect 35236 11940 35240 11996
rect 35176 11936 35240 11940
rect 65656 11996 65720 12000
rect 65656 11940 65660 11996
rect 65660 11940 65716 11996
rect 65716 11940 65720 11996
rect 65656 11936 65720 11940
rect 65736 11996 65800 12000
rect 65736 11940 65740 11996
rect 65740 11940 65796 11996
rect 65796 11940 65800 11996
rect 65736 11936 65800 11940
rect 65816 11996 65880 12000
rect 65816 11940 65820 11996
rect 65820 11940 65876 11996
rect 65876 11940 65880 11996
rect 65816 11936 65880 11940
rect 65896 11996 65960 12000
rect 65896 11940 65900 11996
rect 65900 11940 65956 11996
rect 65956 11940 65960 11996
rect 65896 11936 65960 11940
rect 96376 11996 96440 12000
rect 96376 11940 96380 11996
rect 96380 11940 96436 11996
rect 96436 11940 96440 11996
rect 96376 11936 96440 11940
rect 96456 11996 96520 12000
rect 96456 11940 96460 11996
rect 96460 11940 96516 11996
rect 96516 11940 96520 11996
rect 96456 11936 96520 11940
rect 96536 11996 96600 12000
rect 96536 11940 96540 11996
rect 96540 11940 96596 11996
rect 96596 11940 96600 11996
rect 96536 11936 96600 11940
rect 96616 11996 96680 12000
rect 96616 11940 96620 11996
rect 96620 11940 96676 11996
rect 96676 11940 96680 11996
rect 96616 11936 96680 11940
rect 127096 11996 127160 12000
rect 127096 11940 127100 11996
rect 127100 11940 127156 11996
rect 127156 11940 127160 11996
rect 127096 11936 127160 11940
rect 127176 11996 127240 12000
rect 127176 11940 127180 11996
rect 127180 11940 127236 11996
rect 127236 11940 127240 11996
rect 127176 11936 127240 11940
rect 127256 11996 127320 12000
rect 127256 11940 127260 11996
rect 127260 11940 127316 11996
rect 127316 11940 127320 11996
rect 127256 11936 127320 11940
rect 127336 11996 127400 12000
rect 127336 11940 127340 11996
rect 127340 11940 127396 11996
rect 127396 11940 127400 11996
rect 127336 11936 127400 11940
rect 157816 11996 157880 12000
rect 157816 11940 157820 11996
rect 157820 11940 157876 11996
rect 157876 11940 157880 11996
rect 157816 11936 157880 11940
rect 157896 11996 157960 12000
rect 157896 11940 157900 11996
rect 157900 11940 157956 11996
rect 157956 11940 157960 11996
rect 157896 11936 157960 11940
rect 157976 11996 158040 12000
rect 157976 11940 157980 11996
rect 157980 11940 158036 11996
rect 158036 11940 158040 11996
rect 157976 11936 158040 11940
rect 158056 11996 158120 12000
rect 158056 11940 158060 11996
rect 158060 11940 158116 11996
rect 158116 11940 158120 11996
rect 158056 11936 158120 11940
rect 19576 11452 19640 11456
rect 19576 11396 19580 11452
rect 19580 11396 19636 11452
rect 19636 11396 19640 11452
rect 19576 11392 19640 11396
rect 19656 11452 19720 11456
rect 19656 11396 19660 11452
rect 19660 11396 19716 11452
rect 19716 11396 19720 11452
rect 19656 11392 19720 11396
rect 19736 11452 19800 11456
rect 19736 11396 19740 11452
rect 19740 11396 19796 11452
rect 19796 11396 19800 11452
rect 19736 11392 19800 11396
rect 19816 11452 19880 11456
rect 19816 11396 19820 11452
rect 19820 11396 19876 11452
rect 19876 11396 19880 11452
rect 19816 11392 19880 11396
rect 50296 11452 50360 11456
rect 50296 11396 50300 11452
rect 50300 11396 50356 11452
rect 50356 11396 50360 11452
rect 50296 11392 50360 11396
rect 50376 11452 50440 11456
rect 50376 11396 50380 11452
rect 50380 11396 50436 11452
rect 50436 11396 50440 11452
rect 50376 11392 50440 11396
rect 50456 11452 50520 11456
rect 50456 11396 50460 11452
rect 50460 11396 50516 11452
rect 50516 11396 50520 11452
rect 50456 11392 50520 11396
rect 50536 11452 50600 11456
rect 50536 11396 50540 11452
rect 50540 11396 50596 11452
rect 50596 11396 50600 11452
rect 50536 11392 50600 11396
rect 81016 11452 81080 11456
rect 81016 11396 81020 11452
rect 81020 11396 81076 11452
rect 81076 11396 81080 11452
rect 81016 11392 81080 11396
rect 81096 11452 81160 11456
rect 81096 11396 81100 11452
rect 81100 11396 81156 11452
rect 81156 11396 81160 11452
rect 81096 11392 81160 11396
rect 81176 11452 81240 11456
rect 81176 11396 81180 11452
rect 81180 11396 81236 11452
rect 81236 11396 81240 11452
rect 81176 11392 81240 11396
rect 81256 11452 81320 11456
rect 81256 11396 81260 11452
rect 81260 11396 81316 11452
rect 81316 11396 81320 11452
rect 81256 11392 81320 11396
rect 111736 11452 111800 11456
rect 111736 11396 111740 11452
rect 111740 11396 111796 11452
rect 111796 11396 111800 11452
rect 111736 11392 111800 11396
rect 111816 11452 111880 11456
rect 111816 11396 111820 11452
rect 111820 11396 111876 11452
rect 111876 11396 111880 11452
rect 111816 11392 111880 11396
rect 111896 11452 111960 11456
rect 111896 11396 111900 11452
rect 111900 11396 111956 11452
rect 111956 11396 111960 11452
rect 111896 11392 111960 11396
rect 111976 11452 112040 11456
rect 111976 11396 111980 11452
rect 111980 11396 112036 11452
rect 112036 11396 112040 11452
rect 111976 11392 112040 11396
rect 142456 11452 142520 11456
rect 142456 11396 142460 11452
rect 142460 11396 142516 11452
rect 142516 11396 142520 11452
rect 142456 11392 142520 11396
rect 142536 11452 142600 11456
rect 142536 11396 142540 11452
rect 142540 11396 142596 11452
rect 142596 11396 142600 11452
rect 142536 11392 142600 11396
rect 142616 11452 142680 11456
rect 142616 11396 142620 11452
rect 142620 11396 142676 11452
rect 142676 11396 142680 11452
rect 142616 11392 142680 11396
rect 142696 11452 142760 11456
rect 142696 11396 142700 11452
rect 142700 11396 142756 11452
rect 142756 11396 142760 11452
rect 142696 11392 142760 11396
rect 173176 11452 173240 11456
rect 173176 11396 173180 11452
rect 173180 11396 173236 11452
rect 173236 11396 173240 11452
rect 173176 11392 173240 11396
rect 173256 11452 173320 11456
rect 173256 11396 173260 11452
rect 173260 11396 173316 11452
rect 173316 11396 173320 11452
rect 173256 11392 173320 11396
rect 173336 11452 173400 11456
rect 173336 11396 173340 11452
rect 173340 11396 173396 11452
rect 173396 11396 173400 11452
rect 173336 11392 173400 11396
rect 173416 11452 173480 11456
rect 173416 11396 173420 11452
rect 173420 11396 173476 11452
rect 173476 11396 173480 11452
rect 173416 11392 173480 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 34936 10908 35000 10912
rect 34936 10852 34940 10908
rect 34940 10852 34996 10908
rect 34996 10852 35000 10908
rect 34936 10848 35000 10852
rect 35016 10908 35080 10912
rect 35016 10852 35020 10908
rect 35020 10852 35076 10908
rect 35076 10852 35080 10908
rect 35016 10848 35080 10852
rect 35096 10908 35160 10912
rect 35096 10852 35100 10908
rect 35100 10852 35156 10908
rect 35156 10852 35160 10908
rect 35096 10848 35160 10852
rect 35176 10908 35240 10912
rect 35176 10852 35180 10908
rect 35180 10852 35236 10908
rect 35236 10852 35240 10908
rect 35176 10848 35240 10852
rect 65656 10908 65720 10912
rect 65656 10852 65660 10908
rect 65660 10852 65716 10908
rect 65716 10852 65720 10908
rect 65656 10848 65720 10852
rect 65736 10908 65800 10912
rect 65736 10852 65740 10908
rect 65740 10852 65796 10908
rect 65796 10852 65800 10908
rect 65736 10848 65800 10852
rect 65816 10908 65880 10912
rect 65816 10852 65820 10908
rect 65820 10852 65876 10908
rect 65876 10852 65880 10908
rect 65816 10848 65880 10852
rect 65896 10908 65960 10912
rect 65896 10852 65900 10908
rect 65900 10852 65956 10908
rect 65956 10852 65960 10908
rect 65896 10848 65960 10852
rect 96376 10908 96440 10912
rect 96376 10852 96380 10908
rect 96380 10852 96436 10908
rect 96436 10852 96440 10908
rect 96376 10848 96440 10852
rect 96456 10908 96520 10912
rect 96456 10852 96460 10908
rect 96460 10852 96516 10908
rect 96516 10852 96520 10908
rect 96456 10848 96520 10852
rect 96536 10908 96600 10912
rect 96536 10852 96540 10908
rect 96540 10852 96596 10908
rect 96596 10852 96600 10908
rect 96536 10848 96600 10852
rect 96616 10908 96680 10912
rect 96616 10852 96620 10908
rect 96620 10852 96676 10908
rect 96676 10852 96680 10908
rect 96616 10848 96680 10852
rect 127096 10908 127160 10912
rect 127096 10852 127100 10908
rect 127100 10852 127156 10908
rect 127156 10852 127160 10908
rect 127096 10848 127160 10852
rect 127176 10908 127240 10912
rect 127176 10852 127180 10908
rect 127180 10852 127236 10908
rect 127236 10852 127240 10908
rect 127176 10848 127240 10852
rect 127256 10908 127320 10912
rect 127256 10852 127260 10908
rect 127260 10852 127316 10908
rect 127316 10852 127320 10908
rect 127256 10848 127320 10852
rect 127336 10908 127400 10912
rect 127336 10852 127340 10908
rect 127340 10852 127396 10908
rect 127396 10852 127400 10908
rect 127336 10848 127400 10852
rect 157816 10908 157880 10912
rect 157816 10852 157820 10908
rect 157820 10852 157876 10908
rect 157876 10852 157880 10908
rect 157816 10848 157880 10852
rect 157896 10908 157960 10912
rect 157896 10852 157900 10908
rect 157900 10852 157956 10908
rect 157956 10852 157960 10908
rect 157896 10848 157960 10852
rect 157976 10908 158040 10912
rect 157976 10852 157980 10908
rect 157980 10852 158036 10908
rect 158036 10852 158040 10908
rect 157976 10848 158040 10852
rect 158056 10908 158120 10912
rect 158056 10852 158060 10908
rect 158060 10852 158116 10908
rect 158116 10852 158120 10908
rect 158056 10848 158120 10852
rect 19576 10364 19640 10368
rect 19576 10308 19580 10364
rect 19580 10308 19636 10364
rect 19636 10308 19640 10364
rect 19576 10304 19640 10308
rect 19656 10364 19720 10368
rect 19656 10308 19660 10364
rect 19660 10308 19716 10364
rect 19716 10308 19720 10364
rect 19656 10304 19720 10308
rect 19736 10364 19800 10368
rect 19736 10308 19740 10364
rect 19740 10308 19796 10364
rect 19796 10308 19800 10364
rect 19736 10304 19800 10308
rect 19816 10364 19880 10368
rect 19816 10308 19820 10364
rect 19820 10308 19876 10364
rect 19876 10308 19880 10364
rect 19816 10304 19880 10308
rect 50296 10364 50360 10368
rect 50296 10308 50300 10364
rect 50300 10308 50356 10364
rect 50356 10308 50360 10364
rect 50296 10304 50360 10308
rect 50376 10364 50440 10368
rect 50376 10308 50380 10364
rect 50380 10308 50436 10364
rect 50436 10308 50440 10364
rect 50376 10304 50440 10308
rect 50456 10364 50520 10368
rect 50456 10308 50460 10364
rect 50460 10308 50516 10364
rect 50516 10308 50520 10364
rect 50456 10304 50520 10308
rect 50536 10364 50600 10368
rect 50536 10308 50540 10364
rect 50540 10308 50596 10364
rect 50596 10308 50600 10364
rect 50536 10304 50600 10308
rect 81016 10364 81080 10368
rect 81016 10308 81020 10364
rect 81020 10308 81076 10364
rect 81076 10308 81080 10364
rect 81016 10304 81080 10308
rect 81096 10364 81160 10368
rect 81096 10308 81100 10364
rect 81100 10308 81156 10364
rect 81156 10308 81160 10364
rect 81096 10304 81160 10308
rect 81176 10364 81240 10368
rect 81176 10308 81180 10364
rect 81180 10308 81236 10364
rect 81236 10308 81240 10364
rect 81176 10304 81240 10308
rect 81256 10364 81320 10368
rect 81256 10308 81260 10364
rect 81260 10308 81316 10364
rect 81316 10308 81320 10364
rect 81256 10304 81320 10308
rect 111736 10364 111800 10368
rect 111736 10308 111740 10364
rect 111740 10308 111796 10364
rect 111796 10308 111800 10364
rect 111736 10304 111800 10308
rect 111816 10364 111880 10368
rect 111816 10308 111820 10364
rect 111820 10308 111876 10364
rect 111876 10308 111880 10364
rect 111816 10304 111880 10308
rect 111896 10364 111960 10368
rect 111896 10308 111900 10364
rect 111900 10308 111956 10364
rect 111956 10308 111960 10364
rect 111896 10304 111960 10308
rect 111976 10364 112040 10368
rect 111976 10308 111980 10364
rect 111980 10308 112036 10364
rect 112036 10308 112040 10364
rect 111976 10304 112040 10308
rect 142456 10364 142520 10368
rect 142456 10308 142460 10364
rect 142460 10308 142516 10364
rect 142516 10308 142520 10364
rect 142456 10304 142520 10308
rect 142536 10364 142600 10368
rect 142536 10308 142540 10364
rect 142540 10308 142596 10364
rect 142596 10308 142600 10364
rect 142536 10304 142600 10308
rect 142616 10364 142680 10368
rect 142616 10308 142620 10364
rect 142620 10308 142676 10364
rect 142676 10308 142680 10364
rect 142616 10304 142680 10308
rect 142696 10364 142760 10368
rect 142696 10308 142700 10364
rect 142700 10308 142756 10364
rect 142756 10308 142760 10364
rect 142696 10304 142760 10308
rect 173176 10364 173240 10368
rect 173176 10308 173180 10364
rect 173180 10308 173236 10364
rect 173236 10308 173240 10364
rect 173176 10304 173240 10308
rect 173256 10364 173320 10368
rect 173256 10308 173260 10364
rect 173260 10308 173316 10364
rect 173316 10308 173320 10364
rect 173256 10304 173320 10308
rect 173336 10364 173400 10368
rect 173336 10308 173340 10364
rect 173340 10308 173396 10364
rect 173396 10308 173400 10364
rect 173336 10304 173400 10308
rect 173416 10364 173480 10368
rect 173416 10308 173420 10364
rect 173420 10308 173476 10364
rect 173476 10308 173480 10364
rect 173416 10304 173480 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 34936 9820 35000 9824
rect 34936 9764 34940 9820
rect 34940 9764 34996 9820
rect 34996 9764 35000 9820
rect 34936 9760 35000 9764
rect 35016 9820 35080 9824
rect 35016 9764 35020 9820
rect 35020 9764 35076 9820
rect 35076 9764 35080 9820
rect 35016 9760 35080 9764
rect 35096 9820 35160 9824
rect 35096 9764 35100 9820
rect 35100 9764 35156 9820
rect 35156 9764 35160 9820
rect 35096 9760 35160 9764
rect 35176 9820 35240 9824
rect 35176 9764 35180 9820
rect 35180 9764 35236 9820
rect 35236 9764 35240 9820
rect 35176 9760 35240 9764
rect 65656 9820 65720 9824
rect 65656 9764 65660 9820
rect 65660 9764 65716 9820
rect 65716 9764 65720 9820
rect 65656 9760 65720 9764
rect 65736 9820 65800 9824
rect 65736 9764 65740 9820
rect 65740 9764 65796 9820
rect 65796 9764 65800 9820
rect 65736 9760 65800 9764
rect 65816 9820 65880 9824
rect 65816 9764 65820 9820
rect 65820 9764 65876 9820
rect 65876 9764 65880 9820
rect 65816 9760 65880 9764
rect 65896 9820 65960 9824
rect 65896 9764 65900 9820
rect 65900 9764 65956 9820
rect 65956 9764 65960 9820
rect 65896 9760 65960 9764
rect 96376 9820 96440 9824
rect 96376 9764 96380 9820
rect 96380 9764 96436 9820
rect 96436 9764 96440 9820
rect 96376 9760 96440 9764
rect 96456 9820 96520 9824
rect 96456 9764 96460 9820
rect 96460 9764 96516 9820
rect 96516 9764 96520 9820
rect 96456 9760 96520 9764
rect 96536 9820 96600 9824
rect 96536 9764 96540 9820
rect 96540 9764 96596 9820
rect 96596 9764 96600 9820
rect 96536 9760 96600 9764
rect 96616 9820 96680 9824
rect 96616 9764 96620 9820
rect 96620 9764 96676 9820
rect 96676 9764 96680 9820
rect 96616 9760 96680 9764
rect 127096 9820 127160 9824
rect 127096 9764 127100 9820
rect 127100 9764 127156 9820
rect 127156 9764 127160 9820
rect 127096 9760 127160 9764
rect 127176 9820 127240 9824
rect 127176 9764 127180 9820
rect 127180 9764 127236 9820
rect 127236 9764 127240 9820
rect 127176 9760 127240 9764
rect 127256 9820 127320 9824
rect 127256 9764 127260 9820
rect 127260 9764 127316 9820
rect 127316 9764 127320 9820
rect 127256 9760 127320 9764
rect 127336 9820 127400 9824
rect 127336 9764 127340 9820
rect 127340 9764 127396 9820
rect 127396 9764 127400 9820
rect 127336 9760 127400 9764
rect 157816 9820 157880 9824
rect 157816 9764 157820 9820
rect 157820 9764 157876 9820
rect 157876 9764 157880 9820
rect 157816 9760 157880 9764
rect 157896 9820 157960 9824
rect 157896 9764 157900 9820
rect 157900 9764 157956 9820
rect 157956 9764 157960 9820
rect 157896 9760 157960 9764
rect 157976 9820 158040 9824
rect 157976 9764 157980 9820
rect 157980 9764 158036 9820
rect 158036 9764 158040 9820
rect 157976 9760 158040 9764
rect 158056 9820 158120 9824
rect 158056 9764 158060 9820
rect 158060 9764 158116 9820
rect 158116 9764 158120 9820
rect 158056 9760 158120 9764
rect 19576 9276 19640 9280
rect 19576 9220 19580 9276
rect 19580 9220 19636 9276
rect 19636 9220 19640 9276
rect 19576 9216 19640 9220
rect 19656 9276 19720 9280
rect 19656 9220 19660 9276
rect 19660 9220 19716 9276
rect 19716 9220 19720 9276
rect 19656 9216 19720 9220
rect 19736 9276 19800 9280
rect 19736 9220 19740 9276
rect 19740 9220 19796 9276
rect 19796 9220 19800 9276
rect 19736 9216 19800 9220
rect 19816 9276 19880 9280
rect 19816 9220 19820 9276
rect 19820 9220 19876 9276
rect 19876 9220 19880 9276
rect 19816 9216 19880 9220
rect 50296 9276 50360 9280
rect 50296 9220 50300 9276
rect 50300 9220 50356 9276
rect 50356 9220 50360 9276
rect 50296 9216 50360 9220
rect 50376 9276 50440 9280
rect 50376 9220 50380 9276
rect 50380 9220 50436 9276
rect 50436 9220 50440 9276
rect 50376 9216 50440 9220
rect 50456 9276 50520 9280
rect 50456 9220 50460 9276
rect 50460 9220 50516 9276
rect 50516 9220 50520 9276
rect 50456 9216 50520 9220
rect 50536 9276 50600 9280
rect 50536 9220 50540 9276
rect 50540 9220 50596 9276
rect 50596 9220 50600 9276
rect 50536 9216 50600 9220
rect 81016 9276 81080 9280
rect 81016 9220 81020 9276
rect 81020 9220 81076 9276
rect 81076 9220 81080 9276
rect 81016 9216 81080 9220
rect 81096 9276 81160 9280
rect 81096 9220 81100 9276
rect 81100 9220 81156 9276
rect 81156 9220 81160 9276
rect 81096 9216 81160 9220
rect 81176 9276 81240 9280
rect 81176 9220 81180 9276
rect 81180 9220 81236 9276
rect 81236 9220 81240 9276
rect 81176 9216 81240 9220
rect 81256 9276 81320 9280
rect 81256 9220 81260 9276
rect 81260 9220 81316 9276
rect 81316 9220 81320 9276
rect 81256 9216 81320 9220
rect 111736 9276 111800 9280
rect 111736 9220 111740 9276
rect 111740 9220 111796 9276
rect 111796 9220 111800 9276
rect 111736 9216 111800 9220
rect 111816 9276 111880 9280
rect 111816 9220 111820 9276
rect 111820 9220 111876 9276
rect 111876 9220 111880 9276
rect 111816 9216 111880 9220
rect 111896 9276 111960 9280
rect 111896 9220 111900 9276
rect 111900 9220 111956 9276
rect 111956 9220 111960 9276
rect 111896 9216 111960 9220
rect 111976 9276 112040 9280
rect 111976 9220 111980 9276
rect 111980 9220 112036 9276
rect 112036 9220 112040 9276
rect 111976 9216 112040 9220
rect 142456 9276 142520 9280
rect 142456 9220 142460 9276
rect 142460 9220 142516 9276
rect 142516 9220 142520 9276
rect 142456 9216 142520 9220
rect 142536 9276 142600 9280
rect 142536 9220 142540 9276
rect 142540 9220 142596 9276
rect 142596 9220 142600 9276
rect 142536 9216 142600 9220
rect 142616 9276 142680 9280
rect 142616 9220 142620 9276
rect 142620 9220 142676 9276
rect 142676 9220 142680 9276
rect 142616 9216 142680 9220
rect 142696 9276 142760 9280
rect 142696 9220 142700 9276
rect 142700 9220 142756 9276
rect 142756 9220 142760 9276
rect 142696 9216 142760 9220
rect 173176 9276 173240 9280
rect 173176 9220 173180 9276
rect 173180 9220 173236 9276
rect 173236 9220 173240 9276
rect 173176 9216 173240 9220
rect 173256 9276 173320 9280
rect 173256 9220 173260 9276
rect 173260 9220 173316 9276
rect 173316 9220 173320 9276
rect 173256 9216 173320 9220
rect 173336 9276 173400 9280
rect 173336 9220 173340 9276
rect 173340 9220 173396 9276
rect 173396 9220 173400 9276
rect 173336 9216 173400 9220
rect 173416 9276 173480 9280
rect 173416 9220 173420 9276
rect 173420 9220 173476 9276
rect 173476 9220 173480 9276
rect 173416 9216 173480 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 34936 8732 35000 8736
rect 34936 8676 34940 8732
rect 34940 8676 34996 8732
rect 34996 8676 35000 8732
rect 34936 8672 35000 8676
rect 35016 8732 35080 8736
rect 35016 8676 35020 8732
rect 35020 8676 35076 8732
rect 35076 8676 35080 8732
rect 35016 8672 35080 8676
rect 35096 8732 35160 8736
rect 35096 8676 35100 8732
rect 35100 8676 35156 8732
rect 35156 8676 35160 8732
rect 35096 8672 35160 8676
rect 35176 8732 35240 8736
rect 35176 8676 35180 8732
rect 35180 8676 35236 8732
rect 35236 8676 35240 8732
rect 35176 8672 35240 8676
rect 65656 8732 65720 8736
rect 65656 8676 65660 8732
rect 65660 8676 65716 8732
rect 65716 8676 65720 8732
rect 65656 8672 65720 8676
rect 65736 8732 65800 8736
rect 65736 8676 65740 8732
rect 65740 8676 65796 8732
rect 65796 8676 65800 8732
rect 65736 8672 65800 8676
rect 65816 8732 65880 8736
rect 65816 8676 65820 8732
rect 65820 8676 65876 8732
rect 65876 8676 65880 8732
rect 65816 8672 65880 8676
rect 65896 8732 65960 8736
rect 65896 8676 65900 8732
rect 65900 8676 65956 8732
rect 65956 8676 65960 8732
rect 65896 8672 65960 8676
rect 96376 8732 96440 8736
rect 96376 8676 96380 8732
rect 96380 8676 96436 8732
rect 96436 8676 96440 8732
rect 96376 8672 96440 8676
rect 96456 8732 96520 8736
rect 96456 8676 96460 8732
rect 96460 8676 96516 8732
rect 96516 8676 96520 8732
rect 96456 8672 96520 8676
rect 96536 8732 96600 8736
rect 96536 8676 96540 8732
rect 96540 8676 96596 8732
rect 96596 8676 96600 8732
rect 96536 8672 96600 8676
rect 96616 8732 96680 8736
rect 96616 8676 96620 8732
rect 96620 8676 96676 8732
rect 96676 8676 96680 8732
rect 96616 8672 96680 8676
rect 127096 8732 127160 8736
rect 127096 8676 127100 8732
rect 127100 8676 127156 8732
rect 127156 8676 127160 8732
rect 127096 8672 127160 8676
rect 127176 8732 127240 8736
rect 127176 8676 127180 8732
rect 127180 8676 127236 8732
rect 127236 8676 127240 8732
rect 127176 8672 127240 8676
rect 127256 8732 127320 8736
rect 127256 8676 127260 8732
rect 127260 8676 127316 8732
rect 127316 8676 127320 8732
rect 127256 8672 127320 8676
rect 127336 8732 127400 8736
rect 127336 8676 127340 8732
rect 127340 8676 127396 8732
rect 127396 8676 127400 8732
rect 127336 8672 127400 8676
rect 157816 8732 157880 8736
rect 157816 8676 157820 8732
rect 157820 8676 157876 8732
rect 157876 8676 157880 8732
rect 157816 8672 157880 8676
rect 157896 8732 157960 8736
rect 157896 8676 157900 8732
rect 157900 8676 157956 8732
rect 157956 8676 157960 8732
rect 157896 8672 157960 8676
rect 157976 8732 158040 8736
rect 157976 8676 157980 8732
rect 157980 8676 158036 8732
rect 158036 8676 158040 8732
rect 157976 8672 158040 8676
rect 158056 8732 158120 8736
rect 158056 8676 158060 8732
rect 158060 8676 158116 8732
rect 158116 8676 158120 8732
rect 158056 8672 158120 8676
rect 19576 8188 19640 8192
rect 19576 8132 19580 8188
rect 19580 8132 19636 8188
rect 19636 8132 19640 8188
rect 19576 8128 19640 8132
rect 19656 8188 19720 8192
rect 19656 8132 19660 8188
rect 19660 8132 19716 8188
rect 19716 8132 19720 8188
rect 19656 8128 19720 8132
rect 19736 8188 19800 8192
rect 19736 8132 19740 8188
rect 19740 8132 19796 8188
rect 19796 8132 19800 8188
rect 19736 8128 19800 8132
rect 19816 8188 19880 8192
rect 19816 8132 19820 8188
rect 19820 8132 19876 8188
rect 19876 8132 19880 8188
rect 19816 8128 19880 8132
rect 50296 8188 50360 8192
rect 50296 8132 50300 8188
rect 50300 8132 50356 8188
rect 50356 8132 50360 8188
rect 50296 8128 50360 8132
rect 50376 8188 50440 8192
rect 50376 8132 50380 8188
rect 50380 8132 50436 8188
rect 50436 8132 50440 8188
rect 50376 8128 50440 8132
rect 50456 8188 50520 8192
rect 50456 8132 50460 8188
rect 50460 8132 50516 8188
rect 50516 8132 50520 8188
rect 50456 8128 50520 8132
rect 50536 8188 50600 8192
rect 50536 8132 50540 8188
rect 50540 8132 50596 8188
rect 50596 8132 50600 8188
rect 50536 8128 50600 8132
rect 81016 8188 81080 8192
rect 81016 8132 81020 8188
rect 81020 8132 81076 8188
rect 81076 8132 81080 8188
rect 81016 8128 81080 8132
rect 81096 8188 81160 8192
rect 81096 8132 81100 8188
rect 81100 8132 81156 8188
rect 81156 8132 81160 8188
rect 81096 8128 81160 8132
rect 81176 8188 81240 8192
rect 81176 8132 81180 8188
rect 81180 8132 81236 8188
rect 81236 8132 81240 8188
rect 81176 8128 81240 8132
rect 81256 8188 81320 8192
rect 81256 8132 81260 8188
rect 81260 8132 81316 8188
rect 81316 8132 81320 8188
rect 81256 8128 81320 8132
rect 111736 8188 111800 8192
rect 111736 8132 111740 8188
rect 111740 8132 111796 8188
rect 111796 8132 111800 8188
rect 111736 8128 111800 8132
rect 111816 8188 111880 8192
rect 111816 8132 111820 8188
rect 111820 8132 111876 8188
rect 111876 8132 111880 8188
rect 111816 8128 111880 8132
rect 111896 8188 111960 8192
rect 111896 8132 111900 8188
rect 111900 8132 111956 8188
rect 111956 8132 111960 8188
rect 111896 8128 111960 8132
rect 111976 8188 112040 8192
rect 111976 8132 111980 8188
rect 111980 8132 112036 8188
rect 112036 8132 112040 8188
rect 111976 8128 112040 8132
rect 142456 8188 142520 8192
rect 142456 8132 142460 8188
rect 142460 8132 142516 8188
rect 142516 8132 142520 8188
rect 142456 8128 142520 8132
rect 142536 8188 142600 8192
rect 142536 8132 142540 8188
rect 142540 8132 142596 8188
rect 142596 8132 142600 8188
rect 142536 8128 142600 8132
rect 142616 8188 142680 8192
rect 142616 8132 142620 8188
rect 142620 8132 142676 8188
rect 142676 8132 142680 8188
rect 142616 8128 142680 8132
rect 142696 8188 142760 8192
rect 142696 8132 142700 8188
rect 142700 8132 142756 8188
rect 142756 8132 142760 8188
rect 142696 8128 142760 8132
rect 173176 8188 173240 8192
rect 173176 8132 173180 8188
rect 173180 8132 173236 8188
rect 173236 8132 173240 8188
rect 173176 8128 173240 8132
rect 173256 8188 173320 8192
rect 173256 8132 173260 8188
rect 173260 8132 173316 8188
rect 173316 8132 173320 8188
rect 173256 8128 173320 8132
rect 173336 8188 173400 8192
rect 173336 8132 173340 8188
rect 173340 8132 173396 8188
rect 173396 8132 173400 8188
rect 173336 8128 173400 8132
rect 173416 8188 173480 8192
rect 173416 8132 173420 8188
rect 173420 8132 173476 8188
rect 173476 8132 173480 8188
rect 173416 8128 173480 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 34936 7644 35000 7648
rect 34936 7588 34940 7644
rect 34940 7588 34996 7644
rect 34996 7588 35000 7644
rect 34936 7584 35000 7588
rect 35016 7644 35080 7648
rect 35016 7588 35020 7644
rect 35020 7588 35076 7644
rect 35076 7588 35080 7644
rect 35016 7584 35080 7588
rect 35096 7644 35160 7648
rect 35096 7588 35100 7644
rect 35100 7588 35156 7644
rect 35156 7588 35160 7644
rect 35096 7584 35160 7588
rect 35176 7644 35240 7648
rect 35176 7588 35180 7644
rect 35180 7588 35236 7644
rect 35236 7588 35240 7644
rect 35176 7584 35240 7588
rect 65656 7644 65720 7648
rect 65656 7588 65660 7644
rect 65660 7588 65716 7644
rect 65716 7588 65720 7644
rect 65656 7584 65720 7588
rect 65736 7644 65800 7648
rect 65736 7588 65740 7644
rect 65740 7588 65796 7644
rect 65796 7588 65800 7644
rect 65736 7584 65800 7588
rect 65816 7644 65880 7648
rect 65816 7588 65820 7644
rect 65820 7588 65876 7644
rect 65876 7588 65880 7644
rect 65816 7584 65880 7588
rect 65896 7644 65960 7648
rect 65896 7588 65900 7644
rect 65900 7588 65956 7644
rect 65956 7588 65960 7644
rect 65896 7584 65960 7588
rect 96376 7644 96440 7648
rect 96376 7588 96380 7644
rect 96380 7588 96436 7644
rect 96436 7588 96440 7644
rect 96376 7584 96440 7588
rect 96456 7644 96520 7648
rect 96456 7588 96460 7644
rect 96460 7588 96516 7644
rect 96516 7588 96520 7644
rect 96456 7584 96520 7588
rect 96536 7644 96600 7648
rect 96536 7588 96540 7644
rect 96540 7588 96596 7644
rect 96596 7588 96600 7644
rect 96536 7584 96600 7588
rect 96616 7644 96680 7648
rect 96616 7588 96620 7644
rect 96620 7588 96676 7644
rect 96676 7588 96680 7644
rect 96616 7584 96680 7588
rect 127096 7644 127160 7648
rect 127096 7588 127100 7644
rect 127100 7588 127156 7644
rect 127156 7588 127160 7644
rect 127096 7584 127160 7588
rect 127176 7644 127240 7648
rect 127176 7588 127180 7644
rect 127180 7588 127236 7644
rect 127236 7588 127240 7644
rect 127176 7584 127240 7588
rect 127256 7644 127320 7648
rect 127256 7588 127260 7644
rect 127260 7588 127316 7644
rect 127316 7588 127320 7644
rect 127256 7584 127320 7588
rect 127336 7644 127400 7648
rect 127336 7588 127340 7644
rect 127340 7588 127396 7644
rect 127396 7588 127400 7644
rect 127336 7584 127400 7588
rect 157816 7644 157880 7648
rect 157816 7588 157820 7644
rect 157820 7588 157876 7644
rect 157876 7588 157880 7644
rect 157816 7584 157880 7588
rect 157896 7644 157960 7648
rect 157896 7588 157900 7644
rect 157900 7588 157956 7644
rect 157956 7588 157960 7644
rect 157896 7584 157960 7588
rect 157976 7644 158040 7648
rect 157976 7588 157980 7644
rect 157980 7588 158036 7644
rect 158036 7588 158040 7644
rect 157976 7584 158040 7588
rect 158056 7644 158120 7648
rect 158056 7588 158060 7644
rect 158060 7588 158116 7644
rect 158116 7588 158120 7644
rect 158056 7584 158120 7588
rect 19576 7100 19640 7104
rect 19576 7044 19580 7100
rect 19580 7044 19636 7100
rect 19636 7044 19640 7100
rect 19576 7040 19640 7044
rect 19656 7100 19720 7104
rect 19656 7044 19660 7100
rect 19660 7044 19716 7100
rect 19716 7044 19720 7100
rect 19656 7040 19720 7044
rect 19736 7100 19800 7104
rect 19736 7044 19740 7100
rect 19740 7044 19796 7100
rect 19796 7044 19800 7100
rect 19736 7040 19800 7044
rect 19816 7100 19880 7104
rect 19816 7044 19820 7100
rect 19820 7044 19876 7100
rect 19876 7044 19880 7100
rect 19816 7040 19880 7044
rect 50296 7100 50360 7104
rect 50296 7044 50300 7100
rect 50300 7044 50356 7100
rect 50356 7044 50360 7100
rect 50296 7040 50360 7044
rect 50376 7100 50440 7104
rect 50376 7044 50380 7100
rect 50380 7044 50436 7100
rect 50436 7044 50440 7100
rect 50376 7040 50440 7044
rect 50456 7100 50520 7104
rect 50456 7044 50460 7100
rect 50460 7044 50516 7100
rect 50516 7044 50520 7100
rect 50456 7040 50520 7044
rect 50536 7100 50600 7104
rect 50536 7044 50540 7100
rect 50540 7044 50596 7100
rect 50596 7044 50600 7100
rect 50536 7040 50600 7044
rect 81016 7100 81080 7104
rect 81016 7044 81020 7100
rect 81020 7044 81076 7100
rect 81076 7044 81080 7100
rect 81016 7040 81080 7044
rect 81096 7100 81160 7104
rect 81096 7044 81100 7100
rect 81100 7044 81156 7100
rect 81156 7044 81160 7100
rect 81096 7040 81160 7044
rect 81176 7100 81240 7104
rect 81176 7044 81180 7100
rect 81180 7044 81236 7100
rect 81236 7044 81240 7100
rect 81176 7040 81240 7044
rect 81256 7100 81320 7104
rect 81256 7044 81260 7100
rect 81260 7044 81316 7100
rect 81316 7044 81320 7100
rect 81256 7040 81320 7044
rect 111736 7100 111800 7104
rect 111736 7044 111740 7100
rect 111740 7044 111796 7100
rect 111796 7044 111800 7100
rect 111736 7040 111800 7044
rect 111816 7100 111880 7104
rect 111816 7044 111820 7100
rect 111820 7044 111876 7100
rect 111876 7044 111880 7100
rect 111816 7040 111880 7044
rect 111896 7100 111960 7104
rect 111896 7044 111900 7100
rect 111900 7044 111956 7100
rect 111956 7044 111960 7100
rect 111896 7040 111960 7044
rect 111976 7100 112040 7104
rect 111976 7044 111980 7100
rect 111980 7044 112036 7100
rect 112036 7044 112040 7100
rect 111976 7040 112040 7044
rect 142456 7100 142520 7104
rect 142456 7044 142460 7100
rect 142460 7044 142516 7100
rect 142516 7044 142520 7100
rect 142456 7040 142520 7044
rect 142536 7100 142600 7104
rect 142536 7044 142540 7100
rect 142540 7044 142596 7100
rect 142596 7044 142600 7100
rect 142536 7040 142600 7044
rect 142616 7100 142680 7104
rect 142616 7044 142620 7100
rect 142620 7044 142676 7100
rect 142676 7044 142680 7100
rect 142616 7040 142680 7044
rect 142696 7100 142760 7104
rect 142696 7044 142700 7100
rect 142700 7044 142756 7100
rect 142756 7044 142760 7100
rect 142696 7040 142760 7044
rect 173176 7100 173240 7104
rect 173176 7044 173180 7100
rect 173180 7044 173236 7100
rect 173236 7044 173240 7100
rect 173176 7040 173240 7044
rect 173256 7100 173320 7104
rect 173256 7044 173260 7100
rect 173260 7044 173316 7100
rect 173316 7044 173320 7100
rect 173256 7040 173320 7044
rect 173336 7100 173400 7104
rect 173336 7044 173340 7100
rect 173340 7044 173396 7100
rect 173396 7044 173400 7100
rect 173336 7040 173400 7044
rect 173416 7100 173480 7104
rect 173416 7044 173420 7100
rect 173420 7044 173476 7100
rect 173476 7044 173480 7100
rect 173416 7040 173480 7044
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 34936 6556 35000 6560
rect 34936 6500 34940 6556
rect 34940 6500 34996 6556
rect 34996 6500 35000 6556
rect 34936 6496 35000 6500
rect 35016 6556 35080 6560
rect 35016 6500 35020 6556
rect 35020 6500 35076 6556
rect 35076 6500 35080 6556
rect 35016 6496 35080 6500
rect 35096 6556 35160 6560
rect 35096 6500 35100 6556
rect 35100 6500 35156 6556
rect 35156 6500 35160 6556
rect 35096 6496 35160 6500
rect 35176 6556 35240 6560
rect 35176 6500 35180 6556
rect 35180 6500 35236 6556
rect 35236 6500 35240 6556
rect 35176 6496 35240 6500
rect 65656 6556 65720 6560
rect 65656 6500 65660 6556
rect 65660 6500 65716 6556
rect 65716 6500 65720 6556
rect 65656 6496 65720 6500
rect 65736 6556 65800 6560
rect 65736 6500 65740 6556
rect 65740 6500 65796 6556
rect 65796 6500 65800 6556
rect 65736 6496 65800 6500
rect 65816 6556 65880 6560
rect 65816 6500 65820 6556
rect 65820 6500 65876 6556
rect 65876 6500 65880 6556
rect 65816 6496 65880 6500
rect 65896 6556 65960 6560
rect 65896 6500 65900 6556
rect 65900 6500 65956 6556
rect 65956 6500 65960 6556
rect 65896 6496 65960 6500
rect 96376 6556 96440 6560
rect 96376 6500 96380 6556
rect 96380 6500 96436 6556
rect 96436 6500 96440 6556
rect 96376 6496 96440 6500
rect 96456 6556 96520 6560
rect 96456 6500 96460 6556
rect 96460 6500 96516 6556
rect 96516 6500 96520 6556
rect 96456 6496 96520 6500
rect 96536 6556 96600 6560
rect 96536 6500 96540 6556
rect 96540 6500 96596 6556
rect 96596 6500 96600 6556
rect 96536 6496 96600 6500
rect 96616 6556 96680 6560
rect 96616 6500 96620 6556
rect 96620 6500 96676 6556
rect 96676 6500 96680 6556
rect 96616 6496 96680 6500
rect 127096 6556 127160 6560
rect 127096 6500 127100 6556
rect 127100 6500 127156 6556
rect 127156 6500 127160 6556
rect 127096 6496 127160 6500
rect 127176 6556 127240 6560
rect 127176 6500 127180 6556
rect 127180 6500 127236 6556
rect 127236 6500 127240 6556
rect 127176 6496 127240 6500
rect 127256 6556 127320 6560
rect 127256 6500 127260 6556
rect 127260 6500 127316 6556
rect 127316 6500 127320 6556
rect 127256 6496 127320 6500
rect 127336 6556 127400 6560
rect 127336 6500 127340 6556
rect 127340 6500 127396 6556
rect 127396 6500 127400 6556
rect 127336 6496 127400 6500
rect 157816 6556 157880 6560
rect 157816 6500 157820 6556
rect 157820 6500 157876 6556
rect 157876 6500 157880 6556
rect 157816 6496 157880 6500
rect 157896 6556 157960 6560
rect 157896 6500 157900 6556
rect 157900 6500 157956 6556
rect 157956 6500 157960 6556
rect 157896 6496 157960 6500
rect 157976 6556 158040 6560
rect 157976 6500 157980 6556
rect 157980 6500 158036 6556
rect 158036 6500 158040 6556
rect 157976 6496 158040 6500
rect 158056 6556 158120 6560
rect 158056 6500 158060 6556
rect 158060 6500 158116 6556
rect 158116 6500 158120 6556
rect 158056 6496 158120 6500
rect 19576 6012 19640 6016
rect 19576 5956 19580 6012
rect 19580 5956 19636 6012
rect 19636 5956 19640 6012
rect 19576 5952 19640 5956
rect 19656 6012 19720 6016
rect 19656 5956 19660 6012
rect 19660 5956 19716 6012
rect 19716 5956 19720 6012
rect 19656 5952 19720 5956
rect 19736 6012 19800 6016
rect 19736 5956 19740 6012
rect 19740 5956 19796 6012
rect 19796 5956 19800 6012
rect 19736 5952 19800 5956
rect 19816 6012 19880 6016
rect 19816 5956 19820 6012
rect 19820 5956 19876 6012
rect 19876 5956 19880 6012
rect 19816 5952 19880 5956
rect 50296 6012 50360 6016
rect 50296 5956 50300 6012
rect 50300 5956 50356 6012
rect 50356 5956 50360 6012
rect 50296 5952 50360 5956
rect 50376 6012 50440 6016
rect 50376 5956 50380 6012
rect 50380 5956 50436 6012
rect 50436 5956 50440 6012
rect 50376 5952 50440 5956
rect 50456 6012 50520 6016
rect 50456 5956 50460 6012
rect 50460 5956 50516 6012
rect 50516 5956 50520 6012
rect 50456 5952 50520 5956
rect 50536 6012 50600 6016
rect 50536 5956 50540 6012
rect 50540 5956 50596 6012
rect 50596 5956 50600 6012
rect 50536 5952 50600 5956
rect 81016 6012 81080 6016
rect 81016 5956 81020 6012
rect 81020 5956 81076 6012
rect 81076 5956 81080 6012
rect 81016 5952 81080 5956
rect 81096 6012 81160 6016
rect 81096 5956 81100 6012
rect 81100 5956 81156 6012
rect 81156 5956 81160 6012
rect 81096 5952 81160 5956
rect 81176 6012 81240 6016
rect 81176 5956 81180 6012
rect 81180 5956 81236 6012
rect 81236 5956 81240 6012
rect 81176 5952 81240 5956
rect 81256 6012 81320 6016
rect 81256 5956 81260 6012
rect 81260 5956 81316 6012
rect 81316 5956 81320 6012
rect 81256 5952 81320 5956
rect 111736 6012 111800 6016
rect 111736 5956 111740 6012
rect 111740 5956 111796 6012
rect 111796 5956 111800 6012
rect 111736 5952 111800 5956
rect 111816 6012 111880 6016
rect 111816 5956 111820 6012
rect 111820 5956 111876 6012
rect 111876 5956 111880 6012
rect 111816 5952 111880 5956
rect 111896 6012 111960 6016
rect 111896 5956 111900 6012
rect 111900 5956 111956 6012
rect 111956 5956 111960 6012
rect 111896 5952 111960 5956
rect 111976 6012 112040 6016
rect 111976 5956 111980 6012
rect 111980 5956 112036 6012
rect 112036 5956 112040 6012
rect 111976 5952 112040 5956
rect 142456 6012 142520 6016
rect 142456 5956 142460 6012
rect 142460 5956 142516 6012
rect 142516 5956 142520 6012
rect 142456 5952 142520 5956
rect 142536 6012 142600 6016
rect 142536 5956 142540 6012
rect 142540 5956 142596 6012
rect 142596 5956 142600 6012
rect 142536 5952 142600 5956
rect 142616 6012 142680 6016
rect 142616 5956 142620 6012
rect 142620 5956 142676 6012
rect 142676 5956 142680 6012
rect 142616 5952 142680 5956
rect 142696 6012 142760 6016
rect 142696 5956 142700 6012
rect 142700 5956 142756 6012
rect 142756 5956 142760 6012
rect 142696 5952 142760 5956
rect 173176 6012 173240 6016
rect 173176 5956 173180 6012
rect 173180 5956 173236 6012
rect 173236 5956 173240 6012
rect 173176 5952 173240 5956
rect 173256 6012 173320 6016
rect 173256 5956 173260 6012
rect 173260 5956 173316 6012
rect 173316 5956 173320 6012
rect 173256 5952 173320 5956
rect 173336 6012 173400 6016
rect 173336 5956 173340 6012
rect 173340 5956 173396 6012
rect 173396 5956 173400 6012
rect 173336 5952 173400 5956
rect 173416 6012 173480 6016
rect 173416 5956 173420 6012
rect 173420 5956 173476 6012
rect 173476 5956 173480 6012
rect 173416 5952 173480 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 34936 5468 35000 5472
rect 34936 5412 34940 5468
rect 34940 5412 34996 5468
rect 34996 5412 35000 5468
rect 34936 5408 35000 5412
rect 35016 5468 35080 5472
rect 35016 5412 35020 5468
rect 35020 5412 35076 5468
rect 35076 5412 35080 5468
rect 35016 5408 35080 5412
rect 35096 5468 35160 5472
rect 35096 5412 35100 5468
rect 35100 5412 35156 5468
rect 35156 5412 35160 5468
rect 35096 5408 35160 5412
rect 35176 5468 35240 5472
rect 35176 5412 35180 5468
rect 35180 5412 35236 5468
rect 35236 5412 35240 5468
rect 35176 5408 35240 5412
rect 65656 5468 65720 5472
rect 65656 5412 65660 5468
rect 65660 5412 65716 5468
rect 65716 5412 65720 5468
rect 65656 5408 65720 5412
rect 65736 5468 65800 5472
rect 65736 5412 65740 5468
rect 65740 5412 65796 5468
rect 65796 5412 65800 5468
rect 65736 5408 65800 5412
rect 65816 5468 65880 5472
rect 65816 5412 65820 5468
rect 65820 5412 65876 5468
rect 65876 5412 65880 5468
rect 65816 5408 65880 5412
rect 65896 5468 65960 5472
rect 65896 5412 65900 5468
rect 65900 5412 65956 5468
rect 65956 5412 65960 5468
rect 65896 5408 65960 5412
rect 96376 5468 96440 5472
rect 96376 5412 96380 5468
rect 96380 5412 96436 5468
rect 96436 5412 96440 5468
rect 96376 5408 96440 5412
rect 96456 5468 96520 5472
rect 96456 5412 96460 5468
rect 96460 5412 96516 5468
rect 96516 5412 96520 5468
rect 96456 5408 96520 5412
rect 96536 5468 96600 5472
rect 96536 5412 96540 5468
rect 96540 5412 96596 5468
rect 96596 5412 96600 5468
rect 96536 5408 96600 5412
rect 96616 5468 96680 5472
rect 96616 5412 96620 5468
rect 96620 5412 96676 5468
rect 96676 5412 96680 5468
rect 96616 5408 96680 5412
rect 127096 5468 127160 5472
rect 127096 5412 127100 5468
rect 127100 5412 127156 5468
rect 127156 5412 127160 5468
rect 127096 5408 127160 5412
rect 127176 5468 127240 5472
rect 127176 5412 127180 5468
rect 127180 5412 127236 5468
rect 127236 5412 127240 5468
rect 127176 5408 127240 5412
rect 127256 5468 127320 5472
rect 127256 5412 127260 5468
rect 127260 5412 127316 5468
rect 127316 5412 127320 5468
rect 127256 5408 127320 5412
rect 127336 5468 127400 5472
rect 127336 5412 127340 5468
rect 127340 5412 127396 5468
rect 127396 5412 127400 5468
rect 127336 5408 127400 5412
rect 157816 5468 157880 5472
rect 157816 5412 157820 5468
rect 157820 5412 157876 5468
rect 157876 5412 157880 5468
rect 157816 5408 157880 5412
rect 157896 5468 157960 5472
rect 157896 5412 157900 5468
rect 157900 5412 157956 5468
rect 157956 5412 157960 5468
rect 157896 5408 157960 5412
rect 157976 5468 158040 5472
rect 157976 5412 157980 5468
rect 157980 5412 158036 5468
rect 158036 5412 158040 5468
rect 157976 5408 158040 5412
rect 158056 5468 158120 5472
rect 158056 5412 158060 5468
rect 158060 5412 158116 5468
rect 158116 5412 158120 5468
rect 158056 5408 158120 5412
rect 19576 4924 19640 4928
rect 19576 4868 19580 4924
rect 19580 4868 19636 4924
rect 19636 4868 19640 4924
rect 19576 4864 19640 4868
rect 19656 4924 19720 4928
rect 19656 4868 19660 4924
rect 19660 4868 19716 4924
rect 19716 4868 19720 4924
rect 19656 4864 19720 4868
rect 19736 4924 19800 4928
rect 19736 4868 19740 4924
rect 19740 4868 19796 4924
rect 19796 4868 19800 4924
rect 19736 4864 19800 4868
rect 19816 4924 19880 4928
rect 19816 4868 19820 4924
rect 19820 4868 19876 4924
rect 19876 4868 19880 4924
rect 19816 4864 19880 4868
rect 50296 4924 50360 4928
rect 50296 4868 50300 4924
rect 50300 4868 50356 4924
rect 50356 4868 50360 4924
rect 50296 4864 50360 4868
rect 50376 4924 50440 4928
rect 50376 4868 50380 4924
rect 50380 4868 50436 4924
rect 50436 4868 50440 4924
rect 50376 4864 50440 4868
rect 50456 4924 50520 4928
rect 50456 4868 50460 4924
rect 50460 4868 50516 4924
rect 50516 4868 50520 4924
rect 50456 4864 50520 4868
rect 50536 4924 50600 4928
rect 50536 4868 50540 4924
rect 50540 4868 50596 4924
rect 50596 4868 50600 4924
rect 50536 4864 50600 4868
rect 81016 4924 81080 4928
rect 81016 4868 81020 4924
rect 81020 4868 81076 4924
rect 81076 4868 81080 4924
rect 81016 4864 81080 4868
rect 81096 4924 81160 4928
rect 81096 4868 81100 4924
rect 81100 4868 81156 4924
rect 81156 4868 81160 4924
rect 81096 4864 81160 4868
rect 81176 4924 81240 4928
rect 81176 4868 81180 4924
rect 81180 4868 81236 4924
rect 81236 4868 81240 4924
rect 81176 4864 81240 4868
rect 81256 4924 81320 4928
rect 81256 4868 81260 4924
rect 81260 4868 81316 4924
rect 81316 4868 81320 4924
rect 81256 4864 81320 4868
rect 111736 4924 111800 4928
rect 111736 4868 111740 4924
rect 111740 4868 111796 4924
rect 111796 4868 111800 4924
rect 111736 4864 111800 4868
rect 111816 4924 111880 4928
rect 111816 4868 111820 4924
rect 111820 4868 111876 4924
rect 111876 4868 111880 4924
rect 111816 4864 111880 4868
rect 111896 4924 111960 4928
rect 111896 4868 111900 4924
rect 111900 4868 111956 4924
rect 111956 4868 111960 4924
rect 111896 4864 111960 4868
rect 111976 4924 112040 4928
rect 111976 4868 111980 4924
rect 111980 4868 112036 4924
rect 112036 4868 112040 4924
rect 111976 4864 112040 4868
rect 142456 4924 142520 4928
rect 142456 4868 142460 4924
rect 142460 4868 142516 4924
rect 142516 4868 142520 4924
rect 142456 4864 142520 4868
rect 142536 4924 142600 4928
rect 142536 4868 142540 4924
rect 142540 4868 142596 4924
rect 142596 4868 142600 4924
rect 142536 4864 142600 4868
rect 142616 4924 142680 4928
rect 142616 4868 142620 4924
rect 142620 4868 142676 4924
rect 142676 4868 142680 4924
rect 142616 4864 142680 4868
rect 142696 4924 142760 4928
rect 142696 4868 142700 4924
rect 142700 4868 142756 4924
rect 142756 4868 142760 4924
rect 142696 4864 142760 4868
rect 173176 4924 173240 4928
rect 173176 4868 173180 4924
rect 173180 4868 173236 4924
rect 173236 4868 173240 4924
rect 173176 4864 173240 4868
rect 173256 4924 173320 4928
rect 173256 4868 173260 4924
rect 173260 4868 173316 4924
rect 173316 4868 173320 4924
rect 173256 4864 173320 4868
rect 173336 4924 173400 4928
rect 173336 4868 173340 4924
rect 173340 4868 173396 4924
rect 173396 4868 173400 4924
rect 173336 4864 173400 4868
rect 173416 4924 173480 4928
rect 173416 4868 173420 4924
rect 173420 4868 173476 4924
rect 173476 4868 173480 4924
rect 173416 4864 173480 4868
rect 80652 4660 80716 4724
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 34936 4380 35000 4384
rect 34936 4324 34940 4380
rect 34940 4324 34996 4380
rect 34996 4324 35000 4380
rect 34936 4320 35000 4324
rect 35016 4380 35080 4384
rect 35016 4324 35020 4380
rect 35020 4324 35076 4380
rect 35076 4324 35080 4380
rect 35016 4320 35080 4324
rect 35096 4380 35160 4384
rect 35096 4324 35100 4380
rect 35100 4324 35156 4380
rect 35156 4324 35160 4380
rect 35096 4320 35160 4324
rect 35176 4380 35240 4384
rect 35176 4324 35180 4380
rect 35180 4324 35236 4380
rect 35236 4324 35240 4380
rect 35176 4320 35240 4324
rect 65656 4380 65720 4384
rect 65656 4324 65660 4380
rect 65660 4324 65716 4380
rect 65716 4324 65720 4380
rect 65656 4320 65720 4324
rect 65736 4380 65800 4384
rect 65736 4324 65740 4380
rect 65740 4324 65796 4380
rect 65796 4324 65800 4380
rect 65736 4320 65800 4324
rect 65816 4380 65880 4384
rect 65816 4324 65820 4380
rect 65820 4324 65876 4380
rect 65876 4324 65880 4380
rect 65816 4320 65880 4324
rect 65896 4380 65960 4384
rect 65896 4324 65900 4380
rect 65900 4324 65956 4380
rect 65956 4324 65960 4380
rect 65896 4320 65960 4324
rect 96376 4380 96440 4384
rect 96376 4324 96380 4380
rect 96380 4324 96436 4380
rect 96436 4324 96440 4380
rect 96376 4320 96440 4324
rect 96456 4380 96520 4384
rect 96456 4324 96460 4380
rect 96460 4324 96516 4380
rect 96516 4324 96520 4380
rect 96456 4320 96520 4324
rect 96536 4380 96600 4384
rect 96536 4324 96540 4380
rect 96540 4324 96596 4380
rect 96596 4324 96600 4380
rect 96536 4320 96600 4324
rect 96616 4380 96680 4384
rect 96616 4324 96620 4380
rect 96620 4324 96676 4380
rect 96676 4324 96680 4380
rect 96616 4320 96680 4324
rect 127096 4380 127160 4384
rect 127096 4324 127100 4380
rect 127100 4324 127156 4380
rect 127156 4324 127160 4380
rect 127096 4320 127160 4324
rect 127176 4380 127240 4384
rect 127176 4324 127180 4380
rect 127180 4324 127236 4380
rect 127236 4324 127240 4380
rect 127176 4320 127240 4324
rect 127256 4380 127320 4384
rect 127256 4324 127260 4380
rect 127260 4324 127316 4380
rect 127316 4324 127320 4380
rect 127256 4320 127320 4324
rect 127336 4380 127400 4384
rect 127336 4324 127340 4380
rect 127340 4324 127396 4380
rect 127396 4324 127400 4380
rect 127336 4320 127400 4324
rect 157816 4380 157880 4384
rect 157816 4324 157820 4380
rect 157820 4324 157876 4380
rect 157876 4324 157880 4380
rect 157816 4320 157880 4324
rect 157896 4380 157960 4384
rect 157896 4324 157900 4380
rect 157900 4324 157956 4380
rect 157956 4324 157960 4380
rect 157896 4320 157960 4324
rect 157976 4380 158040 4384
rect 157976 4324 157980 4380
rect 157980 4324 158036 4380
rect 158036 4324 158040 4380
rect 157976 4320 158040 4324
rect 158056 4380 158120 4384
rect 158056 4324 158060 4380
rect 158060 4324 158116 4380
rect 158116 4324 158120 4380
rect 158056 4320 158120 4324
rect 86540 4252 86604 4316
rect 86724 4040 86788 4044
rect 86724 3984 86774 4040
rect 86774 3984 86788 4040
rect 86724 3980 86788 3984
rect 19576 3836 19640 3840
rect 19576 3780 19580 3836
rect 19580 3780 19636 3836
rect 19636 3780 19640 3836
rect 19576 3776 19640 3780
rect 19656 3836 19720 3840
rect 19656 3780 19660 3836
rect 19660 3780 19716 3836
rect 19716 3780 19720 3836
rect 19656 3776 19720 3780
rect 19736 3836 19800 3840
rect 19736 3780 19740 3836
rect 19740 3780 19796 3836
rect 19796 3780 19800 3836
rect 19736 3776 19800 3780
rect 19816 3836 19880 3840
rect 19816 3780 19820 3836
rect 19820 3780 19876 3836
rect 19876 3780 19880 3836
rect 19816 3776 19880 3780
rect 50296 3836 50360 3840
rect 50296 3780 50300 3836
rect 50300 3780 50356 3836
rect 50356 3780 50360 3836
rect 50296 3776 50360 3780
rect 50376 3836 50440 3840
rect 50376 3780 50380 3836
rect 50380 3780 50436 3836
rect 50436 3780 50440 3836
rect 50376 3776 50440 3780
rect 50456 3836 50520 3840
rect 50456 3780 50460 3836
rect 50460 3780 50516 3836
rect 50516 3780 50520 3836
rect 50456 3776 50520 3780
rect 50536 3836 50600 3840
rect 50536 3780 50540 3836
rect 50540 3780 50596 3836
rect 50596 3780 50600 3836
rect 50536 3776 50600 3780
rect 81016 3836 81080 3840
rect 81016 3780 81020 3836
rect 81020 3780 81076 3836
rect 81076 3780 81080 3836
rect 81016 3776 81080 3780
rect 81096 3836 81160 3840
rect 81096 3780 81100 3836
rect 81100 3780 81156 3836
rect 81156 3780 81160 3836
rect 81096 3776 81160 3780
rect 81176 3836 81240 3840
rect 81176 3780 81180 3836
rect 81180 3780 81236 3836
rect 81236 3780 81240 3836
rect 81176 3776 81240 3780
rect 81256 3836 81320 3840
rect 81256 3780 81260 3836
rect 81260 3780 81316 3836
rect 81316 3780 81320 3836
rect 81256 3776 81320 3780
rect 111736 3836 111800 3840
rect 111736 3780 111740 3836
rect 111740 3780 111796 3836
rect 111796 3780 111800 3836
rect 111736 3776 111800 3780
rect 111816 3836 111880 3840
rect 111816 3780 111820 3836
rect 111820 3780 111876 3836
rect 111876 3780 111880 3836
rect 111816 3776 111880 3780
rect 111896 3836 111960 3840
rect 111896 3780 111900 3836
rect 111900 3780 111956 3836
rect 111956 3780 111960 3836
rect 111896 3776 111960 3780
rect 111976 3836 112040 3840
rect 111976 3780 111980 3836
rect 111980 3780 112036 3836
rect 112036 3780 112040 3836
rect 111976 3776 112040 3780
rect 142456 3836 142520 3840
rect 142456 3780 142460 3836
rect 142460 3780 142516 3836
rect 142516 3780 142520 3836
rect 142456 3776 142520 3780
rect 142536 3836 142600 3840
rect 142536 3780 142540 3836
rect 142540 3780 142596 3836
rect 142596 3780 142600 3836
rect 142536 3776 142600 3780
rect 142616 3836 142680 3840
rect 142616 3780 142620 3836
rect 142620 3780 142676 3836
rect 142676 3780 142680 3836
rect 142616 3776 142680 3780
rect 142696 3836 142760 3840
rect 142696 3780 142700 3836
rect 142700 3780 142756 3836
rect 142756 3780 142760 3836
rect 142696 3776 142760 3780
rect 173176 3836 173240 3840
rect 173176 3780 173180 3836
rect 173180 3780 173236 3836
rect 173236 3780 173240 3836
rect 173176 3776 173240 3780
rect 173256 3836 173320 3840
rect 173256 3780 173260 3836
rect 173260 3780 173316 3836
rect 173316 3780 173320 3836
rect 173256 3776 173320 3780
rect 173336 3836 173400 3840
rect 173336 3780 173340 3836
rect 173340 3780 173396 3836
rect 173396 3780 173400 3836
rect 173336 3776 173400 3780
rect 173416 3836 173480 3840
rect 173416 3780 173420 3836
rect 173420 3780 173476 3836
rect 173476 3780 173480 3836
rect 173416 3776 173480 3780
rect 88380 3708 88444 3772
rect 88748 3572 88812 3636
rect 89668 3572 89732 3636
rect 89852 3572 89916 3636
rect 86172 3436 86236 3500
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 34936 3292 35000 3296
rect 34936 3236 34940 3292
rect 34940 3236 34996 3292
rect 34996 3236 35000 3292
rect 34936 3232 35000 3236
rect 35016 3292 35080 3296
rect 35016 3236 35020 3292
rect 35020 3236 35076 3292
rect 35076 3236 35080 3292
rect 35016 3232 35080 3236
rect 35096 3292 35160 3296
rect 35096 3236 35100 3292
rect 35100 3236 35156 3292
rect 35156 3236 35160 3292
rect 35096 3232 35160 3236
rect 35176 3292 35240 3296
rect 35176 3236 35180 3292
rect 35180 3236 35236 3292
rect 35236 3236 35240 3292
rect 35176 3232 35240 3236
rect 65656 3292 65720 3296
rect 65656 3236 65660 3292
rect 65660 3236 65716 3292
rect 65716 3236 65720 3292
rect 65656 3232 65720 3236
rect 65736 3292 65800 3296
rect 65736 3236 65740 3292
rect 65740 3236 65796 3292
rect 65796 3236 65800 3292
rect 65736 3232 65800 3236
rect 65816 3292 65880 3296
rect 65816 3236 65820 3292
rect 65820 3236 65876 3292
rect 65876 3236 65880 3292
rect 65816 3232 65880 3236
rect 65896 3292 65960 3296
rect 65896 3236 65900 3292
rect 65900 3236 65956 3292
rect 65956 3236 65960 3292
rect 65896 3232 65960 3236
rect 96376 3292 96440 3296
rect 96376 3236 96380 3292
rect 96380 3236 96436 3292
rect 96436 3236 96440 3292
rect 96376 3232 96440 3236
rect 96456 3292 96520 3296
rect 96456 3236 96460 3292
rect 96460 3236 96516 3292
rect 96516 3236 96520 3292
rect 96456 3232 96520 3236
rect 96536 3292 96600 3296
rect 96536 3236 96540 3292
rect 96540 3236 96596 3292
rect 96596 3236 96600 3292
rect 96536 3232 96600 3236
rect 96616 3292 96680 3296
rect 96616 3236 96620 3292
rect 96620 3236 96676 3292
rect 96676 3236 96680 3292
rect 96616 3232 96680 3236
rect 127096 3292 127160 3296
rect 127096 3236 127100 3292
rect 127100 3236 127156 3292
rect 127156 3236 127160 3292
rect 127096 3232 127160 3236
rect 127176 3292 127240 3296
rect 127176 3236 127180 3292
rect 127180 3236 127236 3292
rect 127236 3236 127240 3292
rect 127176 3232 127240 3236
rect 127256 3292 127320 3296
rect 127256 3236 127260 3292
rect 127260 3236 127316 3292
rect 127316 3236 127320 3292
rect 127256 3232 127320 3236
rect 127336 3292 127400 3296
rect 127336 3236 127340 3292
rect 127340 3236 127396 3292
rect 127396 3236 127400 3292
rect 127336 3232 127400 3236
rect 157816 3292 157880 3296
rect 157816 3236 157820 3292
rect 157820 3236 157876 3292
rect 157876 3236 157880 3292
rect 157816 3232 157880 3236
rect 157896 3292 157960 3296
rect 157896 3236 157900 3292
rect 157900 3236 157956 3292
rect 157956 3236 157960 3292
rect 157896 3232 157960 3236
rect 157976 3292 158040 3296
rect 157976 3236 157980 3292
rect 157980 3236 158036 3292
rect 158036 3236 158040 3292
rect 157976 3232 158040 3236
rect 158056 3292 158120 3296
rect 158056 3236 158060 3292
rect 158060 3236 158116 3292
rect 158116 3236 158120 3292
rect 158056 3232 158120 3236
rect 2636 3028 2700 3092
rect 102180 3088 102244 3092
rect 102180 3032 102194 3088
rect 102194 3032 102244 3088
rect 102180 3028 102244 3032
rect 80652 2756 80716 2820
rect 19576 2748 19640 2752
rect 19576 2692 19580 2748
rect 19580 2692 19636 2748
rect 19636 2692 19640 2748
rect 19576 2688 19640 2692
rect 19656 2748 19720 2752
rect 19656 2692 19660 2748
rect 19660 2692 19716 2748
rect 19716 2692 19720 2748
rect 19656 2688 19720 2692
rect 19736 2748 19800 2752
rect 19736 2692 19740 2748
rect 19740 2692 19796 2748
rect 19796 2692 19800 2748
rect 19736 2688 19800 2692
rect 19816 2748 19880 2752
rect 19816 2692 19820 2748
rect 19820 2692 19876 2748
rect 19876 2692 19880 2748
rect 19816 2688 19880 2692
rect 50296 2748 50360 2752
rect 50296 2692 50300 2748
rect 50300 2692 50356 2748
rect 50356 2692 50360 2748
rect 50296 2688 50360 2692
rect 50376 2748 50440 2752
rect 50376 2692 50380 2748
rect 50380 2692 50436 2748
rect 50436 2692 50440 2748
rect 50376 2688 50440 2692
rect 50456 2748 50520 2752
rect 50456 2692 50460 2748
rect 50460 2692 50516 2748
rect 50516 2692 50520 2748
rect 50456 2688 50520 2692
rect 50536 2748 50600 2752
rect 50536 2692 50540 2748
rect 50540 2692 50596 2748
rect 50596 2692 50600 2748
rect 50536 2688 50600 2692
rect 86172 2756 86236 2820
rect 86540 2756 86604 2820
rect 81016 2748 81080 2752
rect 81016 2692 81020 2748
rect 81020 2692 81076 2748
rect 81076 2692 81080 2748
rect 81016 2688 81080 2692
rect 81096 2748 81160 2752
rect 81096 2692 81100 2748
rect 81100 2692 81156 2748
rect 81156 2692 81160 2748
rect 81096 2688 81160 2692
rect 81176 2748 81240 2752
rect 81176 2692 81180 2748
rect 81180 2692 81236 2748
rect 81236 2692 81240 2748
rect 81176 2688 81240 2692
rect 81256 2748 81320 2752
rect 81256 2692 81260 2748
rect 81260 2692 81316 2748
rect 81316 2692 81320 2748
rect 81256 2688 81320 2692
rect 111736 2748 111800 2752
rect 111736 2692 111740 2748
rect 111740 2692 111796 2748
rect 111796 2692 111800 2748
rect 111736 2688 111800 2692
rect 111816 2748 111880 2752
rect 111816 2692 111820 2748
rect 111820 2692 111876 2748
rect 111876 2692 111880 2748
rect 111816 2688 111880 2692
rect 111896 2748 111960 2752
rect 111896 2692 111900 2748
rect 111900 2692 111956 2748
rect 111956 2692 111960 2748
rect 111896 2688 111960 2692
rect 111976 2748 112040 2752
rect 111976 2692 111980 2748
rect 111980 2692 112036 2748
rect 112036 2692 112040 2748
rect 111976 2688 112040 2692
rect 142456 2748 142520 2752
rect 142456 2692 142460 2748
rect 142460 2692 142516 2748
rect 142516 2692 142520 2748
rect 142456 2688 142520 2692
rect 142536 2748 142600 2752
rect 142536 2692 142540 2748
rect 142540 2692 142596 2748
rect 142596 2692 142600 2748
rect 142536 2688 142600 2692
rect 142616 2748 142680 2752
rect 142616 2692 142620 2748
rect 142620 2692 142676 2748
rect 142676 2692 142680 2748
rect 142616 2688 142680 2692
rect 142696 2748 142760 2752
rect 142696 2692 142700 2748
rect 142700 2692 142756 2748
rect 142756 2692 142760 2748
rect 142696 2688 142760 2692
rect 173176 2748 173240 2752
rect 173176 2692 173180 2748
rect 173180 2692 173236 2748
rect 173236 2692 173240 2748
rect 173176 2688 173240 2692
rect 173256 2748 173320 2752
rect 173256 2692 173260 2748
rect 173260 2692 173316 2748
rect 173316 2692 173320 2748
rect 173256 2688 173320 2692
rect 173336 2748 173400 2752
rect 173336 2692 173340 2748
rect 173340 2692 173396 2748
rect 173396 2692 173400 2748
rect 173336 2688 173400 2692
rect 173416 2748 173480 2752
rect 173416 2692 173420 2748
rect 173420 2692 173476 2748
rect 173476 2692 173480 2748
rect 173416 2688 173480 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 34936 2204 35000 2208
rect 34936 2148 34940 2204
rect 34940 2148 34996 2204
rect 34996 2148 35000 2204
rect 34936 2144 35000 2148
rect 35016 2204 35080 2208
rect 35016 2148 35020 2204
rect 35020 2148 35076 2204
rect 35076 2148 35080 2204
rect 35016 2144 35080 2148
rect 35096 2204 35160 2208
rect 35096 2148 35100 2204
rect 35100 2148 35156 2204
rect 35156 2148 35160 2204
rect 35096 2144 35160 2148
rect 35176 2204 35240 2208
rect 35176 2148 35180 2204
rect 35180 2148 35236 2204
rect 35236 2148 35240 2204
rect 35176 2144 35240 2148
rect 65656 2204 65720 2208
rect 65656 2148 65660 2204
rect 65660 2148 65716 2204
rect 65716 2148 65720 2204
rect 65656 2144 65720 2148
rect 65736 2204 65800 2208
rect 65736 2148 65740 2204
rect 65740 2148 65796 2204
rect 65796 2148 65800 2204
rect 65736 2144 65800 2148
rect 65816 2204 65880 2208
rect 65816 2148 65820 2204
rect 65820 2148 65876 2204
rect 65876 2148 65880 2204
rect 65816 2144 65880 2148
rect 65896 2204 65960 2208
rect 65896 2148 65900 2204
rect 65900 2148 65956 2204
rect 65956 2148 65960 2204
rect 65896 2144 65960 2148
rect 96376 2204 96440 2208
rect 96376 2148 96380 2204
rect 96380 2148 96436 2204
rect 96436 2148 96440 2204
rect 96376 2144 96440 2148
rect 96456 2204 96520 2208
rect 96456 2148 96460 2204
rect 96460 2148 96516 2204
rect 96516 2148 96520 2204
rect 96456 2144 96520 2148
rect 96536 2204 96600 2208
rect 96536 2148 96540 2204
rect 96540 2148 96596 2204
rect 96596 2148 96600 2204
rect 96536 2144 96600 2148
rect 96616 2204 96680 2208
rect 96616 2148 96620 2204
rect 96620 2148 96676 2204
rect 96676 2148 96680 2204
rect 96616 2144 96680 2148
rect 127096 2204 127160 2208
rect 127096 2148 127100 2204
rect 127100 2148 127156 2204
rect 127156 2148 127160 2204
rect 127096 2144 127160 2148
rect 127176 2204 127240 2208
rect 127176 2148 127180 2204
rect 127180 2148 127236 2204
rect 127236 2148 127240 2204
rect 127176 2144 127240 2148
rect 127256 2204 127320 2208
rect 127256 2148 127260 2204
rect 127260 2148 127316 2204
rect 127316 2148 127320 2204
rect 127256 2144 127320 2148
rect 127336 2204 127400 2208
rect 127336 2148 127340 2204
rect 127340 2148 127396 2204
rect 127396 2148 127400 2204
rect 127336 2144 127400 2148
rect 157816 2204 157880 2208
rect 157816 2148 157820 2204
rect 157820 2148 157876 2204
rect 157876 2148 157880 2204
rect 157816 2144 157880 2148
rect 157896 2204 157960 2208
rect 157896 2148 157900 2204
rect 157900 2148 157956 2204
rect 157956 2148 157960 2204
rect 157896 2144 157960 2148
rect 157976 2204 158040 2208
rect 157976 2148 157980 2204
rect 157980 2148 158036 2204
rect 158036 2148 158040 2204
rect 157976 2144 158040 2148
rect 158056 2204 158120 2208
rect 158056 2148 158060 2204
rect 158060 2148 158116 2204
rect 158116 2148 158120 2204
rect 158056 2144 158120 2148
rect 86724 2000 86788 2004
rect 86724 1944 86774 2000
rect 86774 1944 86788 2000
rect 86724 1940 86788 1944
<< metal4 >>
rect 4208 117536 4528 117552
rect 4208 117472 4216 117536
rect 4280 117472 4296 117536
rect 4360 117472 4376 117536
rect 4440 117472 4456 117536
rect 4520 117472 4528 117536
rect 4208 116448 4528 117472
rect 4208 116384 4216 116448
rect 4280 116384 4296 116448
rect 4360 116384 4376 116448
rect 4440 116384 4456 116448
rect 4520 116384 4528 116448
rect 4208 115360 4528 116384
rect 4208 115296 4216 115360
rect 4280 115296 4296 115360
rect 4360 115296 4376 115360
rect 4440 115296 4456 115360
rect 4520 115296 4528 115360
rect 4208 114272 4528 115296
rect 4208 114208 4216 114272
rect 4280 114208 4296 114272
rect 4360 114208 4376 114272
rect 4440 114208 4456 114272
rect 4520 114208 4528 114272
rect 4208 113184 4528 114208
rect 4208 113120 4216 113184
rect 4280 113120 4296 113184
rect 4360 113120 4376 113184
rect 4440 113120 4456 113184
rect 4520 113120 4528 113184
rect 4208 112096 4528 113120
rect 4208 112032 4216 112096
rect 4280 112032 4296 112096
rect 4360 112032 4376 112096
rect 4440 112032 4456 112096
rect 4520 112032 4528 112096
rect 4208 111008 4528 112032
rect 4208 110944 4216 111008
rect 4280 110944 4296 111008
rect 4360 110944 4376 111008
rect 4440 110944 4456 111008
rect 4520 110944 4528 111008
rect 4208 109920 4528 110944
rect 4208 109856 4216 109920
rect 4280 109856 4296 109920
rect 4360 109856 4376 109920
rect 4440 109856 4456 109920
rect 4520 109856 4528 109920
rect 4208 108832 4528 109856
rect 4208 108768 4216 108832
rect 4280 108768 4296 108832
rect 4360 108768 4376 108832
rect 4440 108768 4456 108832
rect 4520 108768 4528 108832
rect 4208 107744 4528 108768
rect 4208 107680 4216 107744
rect 4280 107680 4296 107744
rect 4360 107680 4376 107744
rect 4440 107680 4456 107744
rect 4520 107680 4528 107744
rect 4208 106656 4528 107680
rect 4208 106592 4216 106656
rect 4280 106592 4296 106656
rect 4360 106592 4376 106656
rect 4440 106592 4456 106656
rect 4520 106592 4528 106656
rect 4208 105568 4528 106592
rect 4208 105504 4216 105568
rect 4280 105504 4296 105568
rect 4360 105504 4376 105568
rect 4440 105504 4456 105568
rect 4520 105504 4528 105568
rect 4208 104480 4528 105504
rect 4208 104416 4216 104480
rect 4280 104416 4296 104480
rect 4360 104416 4376 104480
rect 4440 104416 4456 104480
rect 4520 104416 4528 104480
rect 4208 103392 4528 104416
rect 4208 103328 4216 103392
rect 4280 103328 4296 103392
rect 4360 103328 4376 103392
rect 4440 103328 4456 103392
rect 4520 103328 4528 103392
rect 4208 102304 4528 103328
rect 4208 102240 4216 102304
rect 4280 102240 4296 102304
rect 4360 102240 4376 102304
rect 4440 102240 4456 102304
rect 4520 102240 4528 102304
rect 4208 101216 4528 102240
rect 4208 101152 4216 101216
rect 4280 101152 4296 101216
rect 4360 101152 4376 101216
rect 4440 101152 4456 101216
rect 4520 101152 4528 101216
rect 4208 100128 4528 101152
rect 4208 100064 4216 100128
rect 4280 100064 4296 100128
rect 4360 100064 4376 100128
rect 4440 100064 4456 100128
rect 4520 100064 4528 100128
rect 4208 99040 4528 100064
rect 4208 98976 4216 99040
rect 4280 98976 4296 99040
rect 4360 98976 4376 99040
rect 4440 98976 4456 99040
rect 4520 98976 4528 99040
rect 4208 97952 4528 98976
rect 4208 97888 4216 97952
rect 4280 97888 4296 97952
rect 4360 97888 4376 97952
rect 4440 97888 4456 97952
rect 4520 97888 4528 97952
rect 4208 96864 4528 97888
rect 4208 96800 4216 96864
rect 4280 96800 4296 96864
rect 4360 96800 4376 96864
rect 4440 96800 4456 96864
rect 4520 96800 4528 96864
rect 4208 95776 4528 96800
rect 4208 95712 4216 95776
rect 4280 95712 4296 95776
rect 4360 95712 4376 95776
rect 4440 95712 4456 95776
rect 4520 95712 4528 95776
rect 4208 94688 4528 95712
rect 4208 94624 4216 94688
rect 4280 94624 4296 94688
rect 4360 94624 4376 94688
rect 4440 94624 4456 94688
rect 4520 94624 4528 94688
rect 4208 93600 4528 94624
rect 4208 93536 4216 93600
rect 4280 93536 4296 93600
rect 4360 93536 4376 93600
rect 4440 93536 4456 93600
rect 4520 93536 4528 93600
rect 4208 92512 4528 93536
rect 4208 92448 4216 92512
rect 4280 92448 4296 92512
rect 4360 92448 4376 92512
rect 4440 92448 4456 92512
rect 4520 92448 4528 92512
rect 4208 91424 4528 92448
rect 4208 91360 4216 91424
rect 4280 91360 4296 91424
rect 4360 91360 4376 91424
rect 4440 91360 4456 91424
rect 4520 91360 4528 91424
rect 4208 90336 4528 91360
rect 4208 90272 4216 90336
rect 4280 90272 4296 90336
rect 4360 90272 4376 90336
rect 4440 90272 4456 90336
rect 4520 90272 4528 90336
rect 4208 89248 4528 90272
rect 4208 89184 4216 89248
rect 4280 89184 4296 89248
rect 4360 89184 4376 89248
rect 4440 89184 4456 89248
rect 4520 89184 4528 89248
rect 4208 88160 4528 89184
rect 4208 88096 4216 88160
rect 4280 88096 4296 88160
rect 4360 88096 4376 88160
rect 4440 88096 4456 88160
rect 4520 88096 4528 88160
rect 4208 87072 4528 88096
rect 4208 87008 4216 87072
rect 4280 87008 4296 87072
rect 4360 87008 4376 87072
rect 4440 87008 4456 87072
rect 4520 87008 4528 87072
rect 4208 85984 4528 87008
rect 4208 85920 4216 85984
rect 4280 85920 4296 85984
rect 4360 85920 4376 85984
rect 4440 85920 4456 85984
rect 4520 85920 4528 85984
rect 4208 84896 4528 85920
rect 4208 84832 4216 84896
rect 4280 84832 4296 84896
rect 4360 84832 4376 84896
rect 4440 84832 4456 84896
rect 4520 84832 4528 84896
rect 4208 83808 4528 84832
rect 4208 83744 4216 83808
rect 4280 83744 4296 83808
rect 4360 83744 4376 83808
rect 4440 83744 4456 83808
rect 4520 83744 4528 83808
rect 4208 82720 4528 83744
rect 4208 82656 4216 82720
rect 4280 82656 4296 82720
rect 4360 82656 4376 82720
rect 4440 82656 4456 82720
rect 4520 82656 4528 82720
rect 4208 81632 4528 82656
rect 4208 81568 4216 81632
rect 4280 81568 4296 81632
rect 4360 81568 4376 81632
rect 4440 81568 4456 81632
rect 4520 81568 4528 81632
rect 4208 80544 4528 81568
rect 4208 80480 4216 80544
rect 4280 80480 4296 80544
rect 4360 80480 4376 80544
rect 4440 80480 4456 80544
rect 4520 80480 4528 80544
rect 4208 79456 4528 80480
rect 4208 79392 4216 79456
rect 4280 79392 4296 79456
rect 4360 79392 4376 79456
rect 4440 79392 4456 79456
rect 4520 79392 4528 79456
rect 4208 78368 4528 79392
rect 4208 78304 4216 78368
rect 4280 78304 4296 78368
rect 4360 78304 4376 78368
rect 4440 78304 4456 78368
rect 4520 78304 4528 78368
rect 4208 77280 4528 78304
rect 4208 77216 4216 77280
rect 4280 77216 4296 77280
rect 4360 77216 4376 77280
rect 4440 77216 4456 77280
rect 4520 77216 4528 77280
rect 4208 76192 4528 77216
rect 4208 76128 4216 76192
rect 4280 76128 4296 76192
rect 4360 76128 4376 76192
rect 4440 76128 4456 76192
rect 4520 76128 4528 76192
rect 4208 75104 4528 76128
rect 4208 75040 4216 75104
rect 4280 75040 4296 75104
rect 4360 75040 4376 75104
rect 4440 75040 4456 75104
rect 4520 75040 4528 75104
rect 4208 74016 4528 75040
rect 4208 73952 4216 74016
rect 4280 73952 4296 74016
rect 4360 73952 4376 74016
rect 4440 73952 4456 74016
rect 4520 73952 4528 74016
rect 4208 72928 4528 73952
rect 4208 72864 4216 72928
rect 4280 72864 4296 72928
rect 4360 72864 4376 72928
rect 4440 72864 4456 72928
rect 4520 72864 4528 72928
rect 4208 71840 4528 72864
rect 4208 71776 4216 71840
rect 4280 71776 4296 71840
rect 4360 71776 4376 71840
rect 4440 71776 4456 71840
rect 4520 71776 4528 71840
rect 4208 70752 4528 71776
rect 4208 70688 4216 70752
rect 4280 70688 4296 70752
rect 4360 70688 4376 70752
rect 4440 70688 4456 70752
rect 4520 70688 4528 70752
rect 4208 69664 4528 70688
rect 4208 69600 4216 69664
rect 4280 69600 4296 69664
rect 4360 69600 4376 69664
rect 4440 69600 4456 69664
rect 4520 69600 4528 69664
rect 4208 68576 4528 69600
rect 4208 68512 4216 68576
rect 4280 68512 4296 68576
rect 4360 68512 4376 68576
rect 4440 68512 4456 68576
rect 4520 68512 4528 68576
rect 4208 67488 4528 68512
rect 4208 67424 4216 67488
rect 4280 67424 4296 67488
rect 4360 67424 4376 67488
rect 4440 67424 4456 67488
rect 4520 67424 4528 67488
rect 4208 66400 4528 67424
rect 4208 66336 4216 66400
rect 4280 66336 4296 66400
rect 4360 66336 4376 66400
rect 4440 66336 4456 66400
rect 4520 66336 4528 66400
rect 4208 65312 4528 66336
rect 4208 65248 4216 65312
rect 4280 65248 4296 65312
rect 4360 65248 4376 65312
rect 4440 65248 4456 65312
rect 4520 65248 4528 65312
rect 4208 64224 4528 65248
rect 4208 64160 4216 64224
rect 4280 64160 4296 64224
rect 4360 64160 4376 64224
rect 4440 64160 4456 64224
rect 4520 64160 4528 64224
rect 4208 63136 4528 64160
rect 4208 63072 4216 63136
rect 4280 63072 4296 63136
rect 4360 63072 4376 63136
rect 4440 63072 4456 63136
rect 4520 63072 4528 63136
rect 4208 62048 4528 63072
rect 4208 61984 4216 62048
rect 4280 61984 4296 62048
rect 4360 61984 4376 62048
rect 4440 61984 4456 62048
rect 4520 61984 4528 62048
rect 4208 60960 4528 61984
rect 4208 60896 4216 60960
rect 4280 60896 4296 60960
rect 4360 60896 4376 60960
rect 4440 60896 4456 60960
rect 4520 60896 4528 60960
rect 4208 59872 4528 60896
rect 4208 59808 4216 59872
rect 4280 59808 4296 59872
rect 4360 59808 4376 59872
rect 4440 59808 4456 59872
rect 4520 59808 4528 59872
rect 4208 58784 4528 59808
rect 4208 58720 4216 58784
rect 4280 58720 4296 58784
rect 4360 58720 4376 58784
rect 4440 58720 4456 58784
rect 4520 58720 4528 58784
rect 4208 57696 4528 58720
rect 4208 57632 4216 57696
rect 4280 57632 4296 57696
rect 4360 57632 4376 57696
rect 4440 57632 4456 57696
rect 4520 57632 4528 57696
rect 4208 56608 4528 57632
rect 4208 56544 4216 56608
rect 4280 56544 4296 56608
rect 4360 56544 4376 56608
rect 4440 56544 4456 56608
rect 4520 56544 4528 56608
rect 4208 55520 4528 56544
rect 4208 55456 4216 55520
rect 4280 55456 4296 55520
rect 4360 55456 4376 55520
rect 4440 55456 4456 55520
rect 4520 55456 4528 55520
rect 4208 54432 4528 55456
rect 4208 54368 4216 54432
rect 4280 54368 4296 54432
rect 4360 54368 4376 54432
rect 4440 54368 4456 54432
rect 4520 54368 4528 54432
rect 4208 53344 4528 54368
rect 4208 53280 4216 53344
rect 4280 53280 4296 53344
rect 4360 53280 4376 53344
rect 4440 53280 4456 53344
rect 4520 53280 4528 53344
rect 4208 52256 4528 53280
rect 4208 52192 4216 52256
rect 4280 52192 4296 52256
rect 4360 52192 4376 52256
rect 4440 52192 4456 52256
rect 4520 52192 4528 52256
rect 4208 51168 4528 52192
rect 4208 51104 4216 51168
rect 4280 51104 4296 51168
rect 4360 51104 4376 51168
rect 4440 51104 4456 51168
rect 4520 51104 4528 51168
rect 4208 50080 4528 51104
rect 4208 50016 4216 50080
rect 4280 50016 4296 50080
rect 4360 50016 4376 50080
rect 4440 50016 4456 50080
rect 4520 50016 4528 50080
rect 4208 48992 4528 50016
rect 4208 48928 4216 48992
rect 4280 48928 4296 48992
rect 4360 48928 4376 48992
rect 4440 48928 4456 48992
rect 4520 48928 4528 48992
rect 4208 47904 4528 48928
rect 4208 47840 4216 47904
rect 4280 47840 4296 47904
rect 4360 47840 4376 47904
rect 4440 47840 4456 47904
rect 4520 47840 4528 47904
rect 4208 46816 4528 47840
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 45728 4528 46752
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 44640 4528 45664
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 43552 4528 44576
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 42464 4528 43488
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 41376 4528 42400
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 40288 4528 41312
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 39200 4528 40224
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 38112 4528 39136
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 37024 4528 38048
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 35936 4528 36960
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5472 4528 6496
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4868 2176 5188 117504
rect 5528 2176 5848 117504
rect 6188 2176 6508 117504
rect 19568 116992 19888 117552
rect 34928 117536 35248 117552
rect 19568 116928 19576 116992
rect 19640 116928 19656 116992
rect 19720 116928 19736 116992
rect 19800 116928 19816 116992
rect 19880 116928 19888 116992
rect 19568 115904 19888 116928
rect 19568 115840 19576 115904
rect 19640 115840 19656 115904
rect 19720 115840 19736 115904
rect 19800 115840 19816 115904
rect 19880 115840 19888 115904
rect 19568 114816 19888 115840
rect 19568 114752 19576 114816
rect 19640 114752 19656 114816
rect 19720 114752 19736 114816
rect 19800 114752 19816 114816
rect 19880 114752 19888 114816
rect 19568 113728 19888 114752
rect 19568 113664 19576 113728
rect 19640 113664 19656 113728
rect 19720 113664 19736 113728
rect 19800 113664 19816 113728
rect 19880 113664 19888 113728
rect 19568 112640 19888 113664
rect 19568 112576 19576 112640
rect 19640 112576 19656 112640
rect 19720 112576 19736 112640
rect 19800 112576 19816 112640
rect 19880 112576 19888 112640
rect 19568 111552 19888 112576
rect 19568 111488 19576 111552
rect 19640 111488 19656 111552
rect 19720 111488 19736 111552
rect 19800 111488 19816 111552
rect 19880 111488 19888 111552
rect 19568 110464 19888 111488
rect 19568 110400 19576 110464
rect 19640 110400 19656 110464
rect 19720 110400 19736 110464
rect 19800 110400 19816 110464
rect 19880 110400 19888 110464
rect 19568 109376 19888 110400
rect 19568 109312 19576 109376
rect 19640 109312 19656 109376
rect 19720 109312 19736 109376
rect 19800 109312 19816 109376
rect 19880 109312 19888 109376
rect 19568 108288 19888 109312
rect 19568 108224 19576 108288
rect 19640 108224 19656 108288
rect 19720 108224 19736 108288
rect 19800 108224 19816 108288
rect 19880 108224 19888 108288
rect 19568 107200 19888 108224
rect 19568 107136 19576 107200
rect 19640 107136 19656 107200
rect 19720 107136 19736 107200
rect 19800 107136 19816 107200
rect 19880 107136 19888 107200
rect 19568 106112 19888 107136
rect 19568 106048 19576 106112
rect 19640 106048 19656 106112
rect 19720 106048 19736 106112
rect 19800 106048 19816 106112
rect 19880 106048 19888 106112
rect 19568 105024 19888 106048
rect 19568 104960 19576 105024
rect 19640 104960 19656 105024
rect 19720 104960 19736 105024
rect 19800 104960 19816 105024
rect 19880 104960 19888 105024
rect 19568 103936 19888 104960
rect 19568 103872 19576 103936
rect 19640 103872 19656 103936
rect 19720 103872 19736 103936
rect 19800 103872 19816 103936
rect 19880 103872 19888 103936
rect 19568 102848 19888 103872
rect 19568 102784 19576 102848
rect 19640 102784 19656 102848
rect 19720 102784 19736 102848
rect 19800 102784 19816 102848
rect 19880 102784 19888 102848
rect 19568 101760 19888 102784
rect 19568 101696 19576 101760
rect 19640 101696 19656 101760
rect 19720 101696 19736 101760
rect 19800 101696 19816 101760
rect 19880 101696 19888 101760
rect 19568 100672 19888 101696
rect 19568 100608 19576 100672
rect 19640 100608 19656 100672
rect 19720 100608 19736 100672
rect 19800 100608 19816 100672
rect 19880 100608 19888 100672
rect 19568 99584 19888 100608
rect 19568 99520 19576 99584
rect 19640 99520 19656 99584
rect 19720 99520 19736 99584
rect 19800 99520 19816 99584
rect 19880 99520 19888 99584
rect 19568 98496 19888 99520
rect 19568 98432 19576 98496
rect 19640 98432 19656 98496
rect 19720 98432 19736 98496
rect 19800 98432 19816 98496
rect 19880 98432 19888 98496
rect 19568 97408 19888 98432
rect 19568 97344 19576 97408
rect 19640 97344 19656 97408
rect 19720 97344 19736 97408
rect 19800 97344 19816 97408
rect 19880 97344 19888 97408
rect 19568 96320 19888 97344
rect 19568 96256 19576 96320
rect 19640 96256 19656 96320
rect 19720 96256 19736 96320
rect 19800 96256 19816 96320
rect 19880 96256 19888 96320
rect 19568 95232 19888 96256
rect 19568 95168 19576 95232
rect 19640 95168 19656 95232
rect 19720 95168 19736 95232
rect 19800 95168 19816 95232
rect 19880 95168 19888 95232
rect 19568 94144 19888 95168
rect 19568 94080 19576 94144
rect 19640 94080 19656 94144
rect 19720 94080 19736 94144
rect 19800 94080 19816 94144
rect 19880 94080 19888 94144
rect 19568 93056 19888 94080
rect 19568 92992 19576 93056
rect 19640 92992 19656 93056
rect 19720 92992 19736 93056
rect 19800 92992 19816 93056
rect 19880 92992 19888 93056
rect 19568 91968 19888 92992
rect 19568 91904 19576 91968
rect 19640 91904 19656 91968
rect 19720 91904 19736 91968
rect 19800 91904 19816 91968
rect 19880 91904 19888 91968
rect 19568 90880 19888 91904
rect 19568 90816 19576 90880
rect 19640 90816 19656 90880
rect 19720 90816 19736 90880
rect 19800 90816 19816 90880
rect 19880 90816 19888 90880
rect 19568 89792 19888 90816
rect 19568 89728 19576 89792
rect 19640 89728 19656 89792
rect 19720 89728 19736 89792
rect 19800 89728 19816 89792
rect 19880 89728 19888 89792
rect 19568 88704 19888 89728
rect 19568 88640 19576 88704
rect 19640 88640 19656 88704
rect 19720 88640 19736 88704
rect 19800 88640 19816 88704
rect 19880 88640 19888 88704
rect 19568 87616 19888 88640
rect 19568 87552 19576 87616
rect 19640 87552 19656 87616
rect 19720 87552 19736 87616
rect 19800 87552 19816 87616
rect 19880 87552 19888 87616
rect 19568 86528 19888 87552
rect 19568 86464 19576 86528
rect 19640 86464 19656 86528
rect 19720 86464 19736 86528
rect 19800 86464 19816 86528
rect 19880 86464 19888 86528
rect 19568 85440 19888 86464
rect 19568 85376 19576 85440
rect 19640 85376 19656 85440
rect 19720 85376 19736 85440
rect 19800 85376 19816 85440
rect 19880 85376 19888 85440
rect 19568 84352 19888 85376
rect 19568 84288 19576 84352
rect 19640 84288 19656 84352
rect 19720 84288 19736 84352
rect 19800 84288 19816 84352
rect 19880 84288 19888 84352
rect 19568 83264 19888 84288
rect 19568 83200 19576 83264
rect 19640 83200 19656 83264
rect 19720 83200 19736 83264
rect 19800 83200 19816 83264
rect 19880 83200 19888 83264
rect 19568 82176 19888 83200
rect 19568 82112 19576 82176
rect 19640 82112 19656 82176
rect 19720 82112 19736 82176
rect 19800 82112 19816 82176
rect 19880 82112 19888 82176
rect 19568 81088 19888 82112
rect 19568 81024 19576 81088
rect 19640 81024 19656 81088
rect 19720 81024 19736 81088
rect 19800 81024 19816 81088
rect 19880 81024 19888 81088
rect 19568 80000 19888 81024
rect 19568 79936 19576 80000
rect 19640 79936 19656 80000
rect 19720 79936 19736 80000
rect 19800 79936 19816 80000
rect 19880 79936 19888 80000
rect 19568 78912 19888 79936
rect 19568 78848 19576 78912
rect 19640 78848 19656 78912
rect 19720 78848 19736 78912
rect 19800 78848 19816 78912
rect 19880 78848 19888 78912
rect 19568 77824 19888 78848
rect 19568 77760 19576 77824
rect 19640 77760 19656 77824
rect 19720 77760 19736 77824
rect 19800 77760 19816 77824
rect 19880 77760 19888 77824
rect 19568 76736 19888 77760
rect 19568 76672 19576 76736
rect 19640 76672 19656 76736
rect 19720 76672 19736 76736
rect 19800 76672 19816 76736
rect 19880 76672 19888 76736
rect 19568 75648 19888 76672
rect 19568 75584 19576 75648
rect 19640 75584 19656 75648
rect 19720 75584 19736 75648
rect 19800 75584 19816 75648
rect 19880 75584 19888 75648
rect 19568 74560 19888 75584
rect 19568 74496 19576 74560
rect 19640 74496 19656 74560
rect 19720 74496 19736 74560
rect 19800 74496 19816 74560
rect 19880 74496 19888 74560
rect 19568 73472 19888 74496
rect 19568 73408 19576 73472
rect 19640 73408 19656 73472
rect 19720 73408 19736 73472
rect 19800 73408 19816 73472
rect 19880 73408 19888 73472
rect 19568 72384 19888 73408
rect 19568 72320 19576 72384
rect 19640 72320 19656 72384
rect 19720 72320 19736 72384
rect 19800 72320 19816 72384
rect 19880 72320 19888 72384
rect 19568 71296 19888 72320
rect 19568 71232 19576 71296
rect 19640 71232 19656 71296
rect 19720 71232 19736 71296
rect 19800 71232 19816 71296
rect 19880 71232 19888 71296
rect 19568 70208 19888 71232
rect 19568 70144 19576 70208
rect 19640 70144 19656 70208
rect 19720 70144 19736 70208
rect 19800 70144 19816 70208
rect 19880 70144 19888 70208
rect 19568 69120 19888 70144
rect 19568 69056 19576 69120
rect 19640 69056 19656 69120
rect 19720 69056 19736 69120
rect 19800 69056 19816 69120
rect 19880 69056 19888 69120
rect 19568 68032 19888 69056
rect 19568 67968 19576 68032
rect 19640 67968 19656 68032
rect 19720 67968 19736 68032
rect 19800 67968 19816 68032
rect 19880 67968 19888 68032
rect 19568 66944 19888 67968
rect 19568 66880 19576 66944
rect 19640 66880 19656 66944
rect 19720 66880 19736 66944
rect 19800 66880 19816 66944
rect 19880 66880 19888 66944
rect 19568 65856 19888 66880
rect 19568 65792 19576 65856
rect 19640 65792 19656 65856
rect 19720 65792 19736 65856
rect 19800 65792 19816 65856
rect 19880 65792 19888 65856
rect 19568 64768 19888 65792
rect 19568 64704 19576 64768
rect 19640 64704 19656 64768
rect 19720 64704 19736 64768
rect 19800 64704 19816 64768
rect 19880 64704 19888 64768
rect 19568 63680 19888 64704
rect 19568 63616 19576 63680
rect 19640 63616 19656 63680
rect 19720 63616 19736 63680
rect 19800 63616 19816 63680
rect 19880 63616 19888 63680
rect 19568 62592 19888 63616
rect 19568 62528 19576 62592
rect 19640 62528 19656 62592
rect 19720 62528 19736 62592
rect 19800 62528 19816 62592
rect 19880 62528 19888 62592
rect 19568 61504 19888 62528
rect 19568 61440 19576 61504
rect 19640 61440 19656 61504
rect 19720 61440 19736 61504
rect 19800 61440 19816 61504
rect 19880 61440 19888 61504
rect 19568 60416 19888 61440
rect 19568 60352 19576 60416
rect 19640 60352 19656 60416
rect 19720 60352 19736 60416
rect 19800 60352 19816 60416
rect 19880 60352 19888 60416
rect 19568 59328 19888 60352
rect 19568 59264 19576 59328
rect 19640 59264 19656 59328
rect 19720 59264 19736 59328
rect 19800 59264 19816 59328
rect 19880 59264 19888 59328
rect 19568 58240 19888 59264
rect 19568 58176 19576 58240
rect 19640 58176 19656 58240
rect 19720 58176 19736 58240
rect 19800 58176 19816 58240
rect 19880 58176 19888 58240
rect 19568 57152 19888 58176
rect 19568 57088 19576 57152
rect 19640 57088 19656 57152
rect 19720 57088 19736 57152
rect 19800 57088 19816 57152
rect 19880 57088 19888 57152
rect 19568 56064 19888 57088
rect 19568 56000 19576 56064
rect 19640 56000 19656 56064
rect 19720 56000 19736 56064
rect 19800 56000 19816 56064
rect 19880 56000 19888 56064
rect 19568 54976 19888 56000
rect 19568 54912 19576 54976
rect 19640 54912 19656 54976
rect 19720 54912 19736 54976
rect 19800 54912 19816 54976
rect 19880 54912 19888 54976
rect 19568 53888 19888 54912
rect 19568 53824 19576 53888
rect 19640 53824 19656 53888
rect 19720 53824 19736 53888
rect 19800 53824 19816 53888
rect 19880 53824 19888 53888
rect 19568 52800 19888 53824
rect 19568 52736 19576 52800
rect 19640 52736 19656 52800
rect 19720 52736 19736 52800
rect 19800 52736 19816 52800
rect 19880 52736 19888 52800
rect 19568 51712 19888 52736
rect 19568 51648 19576 51712
rect 19640 51648 19656 51712
rect 19720 51648 19736 51712
rect 19800 51648 19816 51712
rect 19880 51648 19888 51712
rect 19568 50624 19888 51648
rect 19568 50560 19576 50624
rect 19640 50560 19656 50624
rect 19720 50560 19736 50624
rect 19800 50560 19816 50624
rect 19880 50560 19888 50624
rect 19568 49536 19888 50560
rect 19568 49472 19576 49536
rect 19640 49472 19656 49536
rect 19720 49472 19736 49536
rect 19800 49472 19816 49536
rect 19880 49472 19888 49536
rect 19568 48448 19888 49472
rect 19568 48384 19576 48448
rect 19640 48384 19656 48448
rect 19720 48384 19736 48448
rect 19800 48384 19816 48448
rect 19880 48384 19888 48448
rect 19568 47360 19888 48384
rect 19568 47296 19576 47360
rect 19640 47296 19656 47360
rect 19720 47296 19736 47360
rect 19800 47296 19816 47360
rect 19880 47296 19888 47360
rect 19568 46272 19888 47296
rect 19568 46208 19576 46272
rect 19640 46208 19656 46272
rect 19720 46208 19736 46272
rect 19800 46208 19816 46272
rect 19880 46208 19888 46272
rect 19568 45184 19888 46208
rect 19568 45120 19576 45184
rect 19640 45120 19656 45184
rect 19720 45120 19736 45184
rect 19800 45120 19816 45184
rect 19880 45120 19888 45184
rect 19568 44096 19888 45120
rect 19568 44032 19576 44096
rect 19640 44032 19656 44096
rect 19720 44032 19736 44096
rect 19800 44032 19816 44096
rect 19880 44032 19888 44096
rect 19568 43008 19888 44032
rect 19568 42944 19576 43008
rect 19640 42944 19656 43008
rect 19720 42944 19736 43008
rect 19800 42944 19816 43008
rect 19880 42944 19888 43008
rect 19568 41920 19888 42944
rect 19568 41856 19576 41920
rect 19640 41856 19656 41920
rect 19720 41856 19736 41920
rect 19800 41856 19816 41920
rect 19880 41856 19888 41920
rect 19568 40832 19888 41856
rect 19568 40768 19576 40832
rect 19640 40768 19656 40832
rect 19720 40768 19736 40832
rect 19800 40768 19816 40832
rect 19880 40768 19888 40832
rect 19568 39744 19888 40768
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 19568 38656 19888 39680
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 37568 19888 38592
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 36480 19888 37504
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 35392 19888 36416
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 34304 19888 35328
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 33216 19888 34240
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 32128 19888 33152
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 31040 19888 32064
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 29952 19888 30976
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 28864 19888 29888
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 27776 19888 28800
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 26688 19888 27712
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 25600 19888 26624
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 24512 19888 25536
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 23424 19888 24448
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 22336 19888 23360
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 21248 19888 22272
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 20160 19888 21184
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 19072 19888 20096
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 17984 19888 19008
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 16896 19888 17920
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 15808 19888 16832
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 14720 19888 15744
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 13632 19888 14656
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 12544 19888 13568
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 11456 19888 12480
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 10368 19888 11392
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 9280 19888 10304
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 8192 19888 9216
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 7104 19888 8128
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 6016 19888 7040
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 4928 19888 5952
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 3840 19888 4864
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 2752 19888 3776
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 4208 2128 4528 2144
rect 19568 2128 19888 2688
rect 20228 2176 20548 117504
rect 20888 2176 21208 117504
rect 21548 2176 21868 117504
rect 34928 117472 34936 117536
rect 35000 117472 35016 117536
rect 35080 117472 35096 117536
rect 35160 117472 35176 117536
rect 35240 117472 35248 117536
rect 34928 116448 35248 117472
rect 34928 116384 34936 116448
rect 35000 116384 35016 116448
rect 35080 116384 35096 116448
rect 35160 116384 35176 116448
rect 35240 116384 35248 116448
rect 34928 115360 35248 116384
rect 34928 115296 34936 115360
rect 35000 115296 35016 115360
rect 35080 115296 35096 115360
rect 35160 115296 35176 115360
rect 35240 115296 35248 115360
rect 34928 114272 35248 115296
rect 34928 114208 34936 114272
rect 35000 114208 35016 114272
rect 35080 114208 35096 114272
rect 35160 114208 35176 114272
rect 35240 114208 35248 114272
rect 34928 113184 35248 114208
rect 34928 113120 34936 113184
rect 35000 113120 35016 113184
rect 35080 113120 35096 113184
rect 35160 113120 35176 113184
rect 35240 113120 35248 113184
rect 34928 112096 35248 113120
rect 34928 112032 34936 112096
rect 35000 112032 35016 112096
rect 35080 112032 35096 112096
rect 35160 112032 35176 112096
rect 35240 112032 35248 112096
rect 34928 111008 35248 112032
rect 34928 110944 34936 111008
rect 35000 110944 35016 111008
rect 35080 110944 35096 111008
rect 35160 110944 35176 111008
rect 35240 110944 35248 111008
rect 34928 109920 35248 110944
rect 34928 109856 34936 109920
rect 35000 109856 35016 109920
rect 35080 109856 35096 109920
rect 35160 109856 35176 109920
rect 35240 109856 35248 109920
rect 34928 108832 35248 109856
rect 34928 108768 34936 108832
rect 35000 108768 35016 108832
rect 35080 108768 35096 108832
rect 35160 108768 35176 108832
rect 35240 108768 35248 108832
rect 34928 107744 35248 108768
rect 34928 107680 34936 107744
rect 35000 107680 35016 107744
rect 35080 107680 35096 107744
rect 35160 107680 35176 107744
rect 35240 107680 35248 107744
rect 34928 106656 35248 107680
rect 34928 106592 34936 106656
rect 35000 106592 35016 106656
rect 35080 106592 35096 106656
rect 35160 106592 35176 106656
rect 35240 106592 35248 106656
rect 34928 105568 35248 106592
rect 34928 105504 34936 105568
rect 35000 105504 35016 105568
rect 35080 105504 35096 105568
rect 35160 105504 35176 105568
rect 35240 105504 35248 105568
rect 34928 104480 35248 105504
rect 34928 104416 34936 104480
rect 35000 104416 35016 104480
rect 35080 104416 35096 104480
rect 35160 104416 35176 104480
rect 35240 104416 35248 104480
rect 34928 103392 35248 104416
rect 34928 103328 34936 103392
rect 35000 103328 35016 103392
rect 35080 103328 35096 103392
rect 35160 103328 35176 103392
rect 35240 103328 35248 103392
rect 34928 102304 35248 103328
rect 34928 102240 34936 102304
rect 35000 102240 35016 102304
rect 35080 102240 35096 102304
rect 35160 102240 35176 102304
rect 35240 102240 35248 102304
rect 34928 101216 35248 102240
rect 34928 101152 34936 101216
rect 35000 101152 35016 101216
rect 35080 101152 35096 101216
rect 35160 101152 35176 101216
rect 35240 101152 35248 101216
rect 34928 100128 35248 101152
rect 34928 100064 34936 100128
rect 35000 100064 35016 100128
rect 35080 100064 35096 100128
rect 35160 100064 35176 100128
rect 35240 100064 35248 100128
rect 34928 99040 35248 100064
rect 34928 98976 34936 99040
rect 35000 98976 35016 99040
rect 35080 98976 35096 99040
rect 35160 98976 35176 99040
rect 35240 98976 35248 99040
rect 34928 97952 35248 98976
rect 34928 97888 34936 97952
rect 35000 97888 35016 97952
rect 35080 97888 35096 97952
rect 35160 97888 35176 97952
rect 35240 97888 35248 97952
rect 34928 96864 35248 97888
rect 34928 96800 34936 96864
rect 35000 96800 35016 96864
rect 35080 96800 35096 96864
rect 35160 96800 35176 96864
rect 35240 96800 35248 96864
rect 34928 95776 35248 96800
rect 34928 95712 34936 95776
rect 35000 95712 35016 95776
rect 35080 95712 35096 95776
rect 35160 95712 35176 95776
rect 35240 95712 35248 95776
rect 34928 94688 35248 95712
rect 34928 94624 34936 94688
rect 35000 94624 35016 94688
rect 35080 94624 35096 94688
rect 35160 94624 35176 94688
rect 35240 94624 35248 94688
rect 34928 93600 35248 94624
rect 34928 93536 34936 93600
rect 35000 93536 35016 93600
rect 35080 93536 35096 93600
rect 35160 93536 35176 93600
rect 35240 93536 35248 93600
rect 34928 92512 35248 93536
rect 34928 92448 34936 92512
rect 35000 92448 35016 92512
rect 35080 92448 35096 92512
rect 35160 92448 35176 92512
rect 35240 92448 35248 92512
rect 34928 91424 35248 92448
rect 34928 91360 34936 91424
rect 35000 91360 35016 91424
rect 35080 91360 35096 91424
rect 35160 91360 35176 91424
rect 35240 91360 35248 91424
rect 34928 90336 35248 91360
rect 34928 90272 34936 90336
rect 35000 90272 35016 90336
rect 35080 90272 35096 90336
rect 35160 90272 35176 90336
rect 35240 90272 35248 90336
rect 34928 89248 35248 90272
rect 34928 89184 34936 89248
rect 35000 89184 35016 89248
rect 35080 89184 35096 89248
rect 35160 89184 35176 89248
rect 35240 89184 35248 89248
rect 34928 88160 35248 89184
rect 34928 88096 34936 88160
rect 35000 88096 35016 88160
rect 35080 88096 35096 88160
rect 35160 88096 35176 88160
rect 35240 88096 35248 88160
rect 34928 87072 35248 88096
rect 34928 87008 34936 87072
rect 35000 87008 35016 87072
rect 35080 87008 35096 87072
rect 35160 87008 35176 87072
rect 35240 87008 35248 87072
rect 34928 85984 35248 87008
rect 34928 85920 34936 85984
rect 35000 85920 35016 85984
rect 35080 85920 35096 85984
rect 35160 85920 35176 85984
rect 35240 85920 35248 85984
rect 34928 84896 35248 85920
rect 34928 84832 34936 84896
rect 35000 84832 35016 84896
rect 35080 84832 35096 84896
rect 35160 84832 35176 84896
rect 35240 84832 35248 84896
rect 34928 83808 35248 84832
rect 34928 83744 34936 83808
rect 35000 83744 35016 83808
rect 35080 83744 35096 83808
rect 35160 83744 35176 83808
rect 35240 83744 35248 83808
rect 34928 82720 35248 83744
rect 34928 82656 34936 82720
rect 35000 82656 35016 82720
rect 35080 82656 35096 82720
rect 35160 82656 35176 82720
rect 35240 82656 35248 82720
rect 34928 81632 35248 82656
rect 34928 81568 34936 81632
rect 35000 81568 35016 81632
rect 35080 81568 35096 81632
rect 35160 81568 35176 81632
rect 35240 81568 35248 81632
rect 34928 80544 35248 81568
rect 34928 80480 34936 80544
rect 35000 80480 35016 80544
rect 35080 80480 35096 80544
rect 35160 80480 35176 80544
rect 35240 80480 35248 80544
rect 34928 79456 35248 80480
rect 34928 79392 34936 79456
rect 35000 79392 35016 79456
rect 35080 79392 35096 79456
rect 35160 79392 35176 79456
rect 35240 79392 35248 79456
rect 34928 78368 35248 79392
rect 34928 78304 34936 78368
rect 35000 78304 35016 78368
rect 35080 78304 35096 78368
rect 35160 78304 35176 78368
rect 35240 78304 35248 78368
rect 34928 77280 35248 78304
rect 34928 77216 34936 77280
rect 35000 77216 35016 77280
rect 35080 77216 35096 77280
rect 35160 77216 35176 77280
rect 35240 77216 35248 77280
rect 34928 76192 35248 77216
rect 34928 76128 34936 76192
rect 35000 76128 35016 76192
rect 35080 76128 35096 76192
rect 35160 76128 35176 76192
rect 35240 76128 35248 76192
rect 34928 75104 35248 76128
rect 34928 75040 34936 75104
rect 35000 75040 35016 75104
rect 35080 75040 35096 75104
rect 35160 75040 35176 75104
rect 35240 75040 35248 75104
rect 34928 74016 35248 75040
rect 34928 73952 34936 74016
rect 35000 73952 35016 74016
rect 35080 73952 35096 74016
rect 35160 73952 35176 74016
rect 35240 73952 35248 74016
rect 34928 72928 35248 73952
rect 34928 72864 34936 72928
rect 35000 72864 35016 72928
rect 35080 72864 35096 72928
rect 35160 72864 35176 72928
rect 35240 72864 35248 72928
rect 34928 71840 35248 72864
rect 34928 71776 34936 71840
rect 35000 71776 35016 71840
rect 35080 71776 35096 71840
rect 35160 71776 35176 71840
rect 35240 71776 35248 71840
rect 34928 70752 35248 71776
rect 34928 70688 34936 70752
rect 35000 70688 35016 70752
rect 35080 70688 35096 70752
rect 35160 70688 35176 70752
rect 35240 70688 35248 70752
rect 34928 69664 35248 70688
rect 34928 69600 34936 69664
rect 35000 69600 35016 69664
rect 35080 69600 35096 69664
rect 35160 69600 35176 69664
rect 35240 69600 35248 69664
rect 34928 68576 35248 69600
rect 34928 68512 34936 68576
rect 35000 68512 35016 68576
rect 35080 68512 35096 68576
rect 35160 68512 35176 68576
rect 35240 68512 35248 68576
rect 34928 67488 35248 68512
rect 34928 67424 34936 67488
rect 35000 67424 35016 67488
rect 35080 67424 35096 67488
rect 35160 67424 35176 67488
rect 35240 67424 35248 67488
rect 34928 66400 35248 67424
rect 34928 66336 34936 66400
rect 35000 66336 35016 66400
rect 35080 66336 35096 66400
rect 35160 66336 35176 66400
rect 35240 66336 35248 66400
rect 34928 65312 35248 66336
rect 34928 65248 34936 65312
rect 35000 65248 35016 65312
rect 35080 65248 35096 65312
rect 35160 65248 35176 65312
rect 35240 65248 35248 65312
rect 34928 64224 35248 65248
rect 34928 64160 34936 64224
rect 35000 64160 35016 64224
rect 35080 64160 35096 64224
rect 35160 64160 35176 64224
rect 35240 64160 35248 64224
rect 34928 63136 35248 64160
rect 34928 63072 34936 63136
rect 35000 63072 35016 63136
rect 35080 63072 35096 63136
rect 35160 63072 35176 63136
rect 35240 63072 35248 63136
rect 34928 62048 35248 63072
rect 34928 61984 34936 62048
rect 35000 61984 35016 62048
rect 35080 61984 35096 62048
rect 35160 61984 35176 62048
rect 35240 61984 35248 62048
rect 34928 60960 35248 61984
rect 34928 60896 34936 60960
rect 35000 60896 35016 60960
rect 35080 60896 35096 60960
rect 35160 60896 35176 60960
rect 35240 60896 35248 60960
rect 34928 59872 35248 60896
rect 34928 59808 34936 59872
rect 35000 59808 35016 59872
rect 35080 59808 35096 59872
rect 35160 59808 35176 59872
rect 35240 59808 35248 59872
rect 34928 58784 35248 59808
rect 34928 58720 34936 58784
rect 35000 58720 35016 58784
rect 35080 58720 35096 58784
rect 35160 58720 35176 58784
rect 35240 58720 35248 58784
rect 34928 57696 35248 58720
rect 34928 57632 34936 57696
rect 35000 57632 35016 57696
rect 35080 57632 35096 57696
rect 35160 57632 35176 57696
rect 35240 57632 35248 57696
rect 34928 56608 35248 57632
rect 34928 56544 34936 56608
rect 35000 56544 35016 56608
rect 35080 56544 35096 56608
rect 35160 56544 35176 56608
rect 35240 56544 35248 56608
rect 34928 55520 35248 56544
rect 34928 55456 34936 55520
rect 35000 55456 35016 55520
rect 35080 55456 35096 55520
rect 35160 55456 35176 55520
rect 35240 55456 35248 55520
rect 34928 54432 35248 55456
rect 34928 54368 34936 54432
rect 35000 54368 35016 54432
rect 35080 54368 35096 54432
rect 35160 54368 35176 54432
rect 35240 54368 35248 54432
rect 34928 53344 35248 54368
rect 34928 53280 34936 53344
rect 35000 53280 35016 53344
rect 35080 53280 35096 53344
rect 35160 53280 35176 53344
rect 35240 53280 35248 53344
rect 34928 52256 35248 53280
rect 34928 52192 34936 52256
rect 35000 52192 35016 52256
rect 35080 52192 35096 52256
rect 35160 52192 35176 52256
rect 35240 52192 35248 52256
rect 34928 51168 35248 52192
rect 34928 51104 34936 51168
rect 35000 51104 35016 51168
rect 35080 51104 35096 51168
rect 35160 51104 35176 51168
rect 35240 51104 35248 51168
rect 34928 50080 35248 51104
rect 34928 50016 34936 50080
rect 35000 50016 35016 50080
rect 35080 50016 35096 50080
rect 35160 50016 35176 50080
rect 35240 50016 35248 50080
rect 34928 48992 35248 50016
rect 34928 48928 34936 48992
rect 35000 48928 35016 48992
rect 35080 48928 35096 48992
rect 35160 48928 35176 48992
rect 35240 48928 35248 48992
rect 34928 47904 35248 48928
rect 34928 47840 34936 47904
rect 35000 47840 35016 47904
rect 35080 47840 35096 47904
rect 35160 47840 35176 47904
rect 35240 47840 35248 47904
rect 34928 46816 35248 47840
rect 34928 46752 34936 46816
rect 35000 46752 35016 46816
rect 35080 46752 35096 46816
rect 35160 46752 35176 46816
rect 35240 46752 35248 46816
rect 34928 45728 35248 46752
rect 34928 45664 34936 45728
rect 35000 45664 35016 45728
rect 35080 45664 35096 45728
rect 35160 45664 35176 45728
rect 35240 45664 35248 45728
rect 34928 44640 35248 45664
rect 34928 44576 34936 44640
rect 35000 44576 35016 44640
rect 35080 44576 35096 44640
rect 35160 44576 35176 44640
rect 35240 44576 35248 44640
rect 34928 43552 35248 44576
rect 34928 43488 34936 43552
rect 35000 43488 35016 43552
rect 35080 43488 35096 43552
rect 35160 43488 35176 43552
rect 35240 43488 35248 43552
rect 34928 42464 35248 43488
rect 34928 42400 34936 42464
rect 35000 42400 35016 42464
rect 35080 42400 35096 42464
rect 35160 42400 35176 42464
rect 35240 42400 35248 42464
rect 34928 41376 35248 42400
rect 34928 41312 34936 41376
rect 35000 41312 35016 41376
rect 35080 41312 35096 41376
rect 35160 41312 35176 41376
rect 35240 41312 35248 41376
rect 34928 40288 35248 41312
rect 34928 40224 34936 40288
rect 35000 40224 35016 40288
rect 35080 40224 35096 40288
rect 35160 40224 35176 40288
rect 35240 40224 35248 40288
rect 34928 39200 35248 40224
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 38112 35248 39136
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 37024 35248 38048
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 35936 35248 36960
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 34848 35248 35872
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 33760 35248 34784
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 32672 35248 33696
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 31584 35248 32608
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 30496 35248 31520
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 29408 35248 30432
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 28320 35248 29344
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 27232 35248 28256
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 26144 35248 27168
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 25056 35248 26080
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 23968 35248 24992
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 22880 35248 23904
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 21792 35248 22816
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 20704 35248 21728
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 19616 35248 20640
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 18528 35248 19552
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 17440 35248 18464
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 16352 35248 17376
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 15264 35248 16288
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 14176 35248 15200
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 13088 35248 14112
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 12000 35248 13024
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 10912 35248 11936
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 9824 35248 10848
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 8736 35248 9760
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 7648 35248 8672
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 6560 35248 7584
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 5472 35248 6496
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 4384 35248 5408
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 3296 35248 4320
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 2208 35248 3232
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 35588 2176 35908 117504
rect 36248 2176 36568 117504
rect 36908 2176 37228 117504
rect 50288 116992 50608 117552
rect 65648 117536 65968 117552
rect 50288 116928 50296 116992
rect 50360 116928 50376 116992
rect 50440 116928 50456 116992
rect 50520 116928 50536 116992
rect 50600 116928 50608 116992
rect 50288 115904 50608 116928
rect 50288 115840 50296 115904
rect 50360 115840 50376 115904
rect 50440 115840 50456 115904
rect 50520 115840 50536 115904
rect 50600 115840 50608 115904
rect 50288 114816 50608 115840
rect 50288 114752 50296 114816
rect 50360 114752 50376 114816
rect 50440 114752 50456 114816
rect 50520 114752 50536 114816
rect 50600 114752 50608 114816
rect 50288 113728 50608 114752
rect 50288 113664 50296 113728
rect 50360 113664 50376 113728
rect 50440 113664 50456 113728
rect 50520 113664 50536 113728
rect 50600 113664 50608 113728
rect 50288 112640 50608 113664
rect 50288 112576 50296 112640
rect 50360 112576 50376 112640
rect 50440 112576 50456 112640
rect 50520 112576 50536 112640
rect 50600 112576 50608 112640
rect 50288 111552 50608 112576
rect 50288 111488 50296 111552
rect 50360 111488 50376 111552
rect 50440 111488 50456 111552
rect 50520 111488 50536 111552
rect 50600 111488 50608 111552
rect 50288 110464 50608 111488
rect 50288 110400 50296 110464
rect 50360 110400 50376 110464
rect 50440 110400 50456 110464
rect 50520 110400 50536 110464
rect 50600 110400 50608 110464
rect 50288 109376 50608 110400
rect 50288 109312 50296 109376
rect 50360 109312 50376 109376
rect 50440 109312 50456 109376
rect 50520 109312 50536 109376
rect 50600 109312 50608 109376
rect 50288 108288 50608 109312
rect 50288 108224 50296 108288
rect 50360 108224 50376 108288
rect 50440 108224 50456 108288
rect 50520 108224 50536 108288
rect 50600 108224 50608 108288
rect 50288 107200 50608 108224
rect 50288 107136 50296 107200
rect 50360 107136 50376 107200
rect 50440 107136 50456 107200
rect 50520 107136 50536 107200
rect 50600 107136 50608 107200
rect 50288 106112 50608 107136
rect 50288 106048 50296 106112
rect 50360 106048 50376 106112
rect 50440 106048 50456 106112
rect 50520 106048 50536 106112
rect 50600 106048 50608 106112
rect 50288 105024 50608 106048
rect 50288 104960 50296 105024
rect 50360 104960 50376 105024
rect 50440 104960 50456 105024
rect 50520 104960 50536 105024
rect 50600 104960 50608 105024
rect 50288 103936 50608 104960
rect 50288 103872 50296 103936
rect 50360 103872 50376 103936
rect 50440 103872 50456 103936
rect 50520 103872 50536 103936
rect 50600 103872 50608 103936
rect 50288 102848 50608 103872
rect 50288 102784 50296 102848
rect 50360 102784 50376 102848
rect 50440 102784 50456 102848
rect 50520 102784 50536 102848
rect 50600 102784 50608 102848
rect 50288 101760 50608 102784
rect 50288 101696 50296 101760
rect 50360 101696 50376 101760
rect 50440 101696 50456 101760
rect 50520 101696 50536 101760
rect 50600 101696 50608 101760
rect 50288 100672 50608 101696
rect 50288 100608 50296 100672
rect 50360 100608 50376 100672
rect 50440 100608 50456 100672
rect 50520 100608 50536 100672
rect 50600 100608 50608 100672
rect 50288 99584 50608 100608
rect 50288 99520 50296 99584
rect 50360 99520 50376 99584
rect 50440 99520 50456 99584
rect 50520 99520 50536 99584
rect 50600 99520 50608 99584
rect 50288 98496 50608 99520
rect 50288 98432 50296 98496
rect 50360 98432 50376 98496
rect 50440 98432 50456 98496
rect 50520 98432 50536 98496
rect 50600 98432 50608 98496
rect 50288 97408 50608 98432
rect 50288 97344 50296 97408
rect 50360 97344 50376 97408
rect 50440 97344 50456 97408
rect 50520 97344 50536 97408
rect 50600 97344 50608 97408
rect 50288 96320 50608 97344
rect 50288 96256 50296 96320
rect 50360 96256 50376 96320
rect 50440 96256 50456 96320
rect 50520 96256 50536 96320
rect 50600 96256 50608 96320
rect 50288 95232 50608 96256
rect 50288 95168 50296 95232
rect 50360 95168 50376 95232
rect 50440 95168 50456 95232
rect 50520 95168 50536 95232
rect 50600 95168 50608 95232
rect 50288 94144 50608 95168
rect 50288 94080 50296 94144
rect 50360 94080 50376 94144
rect 50440 94080 50456 94144
rect 50520 94080 50536 94144
rect 50600 94080 50608 94144
rect 50288 93056 50608 94080
rect 50288 92992 50296 93056
rect 50360 92992 50376 93056
rect 50440 92992 50456 93056
rect 50520 92992 50536 93056
rect 50600 92992 50608 93056
rect 50288 91968 50608 92992
rect 50288 91904 50296 91968
rect 50360 91904 50376 91968
rect 50440 91904 50456 91968
rect 50520 91904 50536 91968
rect 50600 91904 50608 91968
rect 50288 90880 50608 91904
rect 50288 90816 50296 90880
rect 50360 90816 50376 90880
rect 50440 90816 50456 90880
rect 50520 90816 50536 90880
rect 50600 90816 50608 90880
rect 50288 89792 50608 90816
rect 50288 89728 50296 89792
rect 50360 89728 50376 89792
rect 50440 89728 50456 89792
rect 50520 89728 50536 89792
rect 50600 89728 50608 89792
rect 50288 88704 50608 89728
rect 50288 88640 50296 88704
rect 50360 88640 50376 88704
rect 50440 88640 50456 88704
rect 50520 88640 50536 88704
rect 50600 88640 50608 88704
rect 50288 87616 50608 88640
rect 50288 87552 50296 87616
rect 50360 87552 50376 87616
rect 50440 87552 50456 87616
rect 50520 87552 50536 87616
rect 50600 87552 50608 87616
rect 50288 86528 50608 87552
rect 50288 86464 50296 86528
rect 50360 86464 50376 86528
rect 50440 86464 50456 86528
rect 50520 86464 50536 86528
rect 50600 86464 50608 86528
rect 50288 85440 50608 86464
rect 50288 85376 50296 85440
rect 50360 85376 50376 85440
rect 50440 85376 50456 85440
rect 50520 85376 50536 85440
rect 50600 85376 50608 85440
rect 50288 84352 50608 85376
rect 50288 84288 50296 84352
rect 50360 84288 50376 84352
rect 50440 84288 50456 84352
rect 50520 84288 50536 84352
rect 50600 84288 50608 84352
rect 50288 83264 50608 84288
rect 50288 83200 50296 83264
rect 50360 83200 50376 83264
rect 50440 83200 50456 83264
rect 50520 83200 50536 83264
rect 50600 83200 50608 83264
rect 50288 82176 50608 83200
rect 50288 82112 50296 82176
rect 50360 82112 50376 82176
rect 50440 82112 50456 82176
rect 50520 82112 50536 82176
rect 50600 82112 50608 82176
rect 50288 81088 50608 82112
rect 50288 81024 50296 81088
rect 50360 81024 50376 81088
rect 50440 81024 50456 81088
rect 50520 81024 50536 81088
rect 50600 81024 50608 81088
rect 50288 80000 50608 81024
rect 50288 79936 50296 80000
rect 50360 79936 50376 80000
rect 50440 79936 50456 80000
rect 50520 79936 50536 80000
rect 50600 79936 50608 80000
rect 50288 78912 50608 79936
rect 50288 78848 50296 78912
rect 50360 78848 50376 78912
rect 50440 78848 50456 78912
rect 50520 78848 50536 78912
rect 50600 78848 50608 78912
rect 50288 77824 50608 78848
rect 50288 77760 50296 77824
rect 50360 77760 50376 77824
rect 50440 77760 50456 77824
rect 50520 77760 50536 77824
rect 50600 77760 50608 77824
rect 50288 76736 50608 77760
rect 50288 76672 50296 76736
rect 50360 76672 50376 76736
rect 50440 76672 50456 76736
rect 50520 76672 50536 76736
rect 50600 76672 50608 76736
rect 50288 75648 50608 76672
rect 50288 75584 50296 75648
rect 50360 75584 50376 75648
rect 50440 75584 50456 75648
rect 50520 75584 50536 75648
rect 50600 75584 50608 75648
rect 50288 74560 50608 75584
rect 50288 74496 50296 74560
rect 50360 74496 50376 74560
rect 50440 74496 50456 74560
rect 50520 74496 50536 74560
rect 50600 74496 50608 74560
rect 50288 73472 50608 74496
rect 50288 73408 50296 73472
rect 50360 73408 50376 73472
rect 50440 73408 50456 73472
rect 50520 73408 50536 73472
rect 50600 73408 50608 73472
rect 50288 72384 50608 73408
rect 50288 72320 50296 72384
rect 50360 72320 50376 72384
rect 50440 72320 50456 72384
rect 50520 72320 50536 72384
rect 50600 72320 50608 72384
rect 50288 71296 50608 72320
rect 50288 71232 50296 71296
rect 50360 71232 50376 71296
rect 50440 71232 50456 71296
rect 50520 71232 50536 71296
rect 50600 71232 50608 71296
rect 50288 70208 50608 71232
rect 50288 70144 50296 70208
rect 50360 70144 50376 70208
rect 50440 70144 50456 70208
rect 50520 70144 50536 70208
rect 50600 70144 50608 70208
rect 50288 69120 50608 70144
rect 50288 69056 50296 69120
rect 50360 69056 50376 69120
rect 50440 69056 50456 69120
rect 50520 69056 50536 69120
rect 50600 69056 50608 69120
rect 50288 68032 50608 69056
rect 50288 67968 50296 68032
rect 50360 67968 50376 68032
rect 50440 67968 50456 68032
rect 50520 67968 50536 68032
rect 50600 67968 50608 68032
rect 50288 66944 50608 67968
rect 50288 66880 50296 66944
rect 50360 66880 50376 66944
rect 50440 66880 50456 66944
rect 50520 66880 50536 66944
rect 50600 66880 50608 66944
rect 50288 65856 50608 66880
rect 50288 65792 50296 65856
rect 50360 65792 50376 65856
rect 50440 65792 50456 65856
rect 50520 65792 50536 65856
rect 50600 65792 50608 65856
rect 50288 64768 50608 65792
rect 50288 64704 50296 64768
rect 50360 64704 50376 64768
rect 50440 64704 50456 64768
rect 50520 64704 50536 64768
rect 50600 64704 50608 64768
rect 50288 63680 50608 64704
rect 50288 63616 50296 63680
rect 50360 63616 50376 63680
rect 50440 63616 50456 63680
rect 50520 63616 50536 63680
rect 50600 63616 50608 63680
rect 50288 62592 50608 63616
rect 50288 62528 50296 62592
rect 50360 62528 50376 62592
rect 50440 62528 50456 62592
rect 50520 62528 50536 62592
rect 50600 62528 50608 62592
rect 50288 61504 50608 62528
rect 50288 61440 50296 61504
rect 50360 61440 50376 61504
rect 50440 61440 50456 61504
rect 50520 61440 50536 61504
rect 50600 61440 50608 61504
rect 50288 60416 50608 61440
rect 50288 60352 50296 60416
rect 50360 60352 50376 60416
rect 50440 60352 50456 60416
rect 50520 60352 50536 60416
rect 50600 60352 50608 60416
rect 50288 59328 50608 60352
rect 50288 59264 50296 59328
rect 50360 59264 50376 59328
rect 50440 59264 50456 59328
rect 50520 59264 50536 59328
rect 50600 59264 50608 59328
rect 50288 58240 50608 59264
rect 50288 58176 50296 58240
rect 50360 58176 50376 58240
rect 50440 58176 50456 58240
rect 50520 58176 50536 58240
rect 50600 58176 50608 58240
rect 50288 57152 50608 58176
rect 50288 57088 50296 57152
rect 50360 57088 50376 57152
rect 50440 57088 50456 57152
rect 50520 57088 50536 57152
rect 50600 57088 50608 57152
rect 50288 56064 50608 57088
rect 50288 56000 50296 56064
rect 50360 56000 50376 56064
rect 50440 56000 50456 56064
rect 50520 56000 50536 56064
rect 50600 56000 50608 56064
rect 50288 54976 50608 56000
rect 50288 54912 50296 54976
rect 50360 54912 50376 54976
rect 50440 54912 50456 54976
rect 50520 54912 50536 54976
rect 50600 54912 50608 54976
rect 50288 53888 50608 54912
rect 50288 53824 50296 53888
rect 50360 53824 50376 53888
rect 50440 53824 50456 53888
rect 50520 53824 50536 53888
rect 50600 53824 50608 53888
rect 50288 52800 50608 53824
rect 50288 52736 50296 52800
rect 50360 52736 50376 52800
rect 50440 52736 50456 52800
rect 50520 52736 50536 52800
rect 50600 52736 50608 52800
rect 50288 51712 50608 52736
rect 50288 51648 50296 51712
rect 50360 51648 50376 51712
rect 50440 51648 50456 51712
rect 50520 51648 50536 51712
rect 50600 51648 50608 51712
rect 50288 50624 50608 51648
rect 50288 50560 50296 50624
rect 50360 50560 50376 50624
rect 50440 50560 50456 50624
rect 50520 50560 50536 50624
rect 50600 50560 50608 50624
rect 50288 49536 50608 50560
rect 50288 49472 50296 49536
rect 50360 49472 50376 49536
rect 50440 49472 50456 49536
rect 50520 49472 50536 49536
rect 50600 49472 50608 49536
rect 50288 48448 50608 49472
rect 50288 48384 50296 48448
rect 50360 48384 50376 48448
rect 50440 48384 50456 48448
rect 50520 48384 50536 48448
rect 50600 48384 50608 48448
rect 50288 47360 50608 48384
rect 50288 47296 50296 47360
rect 50360 47296 50376 47360
rect 50440 47296 50456 47360
rect 50520 47296 50536 47360
rect 50600 47296 50608 47360
rect 50288 46272 50608 47296
rect 50288 46208 50296 46272
rect 50360 46208 50376 46272
rect 50440 46208 50456 46272
rect 50520 46208 50536 46272
rect 50600 46208 50608 46272
rect 50288 45184 50608 46208
rect 50288 45120 50296 45184
rect 50360 45120 50376 45184
rect 50440 45120 50456 45184
rect 50520 45120 50536 45184
rect 50600 45120 50608 45184
rect 50288 44096 50608 45120
rect 50288 44032 50296 44096
rect 50360 44032 50376 44096
rect 50440 44032 50456 44096
rect 50520 44032 50536 44096
rect 50600 44032 50608 44096
rect 50288 43008 50608 44032
rect 50288 42944 50296 43008
rect 50360 42944 50376 43008
rect 50440 42944 50456 43008
rect 50520 42944 50536 43008
rect 50600 42944 50608 43008
rect 50288 41920 50608 42944
rect 50288 41856 50296 41920
rect 50360 41856 50376 41920
rect 50440 41856 50456 41920
rect 50520 41856 50536 41920
rect 50600 41856 50608 41920
rect 50288 40832 50608 41856
rect 50288 40768 50296 40832
rect 50360 40768 50376 40832
rect 50440 40768 50456 40832
rect 50520 40768 50536 40832
rect 50600 40768 50608 40832
rect 50288 39744 50608 40768
rect 50288 39680 50296 39744
rect 50360 39680 50376 39744
rect 50440 39680 50456 39744
rect 50520 39680 50536 39744
rect 50600 39680 50608 39744
rect 50288 38656 50608 39680
rect 50288 38592 50296 38656
rect 50360 38592 50376 38656
rect 50440 38592 50456 38656
rect 50520 38592 50536 38656
rect 50600 38592 50608 38656
rect 50288 37568 50608 38592
rect 50288 37504 50296 37568
rect 50360 37504 50376 37568
rect 50440 37504 50456 37568
rect 50520 37504 50536 37568
rect 50600 37504 50608 37568
rect 50288 36480 50608 37504
rect 50288 36416 50296 36480
rect 50360 36416 50376 36480
rect 50440 36416 50456 36480
rect 50520 36416 50536 36480
rect 50600 36416 50608 36480
rect 50288 35392 50608 36416
rect 50288 35328 50296 35392
rect 50360 35328 50376 35392
rect 50440 35328 50456 35392
rect 50520 35328 50536 35392
rect 50600 35328 50608 35392
rect 50288 34304 50608 35328
rect 50288 34240 50296 34304
rect 50360 34240 50376 34304
rect 50440 34240 50456 34304
rect 50520 34240 50536 34304
rect 50600 34240 50608 34304
rect 50288 33216 50608 34240
rect 50288 33152 50296 33216
rect 50360 33152 50376 33216
rect 50440 33152 50456 33216
rect 50520 33152 50536 33216
rect 50600 33152 50608 33216
rect 50288 32128 50608 33152
rect 50288 32064 50296 32128
rect 50360 32064 50376 32128
rect 50440 32064 50456 32128
rect 50520 32064 50536 32128
rect 50600 32064 50608 32128
rect 50288 31040 50608 32064
rect 50288 30976 50296 31040
rect 50360 30976 50376 31040
rect 50440 30976 50456 31040
rect 50520 30976 50536 31040
rect 50600 30976 50608 31040
rect 50288 29952 50608 30976
rect 50288 29888 50296 29952
rect 50360 29888 50376 29952
rect 50440 29888 50456 29952
rect 50520 29888 50536 29952
rect 50600 29888 50608 29952
rect 50288 28864 50608 29888
rect 50288 28800 50296 28864
rect 50360 28800 50376 28864
rect 50440 28800 50456 28864
rect 50520 28800 50536 28864
rect 50600 28800 50608 28864
rect 50288 27776 50608 28800
rect 50288 27712 50296 27776
rect 50360 27712 50376 27776
rect 50440 27712 50456 27776
rect 50520 27712 50536 27776
rect 50600 27712 50608 27776
rect 50288 26688 50608 27712
rect 50288 26624 50296 26688
rect 50360 26624 50376 26688
rect 50440 26624 50456 26688
rect 50520 26624 50536 26688
rect 50600 26624 50608 26688
rect 50288 25600 50608 26624
rect 50288 25536 50296 25600
rect 50360 25536 50376 25600
rect 50440 25536 50456 25600
rect 50520 25536 50536 25600
rect 50600 25536 50608 25600
rect 50288 24512 50608 25536
rect 50288 24448 50296 24512
rect 50360 24448 50376 24512
rect 50440 24448 50456 24512
rect 50520 24448 50536 24512
rect 50600 24448 50608 24512
rect 50288 23424 50608 24448
rect 50288 23360 50296 23424
rect 50360 23360 50376 23424
rect 50440 23360 50456 23424
rect 50520 23360 50536 23424
rect 50600 23360 50608 23424
rect 50288 22336 50608 23360
rect 50288 22272 50296 22336
rect 50360 22272 50376 22336
rect 50440 22272 50456 22336
rect 50520 22272 50536 22336
rect 50600 22272 50608 22336
rect 50288 21248 50608 22272
rect 50288 21184 50296 21248
rect 50360 21184 50376 21248
rect 50440 21184 50456 21248
rect 50520 21184 50536 21248
rect 50600 21184 50608 21248
rect 50288 20160 50608 21184
rect 50288 20096 50296 20160
rect 50360 20096 50376 20160
rect 50440 20096 50456 20160
rect 50520 20096 50536 20160
rect 50600 20096 50608 20160
rect 50288 19072 50608 20096
rect 50288 19008 50296 19072
rect 50360 19008 50376 19072
rect 50440 19008 50456 19072
rect 50520 19008 50536 19072
rect 50600 19008 50608 19072
rect 50288 17984 50608 19008
rect 50288 17920 50296 17984
rect 50360 17920 50376 17984
rect 50440 17920 50456 17984
rect 50520 17920 50536 17984
rect 50600 17920 50608 17984
rect 50288 16896 50608 17920
rect 50288 16832 50296 16896
rect 50360 16832 50376 16896
rect 50440 16832 50456 16896
rect 50520 16832 50536 16896
rect 50600 16832 50608 16896
rect 50288 15808 50608 16832
rect 50288 15744 50296 15808
rect 50360 15744 50376 15808
rect 50440 15744 50456 15808
rect 50520 15744 50536 15808
rect 50600 15744 50608 15808
rect 50288 14720 50608 15744
rect 50288 14656 50296 14720
rect 50360 14656 50376 14720
rect 50440 14656 50456 14720
rect 50520 14656 50536 14720
rect 50600 14656 50608 14720
rect 50288 13632 50608 14656
rect 50288 13568 50296 13632
rect 50360 13568 50376 13632
rect 50440 13568 50456 13632
rect 50520 13568 50536 13632
rect 50600 13568 50608 13632
rect 50288 12544 50608 13568
rect 50288 12480 50296 12544
rect 50360 12480 50376 12544
rect 50440 12480 50456 12544
rect 50520 12480 50536 12544
rect 50600 12480 50608 12544
rect 50288 11456 50608 12480
rect 50288 11392 50296 11456
rect 50360 11392 50376 11456
rect 50440 11392 50456 11456
rect 50520 11392 50536 11456
rect 50600 11392 50608 11456
rect 50288 10368 50608 11392
rect 50288 10304 50296 10368
rect 50360 10304 50376 10368
rect 50440 10304 50456 10368
rect 50520 10304 50536 10368
rect 50600 10304 50608 10368
rect 50288 9280 50608 10304
rect 50288 9216 50296 9280
rect 50360 9216 50376 9280
rect 50440 9216 50456 9280
rect 50520 9216 50536 9280
rect 50600 9216 50608 9280
rect 50288 8192 50608 9216
rect 50288 8128 50296 8192
rect 50360 8128 50376 8192
rect 50440 8128 50456 8192
rect 50520 8128 50536 8192
rect 50600 8128 50608 8192
rect 50288 7104 50608 8128
rect 50288 7040 50296 7104
rect 50360 7040 50376 7104
rect 50440 7040 50456 7104
rect 50520 7040 50536 7104
rect 50600 7040 50608 7104
rect 50288 6016 50608 7040
rect 50288 5952 50296 6016
rect 50360 5952 50376 6016
rect 50440 5952 50456 6016
rect 50520 5952 50536 6016
rect 50600 5952 50608 6016
rect 50288 4928 50608 5952
rect 50288 4864 50296 4928
rect 50360 4864 50376 4928
rect 50440 4864 50456 4928
rect 50520 4864 50536 4928
rect 50600 4864 50608 4928
rect 50288 3840 50608 4864
rect 50288 3776 50296 3840
rect 50360 3776 50376 3840
rect 50440 3776 50456 3840
rect 50520 3776 50536 3840
rect 50600 3776 50608 3840
rect 50288 2752 50608 3776
rect 50288 2688 50296 2752
rect 50360 2688 50376 2752
rect 50440 2688 50456 2752
rect 50520 2688 50536 2752
rect 50600 2688 50608 2752
rect 34928 2128 35248 2144
rect 50288 2128 50608 2688
rect 50948 2176 51268 117504
rect 51608 2176 51928 117504
rect 52268 2176 52588 117504
rect 65648 117472 65656 117536
rect 65720 117472 65736 117536
rect 65800 117472 65816 117536
rect 65880 117472 65896 117536
rect 65960 117472 65968 117536
rect 65648 116448 65968 117472
rect 65648 116384 65656 116448
rect 65720 116384 65736 116448
rect 65800 116384 65816 116448
rect 65880 116384 65896 116448
rect 65960 116384 65968 116448
rect 65648 115360 65968 116384
rect 65648 115296 65656 115360
rect 65720 115296 65736 115360
rect 65800 115296 65816 115360
rect 65880 115296 65896 115360
rect 65960 115296 65968 115360
rect 65648 114272 65968 115296
rect 65648 114208 65656 114272
rect 65720 114208 65736 114272
rect 65800 114208 65816 114272
rect 65880 114208 65896 114272
rect 65960 114208 65968 114272
rect 65648 113184 65968 114208
rect 65648 113120 65656 113184
rect 65720 113120 65736 113184
rect 65800 113120 65816 113184
rect 65880 113120 65896 113184
rect 65960 113120 65968 113184
rect 65648 112096 65968 113120
rect 65648 112032 65656 112096
rect 65720 112032 65736 112096
rect 65800 112032 65816 112096
rect 65880 112032 65896 112096
rect 65960 112032 65968 112096
rect 65648 111008 65968 112032
rect 65648 110944 65656 111008
rect 65720 110944 65736 111008
rect 65800 110944 65816 111008
rect 65880 110944 65896 111008
rect 65960 110944 65968 111008
rect 65648 109920 65968 110944
rect 65648 109856 65656 109920
rect 65720 109856 65736 109920
rect 65800 109856 65816 109920
rect 65880 109856 65896 109920
rect 65960 109856 65968 109920
rect 65648 108832 65968 109856
rect 65648 108768 65656 108832
rect 65720 108768 65736 108832
rect 65800 108768 65816 108832
rect 65880 108768 65896 108832
rect 65960 108768 65968 108832
rect 65648 107744 65968 108768
rect 65648 107680 65656 107744
rect 65720 107680 65736 107744
rect 65800 107680 65816 107744
rect 65880 107680 65896 107744
rect 65960 107680 65968 107744
rect 65648 106656 65968 107680
rect 65648 106592 65656 106656
rect 65720 106592 65736 106656
rect 65800 106592 65816 106656
rect 65880 106592 65896 106656
rect 65960 106592 65968 106656
rect 65648 105568 65968 106592
rect 65648 105504 65656 105568
rect 65720 105504 65736 105568
rect 65800 105504 65816 105568
rect 65880 105504 65896 105568
rect 65960 105504 65968 105568
rect 65648 104480 65968 105504
rect 65648 104416 65656 104480
rect 65720 104416 65736 104480
rect 65800 104416 65816 104480
rect 65880 104416 65896 104480
rect 65960 104416 65968 104480
rect 65648 103392 65968 104416
rect 65648 103328 65656 103392
rect 65720 103328 65736 103392
rect 65800 103328 65816 103392
rect 65880 103328 65896 103392
rect 65960 103328 65968 103392
rect 65648 102304 65968 103328
rect 65648 102240 65656 102304
rect 65720 102240 65736 102304
rect 65800 102240 65816 102304
rect 65880 102240 65896 102304
rect 65960 102240 65968 102304
rect 65648 101216 65968 102240
rect 65648 101152 65656 101216
rect 65720 101152 65736 101216
rect 65800 101152 65816 101216
rect 65880 101152 65896 101216
rect 65960 101152 65968 101216
rect 65648 100128 65968 101152
rect 65648 100064 65656 100128
rect 65720 100064 65736 100128
rect 65800 100064 65816 100128
rect 65880 100064 65896 100128
rect 65960 100064 65968 100128
rect 65648 99040 65968 100064
rect 65648 98976 65656 99040
rect 65720 98976 65736 99040
rect 65800 98976 65816 99040
rect 65880 98976 65896 99040
rect 65960 98976 65968 99040
rect 65648 97952 65968 98976
rect 65648 97888 65656 97952
rect 65720 97888 65736 97952
rect 65800 97888 65816 97952
rect 65880 97888 65896 97952
rect 65960 97888 65968 97952
rect 65648 96864 65968 97888
rect 65648 96800 65656 96864
rect 65720 96800 65736 96864
rect 65800 96800 65816 96864
rect 65880 96800 65896 96864
rect 65960 96800 65968 96864
rect 65648 95776 65968 96800
rect 65648 95712 65656 95776
rect 65720 95712 65736 95776
rect 65800 95712 65816 95776
rect 65880 95712 65896 95776
rect 65960 95712 65968 95776
rect 65648 94688 65968 95712
rect 65648 94624 65656 94688
rect 65720 94624 65736 94688
rect 65800 94624 65816 94688
rect 65880 94624 65896 94688
rect 65960 94624 65968 94688
rect 65648 93600 65968 94624
rect 65648 93536 65656 93600
rect 65720 93536 65736 93600
rect 65800 93536 65816 93600
rect 65880 93536 65896 93600
rect 65960 93536 65968 93600
rect 65648 92512 65968 93536
rect 65648 92448 65656 92512
rect 65720 92448 65736 92512
rect 65800 92448 65816 92512
rect 65880 92448 65896 92512
rect 65960 92448 65968 92512
rect 65648 91424 65968 92448
rect 65648 91360 65656 91424
rect 65720 91360 65736 91424
rect 65800 91360 65816 91424
rect 65880 91360 65896 91424
rect 65960 91360 65968 91424
rect 65648 90336 65968 91360
rect 65648 90272 65656 90336
rect 65720 90272 65736 90336
rect 65800 90272 65816 90336
rect 65880 90272 65896 90336
rect 65960 90272 65968 90336
rect 65648 89248 65968 90272
rect 65648 89184 65656 89248
rect 65720 89184 65736 89248
rect 65800 89184 65816 89248
rect 65880 89184 65896 89248
rect 65960 89184 65968 89248
rect 65648 88160 65968 89184
rect 65648 88096 65656 88160
rect 65720 88096 65736 88160
rect 65800 88096 65816 88160
rect 65880 88096 65896 88160
rect 65960 88096 65968 88160
rect 65648 87072 65968 88096
rect 65648 87008 65656 87072
rect 65720 87008 65736 87072
rect 65800 87008 65816 87072
rect 65880 87008 65896 87072
rect 65960 87008 65968 87072
rect 65648 85984 65968 87008
rect 65648 85920 65656 85984
rect 65720 85920 65736 85984
rect 65800 85920 65816 85984
rect 65880 85920 65896 85984
rect 65960 85920 65968 85984
rect 65648 84896 65968 85920
rect 65648 84832 65656 84896
rect 65720 84832 65736 84896
rect 65800 84832 65816 84896
rect 65880 84832 65896 84896
rect 65960 84832 65968 84896
rect 65648 83808 65968 84832
rect 65648 83744 65656 83808
rect 65720 83744 65736 83808
rect 65800 83744 65816 83808
rect 65880 83744 65896 83808
rect 65960 83744 65968 83808
rect 65648 82720 65968 83744
rect 65648 82656 65656 82720
rect 65720 82656 65736 82720
rect 65800 82656 65816 82720
rect 65880 82656 65896 82720
rect 65960 82656 65968 82720
rect 65648 81632 65968 82656
rect 65648 81568 65656 81632
rect 65720 81568 65736 81632
rect 65800 81568 65816 81632
rect 65880 81568 65896 81632
rect 65960 81568 65968 81632
rect 65648 80544 65968 81568
rect 65648 80480 65656 80544
rect 65720 80480 65736 80544
rect 65800 80480 65816 80544
rect 65880 80480 65896 80544
rect 65960 80480 65968 80544
rect 65648 79456 65968 80480
rect 65648 79392 65656 79456
rect 65720 79392 65736 79456
rect 65800 79392 65816 79456
rect 65880 79392 65896 79456
rect 65960 79392 65968 79456
rect 65648 78368 65968 79392
rect 65648 78304 65656 78368
rect 65720 78304 65736 78368
rect 65800 78304 65816 78368
rect 65880 78304 65896 78368
rect 65960 78304 65968 78368
rect 65648 77280 65968 78304
rect 65648 77216 65656 77280
rect 65720 77216 65736 77280
rect 65800 77216 65816 77280
rect 65880 77216 65896 77280
rect 65960 77216 65968 77280
rect 65648 76192 65968 77216
rect 65648 76128 65656 76192
rect 65720 76128 65736 76192
rect 65800 76128 65816 76192
rect 65880 76128 65896 76192
rect 65960 76128 65968 76192
rect 65648 75104 65968 76128
rect 65648 75040 65656 75104
rect 65720 75040 65736 75104
rect 65800 75040 65816 75104
rect 65880 75040 65896 75104
rect 65960 75040 65968 75104
rect 65648 74016 65968 75040
rect 65648 73952 65656 74016
rect 65720 73952 65736 74016
rect 65800 73952 65816 74016
rect 65880 73952 65896 74016
rect 65960 73952 65968 74016
rect 65648 72928 65968 73952
rect 65648 72864 65656 72928
rect 65720 72864 65736 72928
rect 65800 72864 65816 72928
rect 65880 72864 65896 72928
rect 65960 72864 65968 72928
rect 65648 71840 65968 72864
rect 65648 71776 65656 71840
rect 65720 71776 65736 71840
rect 65800 71776 65816 71840
rect 65880 71776 65896 71840
rect 65960 71776 65968 71840
rect 65648 70752 65968 71776
rect 65648 70688 65656 70752
rect 65720 70688 65736 70752
rect 65800 70688 65816 70752
rect 65880 70688 65896 70752
rect 65960 70688 65968 70752
rect 65648 69664 65968 70688
rect 65648 69600 65656 69664
rect 65720 69600 65736 69664
rect 65800 69600 65816 69664
rect 65880 69600 65896 69664
rect 65960 69600 65968 69664
rect 65648 68576 65968 69600
rect 65648 68512 65656 68576
rect 65720 68512 65736 68576
rect 65800 68512 65816 68576
rect 65880 68512 65896 68576
rect 65960 68512 65968 68576
rect 65648 67488 65968 68512
rect 65648 67424 65656 67488
rect 65720 67424 65736 67488
rect 65800 67424 65816 67488
rect 65880 67424 65896 67488
rect 65960 67424 65968 67488
rect 65648 66400 65968 67424
rect 65648 66336 65656 66400
rect 65720 66336 65736 66400
rect 65800 66336 65816 66400
rect 65880 66336 65896 66400
rect 65960 66336 65968 66400
rect 65648 65312 65968 66336
rect 65648 65248 65656 65312
rect 65720 65248 65736 65312
rect 65800 65248 65816 65312
rect 65880 65248 65896 65312
rect 65960 65248 65968 65312
rect 65648 64224 65968 65248
rect 65648 64160 65656 64224
rect 65720 64160 65736 64224
rect 65800 64160 65816 64224
rect 65880 64160 65896 64224
rect 65960 64160 65968 64224
rect 65648 63136 65968 64160
rect 65648 63072 65656 63136
rect 65720 63072 65736 63136
rect 65800 63072 65816 63136
rect 65880 63072 65896 63136
rect 65960 63072 65968 63136
rect 65648 62048 65968 63072
rect 65648 61984 65656 62048
rect 65720 61984 65736 62048
rect 65800 61984 65816 62048
rect 65880 61984 65896 62048
rect 65960 61984 65968 62048
rect 65648 60960 65968 61984
rect 65648 60896 65656 60960
rect 65720 60896 65736 60960
rect 65800 60896 65816 60960
rect 65880 60896 65896 60960
rect 65960 60896 65968 60960
rect 65648 59872 65968 60896
rect 65648 59808 65656 59872
rect 65720 59808 65736 59872
rect 65800 59808 65816 59872
rect 65880 59808 65896 59872
rect 65960 59808 65968 59872
rect 65648 58784 65968 59808
rect 65648 58720 65656 58784
rect 65720 58720 65736 58784
rect 65800 58720 65816 58784
rect 65880 58720 65896 58784
rect 65960 58720 65968 58784
rect 65648 57696 65968 58720
rect 65648 57632 65656 57696
rect 65720 57632 65736 57696
rect 65800 57632 65816 57696
rect 65880 57632 65896 57696
rect 65960 57632 65968 57696
rect 65648 56608 65968 57632
rect 65648 56544 65656 56608
rect 65720 56544 65736 56608
rect 65800 56544 65816 56608
rect 65880 56544 65896 56608
rect 65960 56544 65968 56608
rect 65648 55520 65968 56544
rect 65648 55456 65656 55520
rect 65720 55456 65736 55520
rect 65800 55456 65816 55520
rect 65880 55456 65896 55520
rect 65960 55456 65968 55520
rect 65648 54432 65968 55456
rect 65648 54368 65656 54432
rect 65720 54368 65736 54432
rect 65800 54368 65816 54432
rect 65880 54368 65896 54432
rect 65960 54368 65968 54432
rect 65648 53344 65968 54368
rect 65648 53280 65656 53344
rect 65720 53280 65736 53344
rect 65800 53280 65816 53344
rect 65880 53280 65896 53344
rect 65960 53280 65968 53344
rect 65648 52256 65968 53280
rect 65648 52192 65656 52256
rect 65720 52192 65736 52256
rect 65800 52192 65816 52256
rect 65880 52192 65896 52256
rect 65960 52192 65968 52256
rect 65648 51168 65968 52192
rect 65648 51104 65656 51168
rect 65720 51104 65736 51168
rect 65800 51104 65816 51168
rect 65880 51104 65896 51168
rect 65960 51104 65968 51168
rect 65648 50080 65968 51104
rect 65648 50016 65656 50080
rect 65720 50016 65736 50080
rect 65800 50016 65816 50080
rect 65880 50016 65896 50080
rect 65960 50016 65968 50080
rect 65648 48992 65968 50016
rect 65648 48928 65656 48992
rect 65720 48928 65736 48992
rect 65800 48928 65816 48992
rect 65880 48928 65896 48992
rect 65960 48928 65968 48992
rect 65648 47904 65968 48928
rect 65648 47840 65656 47904
rect 65720 47840 65736 47904
rect 65800 47840 65816 47904
rect 65880 47840 65896 47904
rect 65960 47840 65968 47904
rect 65648 46816 65968 47840
rect 65648 46752 65656 46816
rect 65720 46752 65736 46816
rect 65800 46752 65816 46816
rect 65880 46752 65896 46816
rect 65960 46752 65968 46816
rect 65648 45728 65968 46752
rect 65648 45664 65656 45728
rect 65720 45664 65736 45728
rect 65800 45664 65816 45728
rect 65880 45664 65896 45728
rect 65960 45664 65968 45728
rect 65648 44640 65968 45664
rect 65648 44576 65656 44640
rect 65720 44576 65736 44640
rect 65800 44576 65816 44640
rect 65880 44576 65896 44640
rect 65960 44576 65968 44640
rect 65648 43552 65968 44576
rect 65648 43488 65656 43552
rect 65720 43488 65736 43552
rect 65800 43488 65816 43552
rect 65880 43488 65896 43552
rect 65960 43488 65968 43552
rect 65648 42464 65968 43488
rect 65648 42400 65656 42464
rect 65720 42400 65736 42464
rect 65800 42400 65816 42464
rect 65880 42400 65896 42464
rect 65960 42400 65968 42464
rect 65648 41376 65968 42400
rect 65648 41312 65656 41376
rect 65720 41312 65736 41376
rect 65800 41312 65816 41376
rect 65880 41312 65896 41376
rect 65960 41312 65968 41376
rect 65648 40288 65968 41312
rect 65648 40224 65656 40288
rect 65720 40224 65736 40288
rect 65800 40224 65816 40288
rect 65880 40224 65896 40288
rect 65960 40224 65968 40288
rect 65648 39200 65968 40224
rect 65648 39136 65656 39200
rect 65720 39136 65736 39200
rect 65800 39136 65816 39200
rect 65880 39136 65896 39200
rect 65960 39136 65968 39200
rect 65648 38112 65968 39136
rect 65648 38048 65656 38112
rect 65720 38048 65736 38112
rect 65800 38048 65816 38112
rect 65880 38048 65896 38112
rect 65960 38048 65968 38112
rect 65648 37024 65968 38048
rect 65648 36960 65656 37024
rect 65720 36960 65736 37024
rect 65800 36960 65816 37024
rect 65880 36960 65896 37024
rect 65960 36960 65968 37024
rect 65648 35936 65968 36960
rect 65648 35872 65656 35936
rect 65720 35872 65736 35936
rect 65800 35872 65816 35936
rect 65880 35872 65896 35936
rect 65960 35872 65968 35936
rect 65648 34848 65968 35872
rect 65648 34784 65656 34848
rect 65720 34784 65736 34848
rect 65800 34784 65816 34848
rect 65880 34784 65896 34848
rect 65960 34784 65968 34848
rect 65648 33760 65968 34784
rect 65648 33696 65656 33760
rect 65720 33696 65736 33760
rect 65800 33696 65816 33760
rect 65880 33696 65896 33760
rect 65960 33696 65968 33760
rect 65648 32672 65968 33696
rect 65648 32608 65656 32672
rect 65720 32608 65736 32672
rect 65800 32608 65816 32672
rect 65880 32608 65896 32672
rect 65960 32608 65968 32672
rect 65648 31584 65968 32608
rect 65648 31520 65656 31584
rect 65720 31520 65736 31584
rect 65800 31520 65816 31584
rect 65880 31520 65896 31584
rect 65960 31520 65968 31584
rect 65648 30496 65968 31520
rect 65648 30432 65656 30496
rect 65720 30432 65736 30496
rect 65800 30432 65816 30496
rect 65880 30432 65896 30496
rect 65960 30432 65968 30496
rect 65648 29408 65968 30432
rect 65648 29344 65656 29408
rect 65720 29344 65736 29408
rect 65800 29344 65816 29408
rect 65880 29344 65896 29408
rect 65960 29344 65968 29408
rect 65648 28320 65968 29344
rect 65648 28256 65656 28320
rect 65720 28256 65736 28320
rect 65800 28256 65816 28320
rect 65880 28256 65896 28320
rect 65960 28256 65968 28320
rect 65648 27232 65968 28256
rect 65648 27168 65656 27232
rect 65720 27168 65736 27232
rect 65800 27168 65816 27232
rect 65880 27168 65896 27232
rect 65960 27168 65968 27232
rect 65648 26144 65968 27168
rect 65648 26080 65656 26144
rect 65720 26080 65736 26144
rect 65800 26080 65816 26144
rect 65880 26080 65896 26144
rect 65960 26080 65968 26144
rect 65648 25056 65968 26080
rect 65648 24992 65656 25056
rect 65720 24992 65736 25056
rect 65800 24992 65816 25056
rect 65880 24992 65896 25056
rect 65960 24992 65968 25056
rect 65648 23968 65968 24992
rect 65648 23904 65656 23968
rect 65720 23904 65736 23968
rect 65800 23904 65816 23968
rect 65880 23904 65896 23968
rect 65960 23904 65968 23968
rect 65648 22880 65968 23904
rect 65648 22816 65656 22880
rect 65720 22816 65736 22880
rect 65800 22816 65816 22880
rect 65880 22816 65896 22880
rect 65960 22816 65968 22880
rect 65648 21792 65968 22816
rect 65648 21728 65656 21792
rect 65720 21728 65736 21792
rect 65800 21728 65816 21792
rect 65880 21728 65896 21792
rect 65960 21728 65968 21792
rect 65648 20704 65968 21728
rect 65648 20640 65656 20704
rect 65720 20640 65736 20704
rect 65800 20640 65816 20704
rect 65880 20640 65896 20704
rect 65960 20640 65968 20704
rect 65648 19616 65968 20640
rect 65648 19552 65656 19616
rect 65720 19552 65736 19616
rect 65800 19552 65816 19616
rect 65880 19552 65896 19616
rect 65960 19552 65968 19616
rect 65648 18528 65968 19552
rect 65648 18464 65656 18528
rect 65720 18464 65736 18528
rect 65800 18464 65816 18528
rect 65880 18464 65896 18528
rect 65960 18464 65968 18528
rect 65648 17440 65968 18464
rect 65648 17376 65656 17440
rect 65720 17376 65736 17440
rect 65800 17376 65816 17440
rect 65880 17376 65896 17440
rect 65960 17376 65968 17440
rect 65648 16352 65968 17376
rect 65648 16288 65656 16352
rect 65720 16288 65736 16352
rect 65800 16288 65816 16352
rect 65880 16288 65896 16352
rect 65960 16288 65968 16352
rect 65648 15264 65968 16288
rect 65648 15200 65656 15264
rect 65720 15200 65736 15264
rect 65800 15200 65816 15264
rect 65880 15200 65896 15264
rect 65960 15200 65968 15264
rect 65648 14176 65968 15200
rect 65648 14112 65656 14176
rect 65720 14112 65736 14176
rect 65800 14112 65816 14176
rect 65880 14112 65896 14176
rect 65960 14112 65968 14176
rect 65648 13088 65968 14112
rect 65648 13024 65656 13088
rect 65720 13024 65736 13088
rect 65800 13024 65816 13088
rect 65880 13024 65896 13088
rect 65960 13024 65968 13088
rect 65648 12000 65968 13024
rect 65648 11936 65656 12000
rect 65720 11936 65736 12000
rect 65800 11936 65816 12000
rect 65880 11936 65896 12000
rect 65960 11936 65968 12000
rect 65648 10912 65968 11936
rect 65648 10848 65656 10912
rect 65720 10848 65736 10912
rect 65800 10848 65816 10912
rect 65880 10848 65896 10912
rect 65960 10848 65968 10912
rect 65648 9824 65968 10848
rect 65648 9760 65656 9824
rect 65720 9760 65736 9824
rect 65800 9760 65816 9824
rect 65880 9760 65896 9824
rect 65960 9760 65968 9824
rect 65648 8736 65968 9760
rect 65648 8672 65656 8736
rect 65720 8672 65736 8736
rect 65800 8672 65816 8736
rect 65880 8672 65896 8736
rect 65960 8672 65968 8736
rect 65648 7648 65968 8672
rect 65648 7584 65656 7648
rect 65720 7584 65736 7648
rect 65800 7584 65816 7648
rect 65880 7584 65896 7648
rect 65960 7584 65968 7648
rect 65648 6560 65968 7584
rect 65648 6496 65656 6560
rect 65720 6496 65736 6560
rect 65800 6496 65816 6560
rect 65880 6496 65896 6560
rect 65960 6496 65968 6560
rect 65648 5472 65968 6496
rect 65648 5408 65656 5472
rect 65720 5408 65736 5472
rect 65800 5408 65816 5472
rect 65880 5408 65896 5472
rect 65960 5408 65968 5472
rect 65648 4384 65968 5408
rect 65648 4320 65656 4384
rect 65720 4320 65736 4384
rect 65800 4320 65816 4384
rect 65880 4320 65896 4384
rect 65960 4320 65968 4384
rect 65648 3296 65968 4320
rect 65648 3232 65656 3296
rect 65720 3232 65736 3296
rect 65800 3232 65816 3296
rect 65880 3232 65896 3296
rect 65960 3232 65968 3296
rect 65648 2208 65968 3232
rect 65648 2144 65656 2208
rect 65720 2144 65736 2208
rect 65800 2144 65816 2208
rect 65880 2144 65896 2208
rect 65960 2144 65968 2208
rect 66308 2176 66628 117504
rect 66968 2176 67288 117504
rect 67628 2176 67948 117504
rect 81008 116992 81328 117552
rect 96368 117536 96688 117552
rect 81008 116928 81016 116992
rect 81080 116928 81096 116992
rect 81160 116928 81176 116992
rect 81240 116928 81256 116992
rect 81320 116928 81328 116992
rect 81008 115904 81328 116928
rect 81008 115840 81016 115904
rect 81080 115840 81096 115904
rect 81160 115840 81176 115904
rect 81240 115840 81256 115904
rect 81320 115840 81328 115904
rect 81008 114816 81328 115840
rect 81008 114752 81016 114816
rect 81080 114752 81096 114816
rect 81160 114752 81176 114816
rect 81240 114752 81256 114816
rect 81320 114752 81328 114816
rect 81008 113728 81328 114752
rect 81008 113664 81016 113728
rect 81080 113664 81096 113728
rect 81160 113664 81176 113728
rect 81240 113664 81256 113728
rect 81320 113664 81328 113728
rect 81008 112640 81328 113664
rect 81008 112576 81016 112640
rect 81080 112576 81096 112640
rect 81160 112576 81176 112640
rect 81240 112576 81256 112640
rect 81320 112576 81328 112640
rect 81008 111552 81328 112576
rect 81008 111488 81016 111552
rect 81080 111488 81096 111552
rect 81160 111488 81176 111552
rect 81240 111488 81256 111552
rect 81320 111488 81328 111552
rect 81008 110464 81328 111488
rect 81008 110400 81016 110464
rect 81080 110400 81096 110464
rect 81160 110400 81176 110464
rect 81240 110400 81256 110464
rect 81320 110400 81328 110464
rect 81008 109376 81328 110400
rect 81008 109312 81016 109376
rect 81080 109312 81096 109376
rect 81160 109312 81176 109376
rect 81240 109312 81256 109376
rect 81320 109312 81328 109376
rect 81008 108288 81328 109312
rect 81008 108224 81016 108288
rect 81080 108224 81096 108288
rect 81160 108224 81176 108288
rect 81240 108224 81256 108288
rect 81320 108224 81328 108288
rect 81008 107200 81328 108224
rect 81008 107136 81016 107200
rect 81080 107136 81096 107200
rect 81160 107136 81176 107200
rect 81240 107136 81256 107200
rect 81320 107136 81328 107200
rect 81008 106112 81328 107136
rect 81008 106048 81016 106112
rect 81080 106048 81096 106112
rect 81160 106048 81176 106112
rect 81240 106048 81256 106112
rect 81320 106048 81328 106112
rect 81008 105024 81328 106048
rect 81008 104960 81016 105024
rect 81080 104960 81096 105024
rect 81160 104960 81176 105024
rect 81240 104960 81256 105024
rect 81320 104960 81328 105024
rect 81008 103936 81328 104960
rect 81008 103872 81016 103936
rect 81080 103872 81096 103936
rect 81160 103872 81176 103936
rect 81240 103872 81256 103936
rect 81320 103872 81328 103936
rect 81008 102848 81328 103872
rect 81008 102784 81016 102848
rect 81080 102784 81096 102848
rect 81160 102784 81176 102848
rect 81240 102784 81256 102848
rect 81320 102784 81328 102848
rect 81008 101760 81328 102784
rect 81008 101696 81016 101760
rect 81080 101696 81096 101760
rect 81160 101696 81176 101760
rect 81240 101696 81256 101760
rect 81320 101696 81328 101760
rect 81008 100672 81328 101696
rect 81008 100608 81016 100672
rect 81080 100608 81096 100672
rect 81160 100608 81176 100672
rect 81240 100608 81256 100672
rect 81320 100608 81328 100672
rect 81008 99584 81328 100608
rect 81008 99520 81016 99584
rect 81080 99520 81096 99584
rect 81160 99520 81176 99584
rect 81240 99520 81256 99584
rect 81320 99520 81328 99584
rect 81008 98496 81328 99520
rect 81008 98432 81016 98496
rect 81080 98432 81096 98496
rect 81160 98432 81176 98496
rect 81240 98432 81256 98496
rect 81320 98432 81328 98496
rect 81008 97408 81328 98432
rect 81008 97344 81016 97408
rect 81080 97344 81096 97408
rect 81160 97344 81176 97408
rect 81240 97344 81256 97408
rect 81320 97344 81328 97408
rect 81008 96320 81328 97344
rect 81008 96256 81016 96320
rect 81080 96256 81096 96320
rect 81160 96256 81176 96320
rect 81240 96256 81256 96320
rect 81320 96256 81328 96320
rect 81008 95232 81328 96256
rect 81008 95168 81016 95232
rect 81080 95168 81096 95232
rect 81160 95168 81176 95232
rect 81240 95168 81256 95232
rect 81320 95168 81328 95232
rect 81008 94144 81328 95168
rect 81008 94080 81016 94144
rect 81080 94080 81096 94144
rect 81160 94080 81176 94144
rect 81240 94080 81256 94144
rect 81320 94080 81328 94144
rect 81008 93056 81328 94080
rect 81008 92992 81016 93056
rect 81080 92992 81096 93056
rect 81160 92992 81176 93056
rect 81240 92992 81256 93056
rect 81320 92992 81328 93056
rect 81008 91968 81328 92992
rect 81008 91904 81016 91968
rect 81080 91904 81096 91968
rect 81160 91904 81176 91968
rect 81240 91904 81256 91968
rect 81320 91904 81328 91968
rect 81008 90880 81328 91904
rect 81008 90816 81016 90880
rect 81080 90816 81096 90880
rect 81160 90816 81176 90880
rect 81240 90816 81256 90880
rect 81320 90816 81328 90880
rect 81008 89792 81328 90816
rect 81008 89728 81016 89792
rect 81080 89728 81096 89792
rect 81160 89728 81176 89792
rect 81240 89728 81256 89792
rect 81320 89728 81328 89792
rect 81008 88704 81328 89728
rect 81008 88640 81016 88704
rect 81080 88640 81096 88704
rect 81160 88640 81176 88704
rect 81240 88640 81256 88704
rect 81320 88640 81328 88704
rect 81008 87616 81328 88640
rect 81008 87552 81016 87616
rect 81080 87552 81096 87616
rect 81160 87552 81176 87616
rect 81240 87552 81256 87616
rect 81320 87552 81328 87616
rect 81008 86528 81328 87552
rect 81008 86464 81016 86528
rect 81080 86464 81096 86528
rect 81160 86464 81176 86528
rect 81240 86464 81256 86528
rect 81320 86464 81328 86528
rect 81008 85440 81328 86464
rect 81008 85376 81016 85440
rect 81080 85376 81096 85440
rect 81160 85376 81176 85440
rect 81240 85376 81256 85440
rect 81320 85376 81328 85440
rect 81008 84352 81328 85376
rect 81008 84288 81016 84352
rect 81080 84288 81096 84352
rect 81160 84288 81176 84352
rect 81240 84288 81256 84352
rect 81320 84288 81328 84352
rect 81008 83264 81328 84288
rect 81008 83200 81016 83264
rect 81080 83200 81096 83264
rect 81160 83200 81176 83264
rect 81240 83200 81256 83264
rect 81320 83200 81328 83264
rect 81008 82176 81328 83200
rect 81008 82112 81016 82176
rect 81080 82112 81096 82176
rect 81160 82112 81176 82176
rect 81240 82112 81256 82176
rect 81320 82112 81328 82176
rect 81008 81088 81328 82112
rect 81008 81024 81016 81088
rect 81080 81024 81096 81088
rect 81160 81024 81176 81088
rect 81240 81024 81256 81088
rect 81320 81024 81328 81088
rect 81008 80000 81328 81024
rect 81008 79936 81016 80000
rect 81080 79936 81096 80000
rect 81160 79936 81176 80000
rect 81240 79936 81256 80000
rect 81320 79936 81328 80000
rect 81008 78912 81328 79936
rect 81008 78848 81016 78912
rect 81080 78848 81096 78912
rect 81160 78848 81176 78912
rect 81240 78848 81256 78912
rect 81320 78848 81328 78912
rect 81008 77824 81328 78848
rect 81008 77760 81016 77824
rect 81080 77760 81096 77824
rect 81160 77760 81176 77824
rect 81240 77760 81256 77824
rect 81320 77760 81328 77824
rect 81008 76736 81328 77760
rect 81008 76672 81016 76736
rect 81080 76672 81096 76736
rect 81160 76672 81176 76736
rect 81240 76672 81256 76736
rect 81320 76672 81328 76736
rect 81008 75648 81328 76672
rect 81008 75584 81016 75648
rect 81080 75584 81096 75648
rect 81160 75584 81176 75648
rect 81240 75584 81256 75648
rect 81320 75584 81328 75648
rect 81008 74560 81328 75584
rect 81008 74496 81016 74560
rect 81080 74496 81096 74560
rect 81160 74496 81176 74560
rect 81240 74496 81256 74560
rect 81320 74496 81328 74560
rect 81008 73472 81328 74496
rect 81008 73408 81016 73472
rect 81080 73408 81096 73472
rect 81160 73408 81176 73472
rect 81240 73408 81256 73472
rect 81320 73408 81328 73472
rect 81008 72384 81328 73408
rect 81008 72320 81016 72384
rect 81080 72320 81096 72384
rect 81160 72320 81176 72384
rect 81240 72320 81256 72384
rect 81320 72320 81328 72384
rect 81008 71296 81328 72320
rect 81008 71232 81016 71296
rect 81080 71232 81096 71296
rect 81160 71232 81176 71296
rect 81240 71232 81256 71296
rect 81320 71232 81328 71296
rect 81008 70208 81328 71232
rect 81008 70144 81016 70208
rect 81080 70144 81096 70208
rect 81160 70144 81176 70208
rect 81240 70144 81256 70208
rect 81320 70144 81328 70208
rect 81008 69120 81328 70144
rect 81008 69056 81016 69120
rect 81080 69056 81096 69120
rect 81160 69056 81176 69120
rect 81240 69056 81256 69120
rect 81320 69056 81328 69120
rect 81008 68032 81328 69056
rect 81008 67968 81016 68032
rect 81080 67968 81096 68032
rect 81160 67968 81176 68032
rect 81240 67968 81256 68032
rect 81320 67968 81328 68032
rect 81008 66944 81328 67968
rect 81008 66880 81016 66944
rect 81080 66880 81096 66944
rect 81160 66880 81176 66944
rect 81240 66880 81256 66944
rect 81320 66880 81328 66944
rect 81008 65856 81328 66880
rect 81008 65792 81016 65856
rect 81080 65792 81096 65856
rect 81160 65792 81176 65856
rect 81240 65792 81256 65856
rect 81320 65792 81328 65856
rect 81008 64768 81328 65792
rect 81008 64704 81016 64768
rect 81080 64704 81096 64768
rect 81160 64704 81176 64768
rect 81240 64704 81256 64768
rect 81320 64704 81328 64768
rect 81008 63680 81328 64704
rect 81008 63616 81016 63680
rect 81080 63616 81096 63680
rect 81160 63616 81176 63680
rect 81240 63616 81256 63680
rect 81320 63616 81328 63680
rect 81008 62592 81328 63616
rect 81008 62528 81016 62592
rect 81080 62528 81096 62592
rect 81160 62528 81176 62592
rect 81240 62528 81256 62592
rect 81320 62528 81328 62592
rect 81008 61504 81328 62528
rect 81008 61440 81016 61504
rect 81080 61440 81096 61504
rect 81160 61440 81176 61504
rect 81240 61440 81256 61504
rect 81320 61440 81328 61504
rect 81008 60416 81328 61440
rect 81008 60352 81016 60416
rect 81080 60352 81096 60416
rect 81160 60352 81176 60416
rect 81240 60352 81256 60416
rect 81320 60352 81328 60416
rect 81008 59328 81328 60352
rect 81008 59264 81016 59328
rect 81080 59264 81096 59328
rect 81160 59264 81176 59328
rect 81240 59264 81256 59328
rect 81320 59264 81328 59328
rect 81008 58240 81328 59264
rect 81008 58176 81016 58240
rect 81080 58176 81096 58240
rect 81160 58176 81176 58240
rect 81240 58176 81256 58240
rect 81320 58176 81328 58240
rect 81008 57152 81328 58176
rect 81008 57088 81016 57152
rect 81080 57088 81096 57152
rect 81160 57088 81176 57152
rect 81240 57088 81256 57152
rect 81320 57088 81328 57152
rect 81008 56064 81328 57088
rect 81008 56000 81016 56064
rect 81080 56000 81096 56064
rect 81160 56000 81176 56064
rect 81240 56000 81256 56064
rect 81320 56000 81328 56064
rect 81008 54976 81328 56000
rect 81008 54912 81016 54976
rect 81080 54912 81096 54976
rect 81160 54912 81176 54976
rect 81240 54912 81256 54976
rect 81320 54912 81328 54976
rect 81008 53888 81328 54912
rect 81008 53824 81016 53888
rect 81080 53824 81096 53888
rect 81160 53824 81176 53888
rect 81240 53824 81256 53888
rect 81320 53824 81328 53888
rect 81008 52800 81328 53824
rect 81008 52736 81016 52800
rect 81080 52736 81096 52800
rect 81160 52736 81176 52800
rect 81240 52736 81256 52800
rect 81320 52736 81328 52800
rect 81008 51712 81328 52736
rect 81008 51648 81016 51712
rect 81080 51648 81096 51712
rect 81160 51648 81176 51712
rect 81240 51648 81256 51712
rect 81320 51648 81328 51712
rect 81008 50624 81328 51648
rect 81008 50560 81016 50624
rect 81080 50560 81096 50624
rect 81160 50560 81176 50624
rect 81240 50560 81256 50624
rect 81320 50560 81328 50624
rect 81008 49536 81328 50560
rect 81008 49472 81016 49536
rect 81080 49472 81096 49536
rect 81160 49472 81176 49536
rect 81240 49472 81256 49536
rect 81320 49472 81328 49536
rect 81008 48448 81328 49472
rect 81008 48384 81016 48448
rect 81080 48384 81096 48448
rect 81160 48384 81176 48448
rect 81240 48384 81256 48448
rect 81320 48384 81328 48448
rect 81008 47360 81328 48384
rect 81008 47296 81016 47360
rect 81080 47296 81096 47360
rect 81160 47296 81176 47360
rect 81240 47296 81256 47360
rect 81320 47296 81328 47360
rect 81008 46272 81328 47296
rect 81008 46208 81016 46272
rect 81080 46208 81096 46272
rect 81160 46208 81176 46272
rect 81240 46208 81256 46272
rect 81320 46208 81328 46272
rect 81008 45184 81328 46208
rect 81008 45120 81016 45184
rect 81080 45120 81096 45184
rect 81160 45120 81176 45184
rect 81240 45120 81256 45184
rect 81320 45120 81328 45184
rect 81008 44096 81328 45120
rect 81008 44032 81016 44096
rect 81080 44032 81096 44096
rect 81160 44032 81176 44096
rect 81240 44032 81256 44096
rect 81320 44032 81328 44096
rect 81008 43008 81328 44032
rect 81008 42944 81016 43008
rect 81080 42944 81096 43008
rect 81160 42944 81176 43008
rect 81240 42944 81256 43008
rect 81320 42944 81328 43008
rect 81008 41920 81328 42944
rect 81008 41856 81016 41920
rect 81080 41856 81096 41920
rect 81160 41856 81176 41920
rect 81240 41856 81256 41920
rect 81320 41856 81328 41920
rect 81008 40832 81328 41856
rect 81008 40768 81016 40832
rect 81080 40768 81096 40832
rect 81160 40768 81176 40832
rect 81240 40768 81256 40832
rect 81320 40768 81328 40832
rect 81008 39744 81328 40768
rect 81008 39680 81016 39744
rect 81080 39680 81096 39744
rect 81160 39680 81176 39744
rect 81240 39680 81256 39744
rect 81320 39680 81328 39744
rect 81008 38656 81328 39680
rect 81008 38592 81016 38656
rect 81080 38592 81096 38656
rect 81160 38592 81176 38656
rect 81240 38592 81256 38656
rect 81320 38592 81328 38656
rect 81008 37568 81328 38592
rect 81008 37504 81016 37568
rect 81080 37504 81096 37568
rect 81160 37504 81176 37568
rect 81240 37504 81256 37568
rect 81320 37504 81328 37568
rect 81008 36480 81328 37504
rect 81008 36416 81016 36480
rect 81080 36416 81096 36480
rect 81160 36416 81176 36480
rect 81240 36416 81256 36480
rect 81320 36416 81328 36480
rect 81008 35392 81328 36416
rect 81008 35328 81016 35392
rect 81080 35328 81096 35392
rect 81160 35328 81176 35392
rect 81240 35328 81256 35392
rect 81320 35328 81328 35392
rect 81008 34304 81328 35328
rect 81008 34240 81016 34304
rect 81080 34240 81096 34304
rect 81160 34240 81176 34304
rect 81240 34240 81256 34304
rect 81320 34240 81328 34304
rect 81008 33216 81328 34240
rect 81008 33152 81016 33216
rect 81080 33152 81096 33216
rect 81160 33152 81176 33216
rect 81240 33152 81256 33216
rect 81320 33152 81328 33216
rect 81008 32128 81328 33152
rect 81008 32064 81016 32128
rect 81080 32064 81096 32128
rect 81160 32064 81176 32128
rect 81240 32064 81256 32128
rect 81320 32064 81328 32128
rect 81008 31040 81328 32064
rect 81008 30976 81016 31040
rect 81080 30976 81096 31040
rect 81160 30976 81176 31040
rect 81240 30976 81256 31040
rect 81320 30976 81328 31040
rect 81008 29952 81328 30976
rect 81008 29888 81016 29952
rect 81080 29888 81096 29952
rect 81160 29888 81176 29952
rect 81240 29888 81256 29952
rect 81320 29888 81328 29952
rect 81008 28864 81328 29888
rect 81008 28800 81016 28864
rect 81080 28800 81096 28864
rect 81160 28800 81176 28864
rect 81240 28800 81256 28864
rect 81320 28800 81328 28864
rect 81008 27776 81328 28800
rect 81008 27712 81016 27776
rect 81080 27712 81096 27776
rect 81160 27712 81176 27776
rect 81240 27712 81256 27776
rect 81320 27712 81328 27776
rect 81008 26688 81328 27712
rect 81008 26624 81016 26688
rect 81080 26624 81096 26688
rect 81160 26624 81176 26688
rect 81240 26624 81256 26688
rect 81320 26624 81328 26688
rect 81008 25600 81328 26624
rect 81008 25536 81016 25600
rect 81080 25536 81096 25600
rect 81160 25536 81176 25600
rect 81240 25536 81256 25600
rect 81320 25536 81328 25600
rect 81008 24512 81328 25536
rect 81008 24448 81016 24512
rect 81080 24448 81096 24512
rect 81160 24448 81176 24512
rect 81240 24448 81256 24512
rect 81320 24448 81328 24512
rect 81008 23424 81328 24448
rect 81008 23360 81016 23424
rect 81080 23360 81096 23424
rect 81160 23360 81176 23424
rect 81240 23360 81256 23424
rect 81320 23360 81328 23424
rect 81008 22336 81328 23360
rect 81008 22272 81016 22336
rect 81080 22272 81096 22336
rect 81160 22272 81176 22336
rect 81240 22272 81256 22336
rect 81320 22272 81328 22336
rect 81008 21248 81328 22272
rect 81008 21184 81016 21248
rect 81080 21184 81096 21248
rect 81160 21184 81176 21248
rect 81240 21184 81256 21248
rect 81320 21184 81328 21248
rect 81008 20160 81328 21184
rect 81008 20096 81016 20160
rect 81080 20096 81096 20160
rect 81160 20096 81176 20160
rect 81240 20096 81256 20160
rect 81320 20096 81328 20160
rect 81008 19072 81328 20096
rect 81008 19008 81016 19072
rect 81080 19008 81096 19072
rect 81160 19008 81176 19072
rect 81240 19008 81256 19072
rect 81320 19008 81328 19072
rect 81008 17984 81328 19008
rect 81008 17920 81016 17984
rect 81080 17920 81096 17984
rect 81160 17920 81176 17984
rect 81240 17920 81256 17984
rect 81320 17920 81328 17984
rect 81008 16896 81328 17920
rect 81008 16832 81016 16896
rect 81080 16832 81096 16896
rect 81160 16832 81176 16896
rect 81240 16832 81256 16896
rect 81320 16832 81328 16896
rect 81008 15808 81328 16832
rect 81008 15744 81016 15808
rect 81080 15744 81096 15808
rect 81160 15744 81176 15808
rect 81240 15744 81256 15808
rect 81320 15744 81328 15808
rect 81008 14720 81328 15744
rect 81008 14656 81016 14720
rect 81080 14656 81096 14720
rect 81160 14656 81176 14720
rect 81240 14656 81256 14720
rect 81320 14656 81328 14720
rect 81008 13632 81328 14656
rect 81008 13568 81016 13632
rect 81080 13568 81096 13632
rect 81160 13568 81176 13632
rect 81240 13568 81256 13632
rect 81320 13568 81328 13632
rect 81008 12544 81328 13568
rect 81008 12480 81016 12544
rect 81080 12480 81096 12544
rect 81160 12480 81176 12544
rect 81240 12480 81256 12544
rect 81320 12480 81328 12544
rect 81008 11456 81328 12480
rect 81008 11392 81016 11456
rect 81080 11392 81096 11456
rect 81160 11392 81176 11456
rect 81240 11392 81256 11456
rect 81320 11392 81328 11456
rect 81008 10368 81328 11392
rect 81008 10304 81016 10368
rect 81080 10304 81096 10368
rect 81160 10304 81176 10368
rect 81240 10304 81256 10368
rect 81320 10304 81328 10368
rect 81008 9280 81328 10304
rect 81008 9216 81016 9280
rect 81080 9216 81096 9280
rect 81160 9216 81176 9280
rect 81240 9216 81256 9280
rect 81320 9216 81328 9280
rect 81008 8192 81328 9216
rect 81008 8128 81016 8192
rect 81080 8128 81096 8192
rect 81160 8128 81176 8192
rect 81240 8128 81256 8192
rect 81320 8128 81328 8192
rect 81008 7104 81328 8128
rect 81008 7040 81016 7104
rect 81080 7040 81096 7104
rect 81160 7040 81176 7104
rect 81240 7040 81256 7104
rect 81320 7040 81328 7104
rect 81008 6016 81328 7040
rect 81008 5952 81016 6016
rect 81080 5952 81096 6016
rect 81160 5952 81176 6016
rect 81240 5952 81256 6016
rect 81320 5952 81328 6016
rect 81008 4928 81328 5952
rect 81008 4864 81016 4928
rect 81080 4864 81096 4928
rect 81160 4864 81176 4928
rect 81240 4864 81256 4928
rect 81320 4864 81328 4928
rect 80651 4724 80717 4725
rect 80651 4660 80652 4724
rect 80716 4660 80717 4724
rect 80651 4659 80717 4660
rect 80654 2821 80714 4659
rect 81008 3840 81328 4864
rect 81008 3776 81016 3840
rect 81080 3776 81096 3840
rect 81160 3776 81176 3840
rect 81240 3776 81256 3840
rect 81320 3776 81328 3840
rect 80651 2820 80717 2821
rect 80651 2756 80652 2820
rect 80716 2756 80717 2820
rect 80651 2755 80717 2756
rect 81008 2752 81328 3776
rect 81008 2688 81016 2752
rect 81080 2688 81096 2752
rect 81160 2688 81176 2752
rect 81240 2688 81256 2752
rect 81320 2688 81328 2752
rect 65648 2128 65968 2144
rect 81008 2128 81328 2688
rect 81668 2176 81988 117504
rect 82328 2176 82648 117504
rect 82988 2176 83308 117504
rect 96368 117472 96376 117536
rect 96440 117472 96456 117536
rect 96520 117472 96536 117536
rect 96600 117472 96616 117536
rect 96680 117472 96688 117536
rect 96368 116448 96688 117472
rect 96368 116384 96376 116448
rect 96440 116384 96456 116448
rect 96520 116384 96536 116448
rect 96600 116384 96616 116448
rect 96680 116384 96688 116448
rect 96368 115360 96688 116384
rect 96368 115296 96376 115360
rect 96440 115296 96456 115360
rect 96520 115296 96536 115360
rect 96600 115296 96616 115360
rect 96680 115296 96688 115360
rect 96368 114272 96688 115296
rect 96368 114208 96376 114272
rect 96440 114208 96456 114272
rect 96520 114208 96536 114272
rect 96600 114208 96616 114272
rect 96680 114208 96688 114272
rect 96368 113184 96688 114208
rect 96368 113120 96376 113184
rect 96440 113120 96456 113184
rect 96520 113120 96536 113184
rect 96600 113120 96616 113184
rect 96680 113120 96688 113184
rect 96368 112096 96688 113120
rect 96368 112032 96376 112096
rect 96440 112032 96456 112096
rect 96520 112032 96536 112096
rect 96600 112032 96616 112096
rect 96680 112032 96688 112096
rect 96368 111008 96688 112032
rect 96368 110944 96376 111008
rect 96440 110944 96456 111008
rect 96520 110944 96536 111008
rect 96600 110944 96616 111008
rect 96680 110944 96688 111008
rect 96368 109920 96688 110944
rect 96368 109856 96376 109920
rect 96440 109856 96456 109920
rect 96520 109856 96536 109920
rect 96600 109856 96616 109920
rect 96680 109856 96688 109920
rect 96368 108832 96688 109856
rect 96368 108768 96376 108832
rect 96440 108768 96456 108832
rect 96520 108768 96536 108832
rect 96600 108768 96616 108832
rect 96680 108768 96688 108832
rect 96368 107744 96688 108768
rect 96368 107680 96376 107744
rect 96440 107680 96456 107744
rect 96520 107680 96536 107744
rect 96600 107680 96616 107744
rect 96680 107680 96688 107744
rect 96368 106656 96688 107680
rect 96368 106592 96376 106656
rect 96440 106592 96456 106656
rect 96520 106592 96536 106656
rect 96600 106592 96616 106656
rect 96680 106592 96688 106656
rect 96368 105568 96688 106592
rect 96368 105504 96376 105568
rect 96440 105504 96456 105568
rect 96520 105504 96536 105568
rect 96600 105504 96616 105568
rect 96680 105504 96688 105568
rect 96368 104480 96688 105504
rect 96368 104416 96376 104480
rect 96440 104416 96456 104480
rect 96520 104416 96536 104480
rect 96600 104416 96616 104480
rect 96680 104416 96688 104480
rect 96368 103392 96688 104416
rect 96368 103328 96376 103392
rect 96440 103328 96456 103392
rect 96520 103328 96536 103392
rect 96600 103328 96616 103392
rect 96680 103328 96688 103392
rect 96368 102304 96688 103328
rect 96368 102240 96376 102304
rect 96440 102240 96456 102304
rect 96520 102240 96536 102304
rect 96600 102240 96616 102304
rect 96680 102240 96688 102304
rect 96368 101216 96688 102240
rect 96368 101152 96376 101216
rect 96440 101152 96456 101216
rect 96520 101152 96536 101216
rect 96600 101152 96616 101216
rect 96680 101152 96688 101216
rect 96368 100128 96688 101152
rect 96368 100064 96376 100128
rect 96440 100064 96456 100128
rect 96520 100064 96536 100128
rect 96600 100064 96616 100128
rect 96680 100064 96688 100128
rect 96368 99040 96688 100064
rect 96368 98976 96376 99040
rect 96440 98976 96456 99040
rect 96520 98976 96536 99040
rect 96600 98976 96616 99040
rect 96680 98976 96688 99040
rect 96368 97952 96688 98976
rect 96368 97888 96376 97952
rect 96440 97888 96456 97952
rect 96520 97888 96536 97952
rect 96600 97888 96616 97952
rect 96680 97888 96688 97952
rect 96368 96864 96688 97888
rect 96368 96800 96376 96864
rect 96440 96800 96456 96864
rect 96520 96800 96536 96864
rect 96600 96800 96616 96864
rect 96680 96800 96688 96864
rect 96368 95776 96688 96800
rect 96368 95712 96376 95776
rect 96440 95712 96456 95776
rect 96520 95712 96536 95776
rect 96600 95712 96616 95776
rect 96680 95712 96688 95776
rect 96368 94688 96688 95712
rect 96368 94624 96376 94688
rect 96440 94624 96456 94688
rect 96520 94624 96536 94688
rect 96600 94624 96616 94688
rect 96680 94624 96688 94688
rect 96368 93600 96688 94624
rect 96368 93536 96376 93600
rect 96440 93536 96456 93600
rect 96520 93536 96536 93600
rect 96600 93536 96616 93600
rect 96680 93536 96688 93600
rect 96368 92512 96688 93536
rect 96368 92448 96376 92512
rect 96440 92448 96456 92512
rect 96520 92448 96536 92512
rect 96600 92448 96616 92512
rect 96680 92448 96688 92512
rect 96368 91424 96688 92448
rect 96368 91360 96376 91424
rect 96440 91360 96456 91424
rect 96520 91360 96536 91424
rect 96600 91360 96616 91424
rect 96680 91360 96688 91424
rect 96368 90336 96688 91360
rect 96368 90272 96376 90336
rect 96440 90272 96456 90336
rect 96520 90272 96536 90336
rect 96600 90272 96616 90336
rect 96680 90272 96688 90336
rect 96368 89248 96688 90272
rect 96368 89184 96376 89248
rect 96440 89184 96456 89248
rect 96520 89184 96536 89248
rect 96600 89184 96616 89248
rect 96680 89184 96688 89248
rect 96368 88160 96688 89184
rect 96368 88096 96376 88160
rect 96440 88096 96456 88160
rect 96520 88096 96536 88160
rect 96600 88096 96616 88160
rect 96680 88096 96688 88160
rect 96368 87072 96688 88096
rect 96368 87008 96376 87072
rect 96440 87008 96456 87072
rect 96520 87008 96536 87072
rect 96600 87008 96616 87072
rect 96680 87008 96688 87072
rect 96368 85984 96688 87008
rect 96368 85920 96376 85984
rect 96440 85920 96456 85984
rect 96520 85920 96536 85984
rect 96600 85920 96616 85984
rect 96680 85920 96688 85984
rect 96368 84896 96688 85920
rect 96368 84832 96376 84896
rect 96440 84832 96456 84896
rect 96520 84832 96536 84896
rect 96600 84832 96616 84896
rect 96680 84832 96688 84896
rect 96368 83808 96688 84832
rect 96368 83744 96376 83808
rect 96440 83744 96456 83808
rect 96520 83744 96536 83808
rect 96600 83744 96616 83808
rect 96680 83744 96688 83808
rect 96368 82720 96688 83744
rect 96368 82656 96376 82720
rect 96440 82656 96456 82720
rect 96520 82656 96536 82720
rect 96600 82656 96616 82720
rect 96680 82656 96688 82720
rect 96368 81632 96688 82656
rect 96368 81568 96376 81632
rect 96440 81568 96456 81632
rect 96520 81568 96536 81632
rect 96600 81568 96616 81632
rect 96680 81568 96688 81632
rect 96368 80544 96688 81568
rect 96368 80480 96376 80544
rect 96440 80480 96456 80544
rect 96520 80480 96536 80544
rect 96600 80480 96616 80544
rect 96680 80480 96688 80544
rect 96368 79456 96688 80480
rect 96368 79392 96376 79456
rect 96440 79392 96456 79456
rect 96520 79392 96536 79456
rect 96600 79392 96616 79456
rect 96680 79392 96688 79456
rect 96368 78368 96688 79392
rect 96368 78304 96376 78368
rect 96440 78304 96456 78368
rect 96520 78304 96536 78368
rect 96600 78304 96616 78368
rect 96680 78304 96688 78368
rect 96368 77280 96688 78304
rect 96368 77216 96376 77280
rect 96440 77216 96456 77280
rect 96520 77216 96536 77280
rect 96600 77216 96616 77280
rect 96680 77216 96688 77280
rect 96368 76192 96688 77216
rect 96368 76128 96376 76192
rect 96440 76128 96456 76192
rect 96520 76128 96536 76192
rect 96600 76128 96616 76192
rect 96680 76128 96688 76192
rect 96368 75104 96688 76128
rect 96368 75040 96376 75104
rect 96440 75040 96456 75104
rect 96520 75040 96536 75104
rect 96600 75040 96616 75104
rect 96680 75040 96688 75104
rect 96368 74016 96688 75040
rect 96368 73952 96376 74016
rect 96440 73952 96456 74016
rect 96520 73952 96536 74016
rect 96600 73952 96616 74016
rect 96680 73952 96688 74016
rect 96368 72928 96688 73952
rect 96368 72864 96376 72928
rect 96440 72864 96456 72928
rect 96520 72864 96536 72928
rect 96600 72864 96616 72928
rect 96680 72864 96688 72928
rect 96368 71840 96688 72864
rect 96368 71776 96376 71840
rect 96440 71776 96456 71840
rect 96520 71776 96536 71840
rect 96600 71776 96616 71840
rect 96680 71776 96688 71840
rect 96368 70752 96688 71776
rect 96368 70688 96376 70752
rect 96440 70688 96456 70752
rect 96520 70688 96536 70752
rect 96600 70688 96616 70752
rect 96680 70688 96688 70752
rect 96368 69664 96688 70688
rect 96368 69600 96376 69664
rect 96440 69600 96456 69664
rect 96520 69600 96536 69664
rect 96600 69600 96616 69664
rect 96680 69600 96688 69664
rect 96368 68576 96688 69600
rect 96368 68512 96376 68576
rect 96440 68512 96456 68576
rect 96520 68512 96536 68576
rect 96600 68512 96616 68576
rect 96680 68512 96688 68576
rect 96368 67488 96688 68512
rect 96368 67424 96376 67488
rect 96440 67424 96456 67488
rect 96520 67424 96536 67488
rect 96600 67424 96616 67488
rect 96680 67424 96688 67488
rect 96368 66400 96688 67424
rect 96368 66336 96376 66400
rect 96440 66336 96456 66400
rect 96520 66336 96536 66400
rect 96600 66336 96616 66400
rect 96680 66336 96688 66400
rect 96368 65312 96688 66336
rect 96368 65248 96376 65312
rect 96440 65248 96456 65312
rect 96520 65248 96536 65312
rect 96600 65248 96616 65312
rect 96680 65248 96688 65312
rect 96368 64224 96688 65248
rect 96368 64160 96376 64224
rect 96440 64160 96456 64224
rect 96520 64160 96536 64224
rect 96600 64160 96616 64224
rect 96680 64160 96688 64224
rect 96368 63136 96688 64160
rect 96368 63072 96376 63136
rect 96440 63072 96456 63136
rect 96520 63072 96536 63136
rect 96600 63072 96616 63136
rect 96680 63072 96688 63136
rect 96368 62048 96688 63072
rect 96368 61984 96376 62048
rect 96440 61984 96456 62048
rect 96520 61984 96536 62048
rect 96600 61984 96616 62048
rect 96680 61984 96688 62048
rect 96368 60960 96688 61984
rect 96368 60896 96376 60960
rect 96440 60896 96456 60960
rect 96520 60896 96536 60960
rect 96600 60896 96616 60960
rect 96680 60896 96688 60960
rect 96368 59872 96688 60896
rect 96368 59808 96376 59872
rect 96440 59808 96456 59872
rect 96520 59808 96536 59872
rect 96600 59808 96616 59872
rect 96680 59808 96688 59872
rect 96368 58784 96688 59808
rect 96368 58720 96376 58784
rect 96440 58720 96456 58784
rect 96520 58720 96536 58784
rect 96600 58720 96616 58784
rect 96680 58720 96688 58784
rect 96368 57696 96688 58720
rect 96368 57632 96376 57696
rect 96440 57632 96456 57696
rect 96520 57632 96536 57696
rect 96600 57632 96616 57696
rect 96680 57632 96688 57696
rect 96368 56608 96688 57632
rect 96368 56544 96376 56608
rect 96440 56544 96456 56608
rect 96520 56544 96536 56608
rect 96600 56544 96616 56608
rect 96680 56544 96688 56608
rect 96368 55520 96688 56544
rect 96368 55456 96376 55520
rect 96440 55456 96456 55520
rect 96520 55456 96536 55520
rect 96600 55456 96616 55520
rect 96680 55456 96688 55520
rect 96368 54432 96688 55456
rect 96368 54368 96376 54432
rect 96440 54368 96456 54432
rect 96520 54368 96536 54432
rect 96600 54368 96616 54432
rect 96680 54368 96688 54432
rect 96368 53344 96688 54368
rect 96368 53280 96376 53344
rect 96440 53280 96456 53344
rect 96520 53280 96536 53344
rect 96600 53280 96616 53344
rect 96680 53280 96688 53344
rect 96368 52256 96688 53280
rect 96368 52192 96376 52256
rect 96440 52192 96456 52256
rect 96520 52192 96536 52256
rect 96600 52192 96616 52256
rect 96680 52192 96688 52256
rect 96368 51168 96688 52192
rect 96368 51104 96376 51168
rect 96440 51104 96456 51168
rect 96520 51104 96536 51168
rect 96600 51104 96616 51168
rect 96680 51104 96688 51168
rect 96368 50080 96688 51104
rect 96368 50016 96376 50080
rect 96440 50016 96456 50080
rect 96520 50016 96536 50080
rect 96600 50016 96616 50080
rect 96680 50016 96688 50080
rect 96368 48992 96688 50016
rect 96368 48928 96376 48992
rect 96440 48928 96456 48992
rect 96520 48928 96536 48992
rect 96600 48928 96616 48992
rect 96680 48928 96688 48992
rect 96368 47904 96688 48928
rect 96368 47840 96376 47904
rect 96440 47840 96456 47904
rect 96520 47840 96536 47904
rect 96600 47840 96616 47904
rect 96680 47840 96688 47904
rect 96368 46816 96688 47840
rect 96368 46752 96376 46816
rect 96440 46752 96456 46816
rect 96520 46752 96536 46816
rect 96600 46752 96616 46816
rect 96680 46752 96688 46816
rect 96368 45728 96688 46752
rect 96368 45664 96376 45728
rect 96440 45664 96456 45728
rect 96520 45664 96536 45728
rect 96600 45664 96616 45728
rect 96680 45664 96688 45728
rect 96368 44640 96688 45664
rect 96368 44576 96376 44640
rect 96440 44576 96456 44640
rect 96520 44576 96536 44640
rect 96600 44576 96616 44640
rect 96680 44576 96688 44640
rect 96368 43552 96688 44576
rect 96368 43488 96376 43552
rect 96440 43488 96456 43552
rect 96520 43488 96536 43552
rect 96600 43488 96616 43552
rect 96680 43488 96688 43552
rect 96368 42464 96688 43488
rect 96368 42400 96376 42464
rect 96440 42400 96456 42464
rect 96520 42400 96536 42464
rect 96600 42400 96616 42464
rect 96680 42400 96688 42464
rect 96368 41376 96688 42400
rect 96368 41312 96376 41376
rect 96440 41312 96456 41376
rect 96520 41312 96536 41376
rect 96600 41312 96616 41376
rect 96680 41312 96688 41376
rect 96368 40288 96688 41312
rect 96368 40224 96376 40288
rect 96440 40224 96456 40288
rect 96520 40224 96536 40288
rect 96600 40224 96616 40288
rect 96680 40224 96688 40288
rect 96368 39200 96688 40224
rect 96368 39136 96376 39200
rect 96440 39136 96456 39200
rect 96520 39136 96536 39200
rect 96600 39136 96616 39200
rect 96680 39136 96688 39200
rect 96368 38112 96688 39136
rect 96368 38048 96376 38112
rect 96440 38048 96456 38112
rect 96520 38048 96536 38112
rect 96600 38048 96616 38112
rect 96680 38048 96688 38112
rect 96368 37024 96688 38048
rect 96368 36960 96376 37024
rect 96440 36960 96456 37024
rect 96520 36960 96536 37024
rect 96600 36960 96616 37024
rect 96680 36960 96688 37024
rect 96368 35936 96688 36960
rect 96368 35872 96376 35936
rect 96440 35872 96456 35936
rect 96520 35872 96536 35936
rect 96600 35872 96616 35936
rect 96680 35872 96688 35936
rect 96368 34848 96688 35872
rect 96368 34784 96376 34848
rect 96440 34784 96456 34848
rect 96520 34784 96536 34848
rect 96600 34784 96616 34848
rect 96680 34784 96688 34848
rect 96368 33760 96688 34784
rect 96368 33696 96376 33760
rect 96440 33696 96456 33760
rect 96520 33696 96536 33760
rect 96600 33696 96616 33760
rect 96680 33696 96688 33760
rect 96368 32672 96688 33696
rect 96368 32608 96376 32672
rect 96440 32608 96456 32672
rect 96520 32608 96536 32672
rect 96600 32608 96616 32672
rect 96680 32608 96688 32672
rect 96368 31584 96688 32608
rect 96368 31520 96376 31584
rect 96440 31520 96456 31584
rect 96520 31520 96536 31584
rect 96600 31520 96616 31584
rect 96680 31520 96688 31584
rect 96368 30496 96688 31520
rect 96368 30432 96376 30496
rect 96440 30432 96456 30496
rect 96520 30432 96536 30496
rect 96600 30432 96616 30496
rect 96680 30432 96688 30496
rect 96368 29408 96688 30432
rect 96368 29344 96376 29408
rect 96440 29344 96456 29408
rect 96520 29344 96536 29408
rect 96600 29344 96616 29408
rect 96680 29344 96688 29408
rect 96368 28320 96688 29344
rect 96368 28256 96376 28320
rect 96440 28256 96456 28320
rect 96520 28256 96536 28320
rect 96600 28256 96616 28320
rect 96680 28256 96688 28320
rect 96368 27232 96688 28256
rect 96368 27168 96376 27232
rect 96440 27168 96456 27232
rect 96520 27168 96536 27232
rect 96600 27168 96616 27232
rect 96680 27168 96688 27232
rect 96368 26144 96688 27168
rect 96368 26080 96376 26144
rect 96440 26080 96456 26144
rect 96520 26080 96536 26144
rect 96600 26080 96616 26144
rect 96680 26080 96688 26144
rect 96368 25056 96688 26080
rect 96368 24992 96376 25056
rect 96440 24992 96456 25056
rect 96520 24992 96536 25056
rect 96600 24992 96616 25056
rect 96680 24992 96688 25056
rect 96368 23968 96688 24992
rect 96368 23904 96376 23968
rect 96440 23904 96456 23968
rect 96520 23904 96536 23968
rect 96600 23904 96616 23968
rect 96680 23904 96688 23968
rect 96368 22880 96688 23904
rect 96368 22816 96376 22880
rect 96440 22816 96456 22880
rect 96520 22816 96536 22880
rect 96600 22816 96616 22880
rect 96680 22816 96688 22880
rect 96368 21792 96688 22816
rect 96368 21728 96376 21792
rect 96440 21728 96456 21792
rect 96520 21728 96536 21792
rect 96600 21728 96616 21792
rect 96680 21728 96688 21792
rect 96368 20704 96688 21728
rect 96368 20640 96376 20704
rect 96440 20640 96456 20704
rect 96520 20640 96536 20704
rect 96600 20640 96616 20704
rect 96680 20640 96688 20704
rect 96368 19616 96688 20640
rect 96368 19552 96376 19616
rect 96440 19552 96456 19616
rect 96520 19552 96536 19616
rect 96600 19552 96616 19616
rect 96680 19552 96688 19616
rect 96368 18528 96688 19552
rect 96368 18464 96376 18528
rect 96440 18464 96456 18528
rect 96520 18464 96536 18528
rect 96600 18464 96616 18528
rect 96680 18464 96688 18528
rect 96368 17440 96688 18464
rect 96368 17376 96376 17440
rect 96440 17376 96456 17440
rect 96520 17376 96536 17440
rect 96600 17376 96616 17440
rect 96680 17376 96688 17440
rect 96368 16352 96688 17376
rect 96368 16288 96376 16352
rect 96440 16288 96456 16352
rect 96520 16288 96536 16352
rect 96600 16288 96616 16352
rect 96680 16288 96688 16352
rect 96368 15264 96688 16288
rect 96368 15200 96376 15264
rect 96440 15200 96456 15264
rect 96520 15200 96536 15264
rect 96600 15200 96616 15264
rect 96680 15200 96688 15264
rect 96368 14176 96688 15200
rect 96368 14112 96376 14176
rect 96440 14112 96456 14176
rect 96520 14112 96536 14176
rect 96600 14112 96616 14176
rect 96680 14112 96688 14176
rect 96368 13088 96688 14112
rect 96368 13024 96376 13088
rect 96440 13024 96456 13088
rect 96520 13024 96536 13088
rect 96600 13024 96616 13088
rect 96680 13024 96688 13088
rect 96368 12000 96688 13024
rect 96368 11936 96376 12000
rect 96440 11936 96456 12000
rect 96520 11936 96536 12000
rect 96600 11936 96616 12000
rect 96680 11936 96688 12000
rect 96368 10912 96688 11936
rect 96368 10848 96376 10912
rect 96440 10848 96456 10912
rect 96520 10848 96536 10912
rect 96600 10848 96616 10912
rect 96680 10848 96688 10912
rect 96368 9824 96688 10848
rect 96368 9760 96376 9824
rect 96440 9760 96456 9824
rect 96520 9760 96536 9824
rect 96600 9760 96616 9824
rect 96680 9760 96688 9824
rect 96368 8736 96688 9760
rect 96368 8672 96376 8736
rect 96440 8672 96456 8736
rect 96520 8672 96536 8736
rect 96600 8672 96616 8736
rect 96680 8672 96688 8736
rect 96368 7648 96688 8672
rect 96368 7584 96376 7648
rect 96440 7584 96456 7648
rect 96520 7584 96536 7648
rect 96600 7584 96616 7648
rect 96680 7584 96688 7648
rect 96368 6560 96688 7584
rect 96368 6496 96376 6560
rect 96440 6496 96456 6560
rect 96520 6496 96536 6560
rect 96600 6496 96616 6560
rect 96680 6496 96688 6560
rect 96368 5472 96688 6496
rect 96368 5408 96376 5472
rect 96440 5408 96456 5472
rect 96520 5408 96536 5472
rect 96600 5408 96616 5472
rect 96680 5408 96688 5472
rect 96368 4384 96688 5408
rect 96368 4320 96376 4384
rect 96440 4320 96456 4384
rect 96520 4320 96536 4384
rect 96600 4320 96616 4384
rect 96680 4320 96688 4384
rect 86539 4316 86605 4317
rect 86539 4252 86540 4316
rect 86604 4252 86605 4316
rect 86539 4251 86605 4252
rect 86171 3500 86237 3501
rect 86171 3436 86172 3500
rect 86236 3436 86237 3500
rect 86171 3435 86237 3436
rect 86174 2821 86234 3435
rect 86542 2821 86602 4251
rect 86723 4044 86789 4045
rect 86723 3980 86724 4044
rect 86788 3980 86789 4044
rect 86723 3979 86789 3980
rect 86171 2820 86237 2821
rect 86171 2756 86172 2820
rect 86236 2756 86237 2820
rect 86171 2755 86237 2756
rect 86539 2820 86605 2821
rect 86539 2756 86540 2820
rect 86604 2756 86605 2820
rect 86539 2755 86605 2756
rect 86726 2005 86786 3979
rect 88379 3772 88445 3773
rect 88379 3708 88380 3772
rect 88444 3708 88445 3772
rect 88379 3707 88445 3708
rect 89670 3710 89914 3770
rect 88382 3634 88442 3707
rect 89670 3637 89730 3710
rect 89854 3637 89914 3710
rect 88747 3636 88813 3637
rect 88747 3634 88748 3636
rect 88382 3574 88748 3634
rect 88747 3572 88748 3574
rect 88812 3572 88813 3636
rect 88747 3571 88813 3572
rect 89667 3636 89733 3637
rect 89667 3572 89668 3636
rect 89732 3572 89733 3636
rect 89667 3571 89733 3572
rect 89851 3636 89917 3637
rect 89851 3572 89852 3636
rect 89916 3572 89917 3636
rect 89851 3571 89917 3572
rect 96368 3296 96688 4320
rect 96368 3232 96376 3296
rect 96440 3232 96456 3296
rect 96520 3232 96536 3296
rect 96600 3232 96616 3296
rect 96680 3232 96688 3296
rect 96368 2208 96688 3232
rect 96368 2144 96376 2208
rect 96440 2144 96456 2208
rect 96520 2144 96536 2208
rect 96600 2144 96616 2208
rect 96680 2144 96688 2208
rect 97028 2176 97348 117504
rect 97688 2176 98008 117504
rect 98348 2176 98668 117504
rect 111728 116992 112048 117552
rect 127088 117536 127408 117552
rect 111728 116928 111736 116992
rect 111800 116928 111816 116992
rect 111880 116928 111896 116992
rect 111960 116928 111976 116992
rect 112040 116928 112048 116992
rect 111728 115904 112048 116928
rect 111728 115840 111736 115904
rect 111800 115840 111816 115904
rect 111880 115840 111896 115904
rect 111960 115840 111976 115904
rect 112040 115840 112048 115904
rect 111728 114816 112048 115840
rect 111728 114752 111736 114816
rect 111800 114752 111816 114816
rect 111880 114752 111896 114816
rect 111960 114752 111976 114816
rect 112040 114752 112048 114816
rect 111728 113728 112048 114752
rect 111728 113664 111736 113728
rect 111800 113664 111816 113728
rect 111880 113664 111896 113728
rect 111960 113664 111976 113728
rect 112040 113664 112048 113728
rect 111728 112640 112048 113664
rect 111728 112576 111736 112640
rect 111800 112576 111816 112640
rect 111880 112576 111896 112640
rect 111960 112576 111976 112640
rect 112040 112576 112048 112640
rect 111728 111552 112048 112576
rect 111728 111488 111736 111552
rect 111800 111488 111816 111552
rect 111880 111488 111896 111552
rect 111960 111488 111976 111552
rect 112040 111488 112048 111552
rect 111728 110464 112048 111488
rect 111728 110400 111736 110464
rect 111800 110400 111816 110464
rect 111880 110400 111896 110464
rect 111960 110400 111976 110464
rect 112040 110400 112048 110464
rect 111728 109376 112048 110400
rect 111728 109312 111736 109376
rect 111800 109312 111816 109376
rect 111880 109312 111896 109376
rect 111960 109312 111976 109376
rect 112040 109312 112048 109376
rect 111728 108288 112048 109312
rect 111728 108224 111736 108288
rect 111800 108224 111816 108288
rect 111880 108224 111896 108288
rect 111960 108224 111976 108288
rect 112040 108224 112048 108288
rect 111728 107200 112048 108224
rect 111728 107136 111736 107200
rect 111800 107136 111816 107200
rect 111880 107136 111896 107200
rect 111960 107136 111976 107200
rect 112040 107136 112048 107200
rect 111728 106112 112048 107136
rect 111728 106048 111736 106112
rect 111800 106048 111816 106112
rect 111880 106048 111896 106112
rect 111960 106048 111976 106112
rect 112040 106048 112048 106112
rect 111728 105024 112048 106048
rect 111728 104960 111736 105024
rect 111800 104960 111816 105024
rect 111880 104960 111896 105024
rect 111960 104960 111976 105024
rect 112040 104960 112048 105024
rect 111728 103936 112048 104960
rect 111728 103872 111736 103936
rect 111800 103872 111816 103936
rect 111880 103872 111896 103936
rect 111960 103872 111976 103936
rect 112040 103872 112048 103936
rect 111728 102848 112048 103872
rect 111728 102784 111736 102848
rect 111800 102784 111816 102848
rect 111880 102784 111896 102848
rect 111960 102784 111976 102848
rect 112040 102784 112048 102848
rect 111728 101760 112048 102784
rect 111728 101696 111736 101760
rect 111800 101696 111816 101760
rect 111880 101696 111896 101760
rect 111960 101696 111976 101760
rect 112040 101696 112048 101760
rect 111728 100672 112048 101696
rect 111728 100608 111736 100672
rect 111800 100608 111816 100672
rect 111880 100608 111896 100672
rect 111960 100608 111976 100672
rect 112040 100608 112048 100672
rect 111728 99584 112048 100608
rect 111728 99520 111736 99584
rect 111800 99520 111816 99584
rect 111880 99520 111896 99584
rect 111960 99520 111976 99584
rect 112040 99520 112048 99584
rect 111728 98496 112048 99520
rect 111728 98432 111736 98496
rect 111800 98432 111816 98496
rect 111880 98432 111896 98496
rect 111960 98432 111976 98496
rect 112040 98432 112048 98496
rect 111728 97408 112048 98432
rect 111728 97344 111736 97408
rect 111800 97344 111816 97408
rect 111880 97344 111896 97408
rect 111960 97344 111976 97408
rect 112040 97344 112048 97408
rect 111728 96320 112048 97344
rect 111728 96256 111736 96320
rect 111800 96256 111816 96320
rect 111880 96256 111896 96320
rect 111960 96256 111976 96320
rect 112040 96256 112048 96320
rect 111728 95232 112048 96256
rect 111728 95168 111736 95232
rect 111800 95168 111816 95232
rect 111880 95168 111896 95232
rect 111960 95168 111976 95232
rect 112040 95168 112048 95232
rect 111728 94144 112048 95168
rect 111728 94080 111736 94144
rect 111800 94080 111816 94144
rect 111880 94080 111896 94144
rect 111960 94080 111976 94144
rect 112040 94080 112048 94144
rect 111728 93056 112048 94080
rect 111728 92992 111736 93056
rect 111800 92992 111816 93056
rect 111880 92992 111896 93056
rect 111960 92992 111976 93056
rect 112040 92992 112048 93056
rect 111728 91968 112048 92992
rect 111728 91904 111736 91968
rect 111800 91904 111816 91968
rect 111880 91904 111896 91968
rect 111960 91904 111976 91968
rect 112040 91904 112048 91968
rect 111728 90880 112048 91904
rect 111728 90816 111736 90880
rect 111800 90816 111816 90880
rect 111880 90816 111896 90880
rect 111960 90816 111976 90880
rect 112040 90816 112048 90880
rect 111728 89792 112048 90816
rect 111728 89728 111736 89792
rect 111800 89728 111816 89792
rect 111880 89728 111896 89792
rect 111960 89728 111976 89792
rect 112040 89728 112048 89792
rect 111728 88704 112048 89728
rect 111728 88640 111736 88704
rect 111800 88640 111816 88704
rect 111880 88640 111896 88704
rect 111960 88640 111976 88704
rect 112040 88640 112048 88704
rect 111728 87616 112048 88640
rect 111728 87552 111736 87616
rect 111800 87552 111816 87616
rect 111880 87552 111896 87616
rect 111960 87552 111976 87616
rect 112040 87552 112048 87616
rect 111728 86528 112048 87552
rect 111728 86464 111736 86528
rect 111800 86464 111816 86528
rect 111880 86464 111896 86528
rect 111960 86464 111976 86528
rect 112040 86464 112048 86528
rect 111728 85440 112048 86464
rect 111728 85376 111736 85440
rect 111800 85376 111816 85440
rect 111880 85376 111896 85440
rect 111960 85376 111976 85440
rect 112040 85376 112048 85440
rect 111728 84352 112048 85376
rect 111728 84288 111736 84352
rect 111800 84288 111816 84352
rect 111880 84288 111896 84352
rect 111960 84288 111976 84352
rect 112040 84288 112048 84352
rect 111728 83264 112048 84288
rect 111728 83200 111736 83264
rect 111800 83200 111816 83264
rect 111880 83200 111896 83264
rect 111960 83200 111976 83264
rect 112040 83200 112048 83264
rect 111728 82176 112048 83200
rect 111728 82112 111736 82176
rect 111800 82112 111816 82176
rect 111880 82112 111896 82176
rect 111960 82112 111976 82176
rect 112040 82112 112048 82176
rect 111728 81088 112048 82112
rect 111728 81024 111736 81088
rect 111800 81024 111816 81088
rect 111880 81024 111896 81088
rect 111960 81024 111976 81088
rect 112040 81024 112048 81088
rect 111728 80000 112048 81024
rect 111728 79936 111736 80000
rect 111800 79936 111816 80000
rect 111880 79936 111896 80000
rect 111960 79936 111976 80000
rect 112040 79936 112048 80000
rect 111728 78912 112048 79936
rect 111728 78848 111736 78912
rect 111800 78848 111816 78912
rect 111880 78848 111896 78912
rect 111960 78848 111976 78912
rect 112040 78848 112048 78912
rect 111728 77824 112048 78848
rect 111728 77760 111736 77824
rect 111800 77760 111816 77824
rect 111880 77760 111896 77824
rect 111960 77760 111976 77824
rect 112040 77760 112048 77824
rect 111728 76736 112048 77760
rect 111728 76672 111736 76736
rect 111800 76672 111816 76736
rect 111880 76672 111896 76736
rect 111960 76672 111976 76736
rect 112040 76672 112048 76736
rect 111728 75648 112048 76672
rect 111728 75584 111736 75648
rect 111800 75584 111816 75648
rect 111880 75584 111896 75648
rect 111960 75584 111976 75648
rect 112040 75584 112048 75648
rect 111728 74560 112048 75584
rect 111728 74496 111736 74560
rect 111800 74496 111816 74560
rect 111880 74496 111896 74560
rect 111960 74496 111976 74560
rect 112040 74496 112048 74560
rect 111728 73472 112048 74496
rect 111728 73408 111736 73472
rect 111800 73408 111816 73472
rect 111880 73408 111896 73472
rect 111960 73408 111976 73472
rect 112040 73408 112048 73472
rect 111728 72384 112048 73408
rect 111728 72320 111736 72384
rect 111800 72320 111816 72384
rect 111880 72320 111896 72384
rect 111960 72320 111976 72384
rect 112040 72320 112048 72384
rect 111728 71296 112048 72320
rect 111728 71232 111736 71296
rect 111800 71232 111816 71296
rect 111880 71232 111896 71296
rect 111960 71232 111976 71296
rect 112040 71232 112048 71296
rect 111728 70208 112048 71232
rect 111728 70144 111736 70208
rect 111800 70144 111816 70208
rect 111880 70144 111896 70208
rect 111960 70144 111976 70208
rect 112040 70144 112048 70208
rect 111728 69120 112048 70144
rect 111728 69056 111736 69120
rect 111800 69056 111816 69120
rect 111880 69056 111896 69120
rect 111960 69056 111976 69120
rect 112040 69056 112048 69120
rect 111728 68032 112048 69056
rect 111728 67968 111736 68032
rect 111800 67968 111816 68032
rect 111880 67968 111896 68032
rect 111960 67968 111976 68032
rect 112040 67968 112048 68032
rect 111728 66944 112048 67968
rect 111728 66880 111736 66944
rect 111800 66880 111816 66944
rect 111880 66880 111896 66944
rect 111960 66880 111976 66944
rect 112040 66880 112048 66944
rect 111728 65856 112048 66880
rect 111728 65792 111736 65856
rect 111800 65792 111816 65856
rect 111880 65792 111896 65856
rect 111960 65792 111976 65856
rect 112040 65792 112048 65856
rect 111728 64768 112048 65792
rect 111728 64704 111736 64768
rect 111800 64704 111816 64768
rect 111880 64704 111896 64768
rect 111960 64704 111976 64768
rect 112040 64704 112048 64768
rect 111728 63680 112048 64704
rect 111728 63616 111736 63680
rect 111800 63616 111816 63680
rect 111880 63616 111896 63680
rect 111960 63616 111976 63680
rect 112040 63616 112048 63680
rect 111728 62592 112048 63616
rect 111728 62528 111736 62592
rect 111800 62528 111816 62592
rect 111880 62528 111896 62592
rect 111960 62528 111976 62592
rect 112040 62528 112048 62592
rect 111728 61504 112048 62528
rect 111728 61440 111736 61504
rect 111800 61440 111816 61504
rect 111880 61440 111896 61504
rect 111960 61440 111976 61504
rect 112040 61440 112048 61504
rect 111728 60416 112048 61440
rect 111728 60352 111736 60416
rect 111800 60352 111816 60416
rect 111880 60352 111896 60416
rect 111960 60352 111976 60416
rect 112040 60352 112048 60416
rect 111728 59328 112048 60352
rect 111728 59264 111736 59328
rect 111800 59264 111816 59328
rect 111880 59264 111896 59328
rect 111960 59264 111976 59328
rect 112040 59264 112048 59328
rect 111728 58240 112048 59264
rect 111728 58176 111736 58240
rect 111800 58176 111816 58240
rect 111880 58176 111896 58240
rect 111960 58176 111976 58240
rect 112040 58176 112048 58240
rect 111728 57152 112048 58176
rect 111728 57088 111736 57152
rect 111800 57088 111816 57152
rect 111880 57088 111896 57152
rect 111960 57088 111976 57152
rect 112040 57088 112048 57152
rect 111728 56064 112048 57088
rect 111728 56000 111736 56064
rect 111800 56000 111816 56064
rect 111880 56000 111896 56064
rect 111960 56000 111976 56064
rect 112040 56000 112048 56064
rect 111728 54976 112048 56000
rect 111728 54912 111736 54976
rect 111800 54912 111816 54976
rect 111880 54912 111896 54976
rect 111960 54912 111976 54976
rect 112040 54912 112048 54976
rect 111728 53888 112048 54912
rect 111728 53824 111736 53888
rect 111800 53824 111816 53888
rect 111880 53824 111896 53888
rect 111960 53824 111976 53888
rect 112040 53824 112048 53888
rect 111728 52800 112048 53824
rect 111728 52736 111736 52800
rect 111800 52736 111816 52800
rect 111880 52736 111896 52800
rect 111960 52736 111976 52800
rect 112040 52736 112048 52800
rect 111728 51712 112048 52736
rect 111728 51648 111736 51712
rect 111800 51648 111816 51712
rect 111880 51648 111896 51712
rect 111960 51648 111976 51712
rect 112040 51648 112048 51712
rect 111728 50624 112048 51648
rect 111728 50560 111736 50624
rect 111800 50560 111816 50624
rect 111880 50560 111896 50624
rect 111960 50560 111976 50624
rect 112040 50560 112048 50624
rect 111728 49536 112048 50560
rect 111728 49472 111736 49536
rect 111800 49472 111816 49536
rect 111880 49472 111896 49536
rect 111960 49472 111976 49536
rect 112040 49472 112048 49536
rect 111728 48448 112048 49472
rect 111728 48384 111736 48448
rect 111800 48384 111816 48448
rect 111880 48384 111896 48448
rect 111960 48384 111976 48448
rect 112040 48384 112048 48448
rect 111728 47360 112048 48384
rect 111728 47296 111736 47360
rect 111800 47296 111816 47360
rect 111880 47296 111896 47360
rect 111960 47296 111976 47360
rect 112040 47296 112048 47360
rect 111728 46272 112048 47296
rect 111728 46208 111736 46272
rect 111800 46208 111816 46272
rect 111880 46208 111896 46272
rect 111960 46208 111976 46272
rect 112040 46208 112048 46272
rect 111728 45184 112048 46208
rect 111728 45120 111736 45184
rect 111800 45120 111816 45184
rect 111880 45120 111896 45184
rect 111960 45120 111976 45184
rect 112040 45120 112048 45184
rect 111728 44096 112048 45120
rect 111728 44032 111736 44096
rect 111800 44032 111816 44096
rect 111880 44032 111896 44096
rect 111960 44032 111976 44096
rect 112040 44032 112048 44096
rect 111728 43008 112048 44032
rect 111728 42944 111736 43008
rect 111800 42944 111816 43008
rect 111880 42944 111896 43008
rect 111960 42944 111976 43008
rect 112040 42944 112048 43008
rect 111728 41920 112048 42944
rect 111728 41856 111736 41920
rect 111800 41856 111816 41920
rect 111880 41856 111896 41920
rect 111960 41856 111976 41920
rect 112040 41856 112048 41920
rect 111728 40832 112048 41856
rect 111728 40768 111736 40832
rect 111800 40768 111816 40832
rect 111880 40768 111896 40832
rect 111960 40768 111976 40832
rect 112040 40768 112048 40832
rect 111728 39744 112048 40768
rect 111728 39680 111736 39744
rect 111800 39680 111816 39744
rect 111880 39680 111896 39744
rect 111960 39680 111976 39744
rect 112040 39680 112048 39744
rect 111728 38656 112048 39680
rect 111728 38592 111736 38656
rect 111800 38592 111816 38656
rect 111880 38592 111896 38656
rect 111960 38592 111976 38656
rect 112040 38592 112048 38656
rect 111728 37568 112048 38592
rect 111728 37504 111736 37568
rect 111800 37504 111816 37568
rect 111880 37504 111896 37568
rect 111960 37504 111976 37568
rect 112040 37504 112048 37568
rect 111728 36480 112048 37504
rect 111728 36416 111736 36480
rect 111800 36416 111816 36480
rect 111880 36416 111896 36480
rect 111960 36416 111976 36480
rect 112040 36416 112048 36480
rect 111728 35392 112048 36416
rect 111728 35328 111736 35392
rect 111800 35328 111816 35392
rect 111880 35328 111896 35392
rect 111960 35328 111976 35392
rect 112040 35328 112048 35392
rect 111728 34304 112048 35328
rect 111728 34240 111736 34304
rect 111800 34240 111816 34304
rect 111880 34240 111896 34304
rect 111960 34240 111976 34304
rect 112040 34240 112048 34304
rect 111728 33216 112048 34240
rect 111728 33152 111736 33216
rect 111800 33152 111816 33216
rect 111880 33152 111896 33216
rect 111960 33152 111976 33216
rect 112040 33152 112048 33216
rect 111728 32128 112048 33152
rect 111728 32064 111736 32128
rect 111800 32064 111816 32128
rect 111880 32064 111896 32128
rect 111960 32064 111976 32128
rect 112040 32064 112048 32128
rect 111728 31040 112048 32064
rect 111728 30976 111736 31040
rect 111800 30976 111816 31040
rect 111880 30976 111896 31040
rect 111960 30976 111976 31040
rect 112040 30976 112048 31040
rect 111728 29952 112048 30976
rect 111728 29888 111736 29952
rect 111800 29888 111816 29952
rect 111880 29888 111896 29952
rect 111960 29888 111976 29952
rect 112040 29888 112048 29952
rect 111728 28864 112048 29888
rect 111728 28800 111736 28864
rect 111800 28800 111816 28864
rect 111880 28800 111896 28864
rect 111960 28800 111976 28864
rect 112040 28800 112048 28864
rect 111728 27776 112048 28800
rect 111728 27712 111736 27776
rect 111800 27712 111816 27776
rect 111880 27712 111896 27776
rect 111960 27712 111976 27776
rect 112040 27712 112048 27776
rect 111728 26688 112048 27712
rect 111728 26624 111736 26688
rect 111800 26624 111816 26688
rect 111880 26624 111896 26688
rect 111960 26624 111976 26688
rect 112040 26624 112048 26688
rect 111728 25600 112048 26624
rect 111728 25536 111736 25600
rect 111800 25536 111816 25600
rect 111880 25536 111896 25600
rect 111960 25536 111976 25600
rect 112040 25536 112048 25600
rect 111728 24512 112048 25536
rect 111728 24448 111736 24512
rect 111800 24448 111816 24512
rect 111880 24448 111896 24512
rect 111960 24448 111976 24512
rect 112040 24448 112048 24512
rect 111728 23424 112048 24448
rect 111728 23360 111736 23424
rect 111800 23360 111816 23424
rect 111880 23360 111896 23424
rect 111960 23360 111976 23424
rect 112040 23360 112048 23424
rect 111728 22336 112048 23360
rect 111728 22272 111736 22336
rect 111800 22272 111816 22336
rect 111880 22272 111896 22336
rect 111960 22272 111976 22336
rect 112040 22272 112048 22336
rect 111728 21248 112048 22272
rect 111728 21184 111736 21248
rect 111800 21184 111816 21248
rect 111880 21184 111896 21248
rect 111960 21184 111976 21248
rect 112040 21184 112048 21248
rect 111728 20160 112048 21184
rect 111728 20096 111736 20160
rect 111800 20096 111816 20160
rect 111880 20096 111896 20160
rect 111960 20096 111976 20160
rect 112040 20096 112048 20160
rect 111728 19072 112048 20096
rect 111728 19008 111736 19072
rect 111800 19008 111816 19072
rect 111880 19008 111896 19072
rect 111960 19008 111976 19072
rect 112040 19008 112048 19072
rect 111728 17984 112048 19008
rect 111728 17920 111736 17984
rect 111800 17920 111816 17984
rect 111880 17920 111896 17984
rect 111960 17920 111976 17984
rect 112040 17920 112048 17984
rect 111728 16896 112048 17920
rect 111728 16832 111736 16896
rect 111800 16832 111816 16896
rect 111880 16832 111896 16896
rect 111960 16832 111976 16896
rect 112040 16832 112048 16896
rect 111728 15808 112048 16832
rect 111728 15744 111736 15808
rect 111800 15744 111816 15808
rect 111880 15744 111896 15808
rect 111960 15744 111976 15808
rect 112040 15744 112048 15808
rect 111728 14720 112048 15744
rect 111728 14656 111736 14720
rect 111800 14656 111816 14720
rect 111880 14656 111896 14720
rect 111960 14656 111976 14720
rect 112040 14656 112048 14720
rect 111728 13632 112048 14656
rect 111728 13568 111736 13632
rect 111800 13568 111816 13632
rect 111880 13568 111896 13632
rect 111960 13568 111976 13632
rect 112040 13568 112048 13632
rect 111728 12544 112048 13568
rect 111728 12480 111736 12544
rect 111800 12480 111816 12544
rect 111880 12480 111896 12544
rect 111960 12480 111976 12544
rect 112040 12480 112048 12544
rect 111728 11456 112048 12480
rect 111728 11392 111736 11456
rect 111800 11392 111816 11456
rect 111880 11392 111896 11456
rect 111960 11392 111976 11456
rect 112040 11392 112048 11456
rect 111728 10368 112048 11392
rect 111728 10304 111736 10368
rect 111800 10304 111816 10368
rect 111880 10304 111896 10368
rect 111960 10304 111976 10368
rect 112040 10304 112048 10368
rect 111728 9280 112048 10304
rect 111728 9216 111736 9280
rect 111800 9216 111816 9280
rect 111880 9216 111896 9280
rect 111960 9216 111976 9280
rect 112040 9216 112048 9280
rect 111728 8192 112048 9216
rect 111728 8128 111736 8192
rect 111800 8128 111816 8192
rect 111880 8128 111896 8192
rect 111960 8128 111976 8192
rect 112040 8128 112048 8192
rect 111728 7104 112048 8128
rect 111728 7040 111736 7104
rect 111800 7040 111816 7104
rect 111880 7040 111896 7104
rect 111960 7040 111976 7104
rect 112040 7040 112048 7104
rect 111728 6016 112048 7040
rect 111728 5952 111736 6016
rect 111800 5952 111816 6016
rect 111880 5952 111896 6016
rect 111960 5952 111976 6016
rect 112040 5952 112048 6016
rect 111728 4928 112048 5952
rect 111728 4864 111736 4928
rect 111800 4864 111816 4928
rect 111880 4864 111896 4928
rect 111960 4864 111976 4928
rect 112040 4864 112048 4928
rect 111728 3840 112048 4864
rect 111728 3776 111736 3840
rect 111800 3776 111816 3840
rect 111880 3776 111896 3840
rect 111960 3776 111976 3840
rect 112040 3776 112048 3840
rect 111728 2752 112048 3776
rect 111728 2688 111736 2752
rect 111800 2688 111816 2752
rect 111880 2688 111896 2752
rect 111960 2688 111976 2752
rect 112040 2688 112048 2752
rect 96368 2128 96688 2144
rect 111728 2128 112048 2688
rect 112388 2176 112708 117504
rect 113048 2176 113368 117504
rect 113708 2176 114028 117504
rect 127088 117472 127096 117536
rect 127160 117472 127176 117536
rect 127240 117472 127256 117536
rect 127320 117472 127336 117536
rect 127400 117472 127408 117536
rect 127088 116448 127408 117472
rect 127088 116384 127096 116448
rect 127160 116384 127176 116448
rect 127240 116384 127256 116448
rect 127320 116384 127336 116448
rect 127400 116384 127408 116448
rect 127088 115360 127408 116384
rect 127088 115296 127096 115360
rect 127160 115296 127176 115360
rect 127240 115296 127256 115360
rect 127320 115296 127336 115360
rect 127400 115296 127408 115360
rect 127088 114272 127408 115296
rect 127088 114208 127096 114272
rect 127160 114208 127176 114272
rect 127240 114208 127256 114272
rect 127320 114208 127336 114272
rect 127400 114208 127408 114272
rect 127088 113184 127408 114208
rect 127088 113120 127096 113184
rect 127160 113120 127176 113184
rect 127240 113120 127256 113184
rect 127320 113120 127336 113184
rect 127400 113120 127408 113184
rect 127088 112096 127408 113120
rect 127088 112032 127096 112096
rect 127160 112032 127176 112096
rect 127240 112032 127256 112096
rect 127320 112032 127336 112096
rect 127400 112032 127408 112096
rect 127088 111008 127408 112032
rect 127088 110944 127096 111008
rect 127160 110944 127176 111008
rect 127240 110944 127256 111008
rect 127320 110944 127336 111008
rect 127400 110944 127408 111008
rect 127088 109920 127408 110944
rect 127088 109856 127096 109920
rect 127160 109856 127176 109920
rect 127240 109856 127256 109920
rect 127320 109856 127336 109920
rect 127400 109856 127408 109920
rect 127088 108832 127408 109856
rect 127088 108768 127096 108832
rect 127160 108768 127176 108832
rect 127240 108768 127256 108832
rect 127320 108768 127336 108832
rect 127400 108768 127408 108832
rect 127088 107744 127408 108768
rect 127088 107680 127096 107744
rect 127160 107680 127176 107744
rect 127240 107680 127256 107744
rect 127320 107680 127336 107744
rect 127400 107680 127408 107744
rect 127088 106656 127408 107680
rect 127088 106592 127096 106656
rect 127160 106592 127176 106656
rect 127240 106592 127256 106656
rect 127320 106592 127336 106656
rect 127400 106592 127408 106656
rect 127088 105568 127408 106592
rect 127088 105504 127096 105568
rect 127160 105504 127176 105568
rect 127240 105504 127256 105568
rect 127320 105504 127336 105568
rect 127400 105504 127408 105568
rect 127088 104480 127408 105504
rect 127088 104416 127096 104480
rect 127160 104416 127176 104480
rect 127240 104416 127256 104480
rect 127320 104416 127336 104480
rect 127400 104416 127408 104480
rect 127088 103392 127408 104416
rect 127088 103328 127096 103392
rect 127160 103328 127176 103392
rect 127240 103328 127256 103392
rect 127320 103328 127336 103392
rect 127400 103328 127408 103392
rect 127088 102304 127408 103328
rect 127088 102240 127096 102304
rect 127160 102240 127176 102304
rect 127240 102240 127256 102304
rect 127320 102240 127336 102304
rect 127400 102240 127408 102304
rect 127088 101216 127408 102240
rect 127088 101152 127096 101216
rect 127160 101152 127176 101216
rect 127240 101152 127256 101216
rect 127320 101152 127336 101216
rect 127400 101152 127408 101216
rect 127088 100128 127408 101152
rect 127088 100064 127096 100128
rect 127160 100064 127176 100128
rect 127240 100064 127256 100128
rect 127320 100064 127336 100128
rect 127400 100064 127408 100128
rect 127088 99040 127408 100064
rect 127088 98976 127096 99040
rect 127160 98976 127176 99040
rect 127240 98976 127256 99040
rect 127320 98976 127336 99040
rect 127400 98976 127408 99040
rect 127088 97952 127408 98976
rect 127088 97888 127096 97952
rect 127160 97888 127176 97952
rect 127240 97888 127256 97952
rect 127320 97888 127336 97952
rect 127400 97888 127408 97952
rect 127088 96864 127408 97888
rect 127088 96800 127096 96864
rect 127160 96800 127176 96864
rect 127240 96800 127256 96864
rect 127320 96800 127336 96864
rect 127400 96800 127408 96864
rect 127088 95776 127408 96800
rect 127088 95712 127096 95776
rect 127160 95712 127176 95776
rect 127240 95712 127256 95776
rect 127320 95712 127336 95776
rect 127400 95712 127408 95776
rect 127088 94688 127408 95712
rect 127088 94624 127096 94688
rect 127160 94624 127176 94688
rect 127240 94624 127256 94688
rect 127320 94624 127336 94688
rect 127400 94624 127408 94688
rect 127088 93600 127408 94624
rect 127088 93536 127096 93600
rect 127160 93536 127176 93600
rect 127240 93536 127256 93600
rect 127320 93536 127336 93600
rect 127400 93536 127408 93600
rect 127088 92512 127408 93536
rect 127088 92448 127096 92512
rect 127160 92448 127176 92512
rect 127240 92448 127256 92512
rect 127320 92448 127336 92512
rect 127400 92448 127408 92512
rect 127088 91424 127408 92448
rect 127088 91360 127096 91424
rect 127160 91360 127176 91424
rect 127240 91360 127256 91424
rect 127320 91360 127336 91424
rect 127400 91360 127408 91424
rect 127088 90336 127408 91360
rect 127088 90272 127096 90336
rect 127160 90272 127176 90336
rect 127240 90272 127256 90336
rect 127320 90272 127336 90336
rect 127400 90272 127408 90336
rect 127088 89248 127408 90272
rect 127088 89184 127096 89248
rect 127160 89184 127176 89248
rect 127240 89184 127256 89248
rect 127320 89184 127336 89248
rect 127400 89184 127408 89248
rect 127088 88160 127408 89184
rect 127088 88096 127096 88160
rect 127160 88096 127176 88160
rect 127240 88096 127256 88160
rect 127320 88096 127336 88160
rect 127400 88096 127408 88160
rect 127088 87072 127408 88096
rect 127088 87008 127096 87072
rect 127160 87008 127176 87072
rect 127240 87008 127256 87072
rect 127320 87008 127336 87072
rect 127400 87008 127408 87072
rect 127088 85984 127408 87008
rect 127088 85920 127096 85984
rect 127160 85920 127176 85984
rect 127240 85920 127256 85984
rect 127320 85920 127336 85984
rect 127400 85920 127408 85984
rect 127088 84896 127408 85920
rect 127088 84832 127096 84896
rect 127160 84832 127176 84896
rect 127240 84832 127256 84896
rect 127320 84832 127336 84896
rect 127400 84832 127408 84896
rect 127088 83808 127408 84832
rect 127088 83744 127096 83808
rect 127160 83744 127176 83808
rect 127240 83744 127256 83808
rect 127320 83744 127336 83808
rect 127400 83744 127408 83808
rect 127088 82720 127408 83744
rect 127088 82656 127096 82720
rect 127160 82656 127176 82720
rect 127240 82656 127256 82720
rect 127320 82656 127336 82720
rect 127400 82656 127408 82720
rect 127088 81632 127408 82656
rect 127088 81568 127096 81632
rect 127160 81568 127176 81632
rect 127240 81568 127256 81632
rect 127320 81568 127336 81632
rect 127400 81568 127408 81632
rect 127088 80544 127408 81568
rect 127088 80480 127096 80544
rect 127160 80480 127176 80544
rect 127240 80480 127256 80544
rect 127320 80480 127336 80544
rect 127400 80480 127408 80544
rect 127088 79456 127408 80480
rect 127088 79392 127096 79456
rect 127160 79392 127176 79456
rect 127240 79392 127256 79456
rect 127320 79392 127336 79456
rect 127400 79392 127408 79456
rect 127088 78368 127408 79392
rect 127088 78304 127096 78368
rect 127160 78304 127176 78368
rect 127240 78304 127256 78368
rect 127320 78304 127336 78368
rect 127400 78304 127408 78368
rect 127088 77280 127408 78304
rect 127088 77216 127096 77280
rect 127160 77216 127176 77280
rect 127240 77216 127256 77280
rect 127320 77216 127336 77280
rect 127400 77216 127408 77280
rect 127088 76192 127408 77216
rect 127088 76128 127096 76192
rect 127160 76128 127176 76192
rect 127240 76128 127256 76192
rect 127320 76128 127336 76192
rect 127400 76128 127408 76192
rect 127088 75104 127408 76128
rect 127088 75040 127096 75104
rect 127160 75040 127176 75104
rect 127240 75040 127256 75104
rect 127320 75040 127336 75104
rect 127400 75040 127408 75104
rect 127088 74016 127408 75040
rect 127088 73952 127096 74016
rect 127160 73952 127176 74016
rect 127240 73952 127256 74016
rect 127320 73952 127336 74016
rect 127400 73952 127408 74016
rect 127088 72928 127408 73952
rect 127088 72864 127096 72928
rect 127160 72864 127176 72928
rect 127240 72864 127256 72928
rect 127320 72864 127336 72928
rect 127400 72864 127408 72928
rect 127088 71840 127408 72864
rect 127088 71776 127096 71840
rect 127160 71776 127176 71840
rect 127240 71776 127256 71840
rect 127320 71776 127336 71840
rect 127400 71776 127408 71840
rect 127088 70752 127408 71776
rect 127088 70688 127096 70752
rect 127160 70688 127176 70752
rect 127240 70688 127256 70752
rect 127320 70688 127336 70752
rect 127400 70688 127408 70752
rect 127088 69664 127408 70688
rect 127088 69600 127096 69664
rect 127160 69600 127176 69664
rect 127240 69600 127256 69664
rect 127320 69600 127336 69664
rect 127400 69600 127408 69664
rect 127088 68576 127408 69600
rect 127088 68512 127096 68576
rect 127160 68512 127176 68576
rect 127240 68512 127256 68576
rect 127320 68512 127336 68576
rect 127400 68512 127408 68576
rect 127088 67488 127408 68512
rect 127088 67424 127096 67488
rect 127160 67424 127176 67488
rect 127240 67424 127256 67488
rect 127320 67424 127336 67488
rect 127400 67424 127408 67488
rect 127088 66400 127408 67424
rect 127088 66336 127096 66400
rect 127160 66336 127176 66400
rect 127240 66336 127256 66400
rect 127320 66336 127336 66400
rect 127400 66336 127408 66400
rect 127088 65312 127408 66336
rect 127088 65248 127096 65312
rect 127160 65248 127176 65312
rect 127240 65248 127256 65312
rect 127320 65248 127336 65312
rect 127400 65248 127408 65312
rect 127088 64224 127408 65248
rect 127088 64160 127096 64224
rect 127160 64160 127176 64224
rect 127240 64160 127256 64224
rect 127320 64160 127336 64224
rect 127400 64160 127408 64224
rect 127088 63136 127408 64160
rect 127088 63072 127096 63136
rect 127160 63072 127176 63136
rect 127240 63072 127256 63136
rect 127320 63072 127336 63136
rect 127400 63072 127408 63136
rect 127088 62048 127408 63072
rect 127088 61984 127096 62048
rect 127160 61984 127176 62048
rect 127240 61984 127256 62048
rect 127320 61984 127336 62048
rect 127400 61984 127408 62048
rect 127088 60960 127408 61984
rect 127088 60896 127096 60960
rect 127160 60896 127176 60960
rect 127240 60896 127256 60960
rect 127320 60896 127336 60960
rect 127400 60896 127408 60960
rect 127088 59872 127408 60896
rect 127088 59808 127096 59872
rect 127160 59808 127176 59872
rect 127240 59808 127256 59872
rect 127320 59808 127336 59872
rect 127400 59808 127408 59872
rect 127088 58784 127408 59808
rect 127088 58720 127096 58784
rect 127160 58720 127176 58784
rect 127240 58720 127256 58784
rect 127320 58720 127336 58784
rect 127400 58720 127408 58784
rect 127088 57696 127408 58720
rect 127088 57632 127096 57696
rect 127160 57632 127176 57696
rect 127240 57632 127256 57696
rect 127320 57632 127336 57696
rect 127400 57632 127408 57696
rect 127088 56608 127408 57632
rect 127088 56544 127096 56608
rect 127160 56544 127176 56608
rect 127240 56544 127256 56608
rect 127320 56544 127336 56608
rect 127400 56544 127408 56608
rect 127088 55520 127408 56544
rect 127088 55456 127096 55520
rect 127160 55456 127176 55520
rect 127240 55456 127256 55520
rect 127320 55456 127336 55520
rect 127400 55456 127408 55520
rect 127088 54432 127408 55456
rect 127088 54368 127096 54432
rect 127160 54368 127176 54432
rect 127240 54368 127256 54432
rect 127320 54368 127336 54432
rect 127400 54368 127408 54432
rect 127088 53344 127408 54368
rect 127088 53280 127096 53344
rect 127160 53280 127176 53344
rect 127240 53280 127256 53344
rect 127320 53280 127336 53344
rect 127400 53280 127408 53344
rect 127088 52256 127408 53280
rect 127088 52192 127096 52256
rect 127160 52192 127176 52256
rect 127240 52192 127256 52256
rect 127320 52192 127336 52256
rect 127400 52192 127408 52256
rect 127088 51168 127408 52192
rect 127088 51104 127096 51168
rect 127160 51104 127176 51168
rect 127240 51104 127256 51168
rect 127320 51104 127336 51168
rect 127400 51104 127408 51168
rect 127088 50080 127408 51104
rect 127088 50016 127096 50080
rect 127160 50016 127176 50080
rect 127240 50016 127256 50080
rect 127320 50016 127336 50080
rect 127400 50016 127408 50080
rect 127088 48992 127408 50016
rect 127088 48928 127096 48992
rect 127160 48928 127176 48992
rect 127240 48928 127256 48992
rect 127320 48928 127336 48992
rect 127400 48928 127408 48992
rect 127088 47904 127408 48928
rect 127088 47840 127096 47904
rect 127160 47840 127176 47904
rect 127240 47840 127256 47904
rect 127320 47840 127336 47904
rect 127400 47840 127408 47904
rect 127088 46816 127408 47840
rect 127088 46752 127096 46816
rect 127160 46752 127176 46816
rect 127240 46752 127256 46816
rect 127320 46752 127336 46816
rect 127400 46752 127408 46816
rect 127088 45728 127408 46752
rect 127088 45664 127096 45728
rect 127160 45664 127176 45728
rect 127240 45664 127256 45728
rect 127320 45664 127336 45728
rect 127400 45664 127408 45728
rect 127088 44640 127408 45664
rect 127088 44576 127096 44640
rect 127160 44576 127176 44640
rect 127240 44576 127256 44640
rect 127320 44576 127336 44640
rect 127400 44576 127408 44640
rect 127088 43552 127408 44576
rect 127088 43488 127096 43552
rect 127160 43488 127176 43552
rect 127240 43488 127256 43552
rect 127320 43488 127336 43552
rect 127400 43488 127408 43552
rect 127088 42464 127408 43488
rect 127088 42400 127096 42464
rect 127160 42400 127176 42464
rect 127240 42400 127256 42464
rect 127320 42400 127336 42464
rect 127400 42400 127408 42464
rect 127088 41376 127408 42400
rect 127088 41312 127096 41376
rect 127160 41312 127176 41376
rect 127240 41312 127256 41376
rect 127320 41312 127336 41376
rect 127400 41312 127408 41376
rect 127088 40288 127408 41312
rect 127088 40224 127096 40288
rect 127160 40224 127176 40288
rect 127240 40224 127256 40288
rect 127320 40224 127336 40288
rect 127400 40224 127408 40288
rect 127088 39200 127408 40224
rect 127088 39136 127096 39200
rect 127160 39136 127176 39200
rect 127240 39136 127256 39200
rect 127320 39136 127336 39200
rect 127400 39136 127408 39200
rect 127088 38112 127408 39136
rect 127088 38048 127096 38112
rect 127160 38048 127176 38112
rect 127240 38048 127256 38112
rect 127320 38048 127336 38112
rect 127400 38048 127408 38112
rect 127088 37024 127408 38048
rect 127088 36960 127096 37024
rect 127160 36960 127176 37024
rect 127240 36960 127256 37024
rect 127320 36960 127336 37024
rect 127400 36960 127408 37024
rect 127088 35936 127408 36960
rect 127088 35872 127096 35936
rect 127160 35872 127176 35936
rect 127240 35872 127256 35936
rect 127320 35872 127336 35936
rect 127400 35872 127408 35936
rect 127088 34848 127408 35872
rect 127088 34784 127096 34848
rect 127160 34784 127176 34848
rect 127240 34784 127256 34848
rect 127320 34784 127336 34848
rect 127400 34784 127408 34848
rect 127088 33760 127408 34784
rect 127088 33696 127096 33760
rect 127160 33696 127176 33760
rect 127240 33696 127256 33760
rect 127320 33696 127336 33760
rect 127400 33696 127408 33760
rect 127088 32672 127408 33696
rect 127088 32608 127096 32672
rect 127160 32608 127176 32672
rect 127240 32608 127256 32672
rect 127320 32608 127336 32672
rect 127400 32608 127408 32672
rect 127088 31584 127408 32608
rect 127088 31520 127096 31584
rect 127160 31520 127176 31584
rect 127240 31520 127256 31584
rect 127320 31520 127336 31584
rect 127400 31520 127408 31584
rect 127088 30496 127408 31520
rect 127088 30432 127096 30496
rect 127160 30432 127176 30496
rect 127240 30432 127256 30496
rect 127320 30432 127336 30496
rect 127400 30432 127408 30496
rect 127088 29408 127408 30432
rect 127088 29344 127096 29408
rect 127160 29344 127176 29408
rect 127240 29344 127256 29408
rect 127320 29344 127336 29408
rect 127400 29344 127408 29408
rect 127088 28320 127408 29344
rect 127088 28256 127096 28320
rect 127160 28256 127176 28320
rect 127240 28256 127256 28320
rect 127320 28256 127336 28320
rect 127400 28256 127408 28320
rect 127088 27232 127408 28256
rect 127088 27168 127096 27232
rect 127160 27168 127176 27232
rect 127240 27168 127256 27232
rect 127320 27168 127336 27232
rect 127400 27168 127408 27232
rect 127088 26144 127408 27168
rect 127088 26080 127096 26144
rect 127160 26080 127176 26144
rect 127240 26080 127256 26144
rect 127320 26080 127336 26144
rect 127400 26080 127408 26144
rect 127088 25056 127408 26080
rect 127088 24992 127096 25056
rect 127160 24992 127176 25056
rect 127240 24992 127256 25056
rect 127320 24992 127336 25056
rect 127400 24992 127408 25056
rect 127088 23968 127408 24992
rect 127088 23904 127096 23968
rect 127160 23904 127176 23968
rect 127240 23904 127256 23968
rect 127320 23904 127336 23968
rect 127400 23904 127408 23968
rect 127088 22880 127408 23904
rect 127088 22816 127096 22880
rect 127160 22816 127176 22880
rect 127240 22816 127256 22880
rect 127320 22816 127336 22880
rect 127400 22816 127408 22880
rect 127088 21792 127408 22816
rect 127088 21728 127096 21792
rect 127160 21728 127176 21792
rect 127240 21728 127256 21792
rect 127320 21728 127336 21792
rect 127400 21728 127408 21792
rect 127088 20704 127408 21728
rect 127088 20640 127096 20704
rect 127160 20640 127176 20704
rect 127240 20640 127256 20704
rect 127320 20640 127336 20704
rect 127400 20640 127408 20704
rect 127088 19616 127408 20640
rect 127088 19552 127096 19616
rect 127160 19552 127176 19616
rect 127240 19552 127256 19616
rect 127320 19552 127336 19616
rect 127400 19552 127408 19616
rect 127088 18528 127408 19552
rect 127088 18464 127096 18528
rect 127160 18464 127176 18528
rect 127240 18464 127256 18528
rect 127320 18464 127336 18528
rect 127400 18464 127408 18528
rect 127088 17440 127408 18464
rect 127088 17376 127096 17440
rect 127160 17376 127176 17440
rect 127240 17376 127256 17440
rect 127320 17376 127336 17440
rect 127400 17376 127408 17440
rect 127088 16352 127408 17376
rect 127088 16288 127096 16352
rect 127160 16288 127176 16352
rect 127240 16288 127256 16352
rect 127320 16288 127336 16352
rect 127400 16288 127408 16352
rect 127088 15264 127408 16288
rect 127088 15200 127096 15264
rect 127160 15200 127176 15264
rect 127240 15200 127256 15264
rect 127320 15200 127336 15264
rect 127400 15200 127408 15264
rect 127088 14176 127408 15200
rect 127088 14112 127096 14176
rect 127160 14112 127176 14176
rect 127240 14112 127256 14176
rect 127320 14112 127336 14176
rect 127400 14112 127408 14176
rect 127088 13088 127408 14112
rect 127088 13024 127096 13088
rect 127160 13024 127176 13088
rect 127240 13024 127256 13088
rect 127320 13024 127336 13088
rect 127400 13024 127408 13088
rect 127088 12000 127408 13024
rect 127088 11936 127096 12000
rect 127160 11936 127176 12000
rect 127240 11936 127256 12000
rect 127320 11936 127336 12000
rect 127400 11936 127408 12000
rect 127088 10912 127408 11936
rect 127088 10848 127096 10912
rect 127160 10848 127176 10912
rect 127240 10848 127256 10912
rect 127320 10848 127336 10912
rect 127400 10848 127408 10912
rect 127088 9824 127408 10848
rect 127088 9760 127096 9824
rect 127160 9760 127176 9824
rect 127240 9760 127256 9824
rect 127320 9760 127336 9824
rect 127400 9760 127408 9824
rect 127088 8736 127408 9760
rect 127088 8672 127096 8736
rect 127160 8672 127176 8736
rect 127240 8672 127256 8736
rect 127320 8672 127336 8736
rect 127400 8672 127408 8736
rect 127088 7648 127408 8672
rect 127088 7584 127096 7648
rect 127160 7584 127176 7648
rect 127240 7584 127256 7648
rect 127320 7584 127336 7648
rect 127400 7584 127408 7648
rect 127088 6560 127408 7584
rect 127088 6496 127096 6560
rect 127160 6496 127176 6560
rect 127240 6496 127256 6560
rect 127320 6496 127336 6560
rect 127400 6496 127408 6560
rect 127088 5472 127408 6496
rect 127088 5408 127096 5472
rect 127160 5408 127176 5472
rect 127240 5408 127256 5472
rect 127320 5408 127336 5472
rect 127400 5408 127408 5472
rect 127088 4384 127408 5408
rect 127088 4320 127096 4384
rect 127160 4320 127176 4384
rect 127240 4320 127256 4384
rect 127320 4320 127336 4384
rect 127400 4320 127408 4384
rect 127088 3296 127408 4320
rect 127088 3232 127096 3296
rect 127160 3232 127176 3296
rect 127240 3232 127256 3296
rect 127320 3232 127336 3296
rect 127400 3232 127408 3296
rect 127088 2208 127408 3232
rect 127088 2144 127096 2208
rect 127160 2144 127176 2208
rect 127240 2144 127256 2208
rect 127320 2144 127336 2208
rect 127400 2144 127408 2208
rect 127748 2176 128068 117504
rect 128408 2176 128728 117504
rect 129068 2176 129388 117504
rect 142448 116992 142768 117552
rect 157808 117536 158128 117552
rect 142448 116928 142456 116992
rect 142520 116928 142536 116992
rect 142600 116928 142616 116992
rect 142680 116928 142696 116992
rect 142760 116928 142768 116992
rect 142448 115904 142768 116928
rect 142448 115840 142456 115904
rect 142520 115840 142536 115904
rect 142600 115840 142616 115904
rect 142680 115840 142696 115904
rect 142760 115840 142768 115904
rect 142448 114816 142768 115840
rect 142448 114752 142456 114816
rect 142520 114752 142536 114816
rect 142600 114752 142616 114816
rect 142680 114752 142696 114816
rect 142760 114752 142768 114816
rect 142448 113728 142768 114752
rect 142448 113664 142456 113728
rect 142520 113664 142536 113728
rect 142600 113664 142616 113728
rect 142680 113664 142696 113728
rect 142760 113664 142768 113728
rect 142448 112640 142768 113664
rect 142448 112576 142456 112640
rect 142520 112576 142536 112640
rect 142600 112576 142616 112640
rect 142680 112576 142696 112640
rect 142760 112576 142768 112640
rect 142448 111552 142768 112576
rect 142448 111488 142456 111552
rect 142520 111488 142536 111552
rect 142600 111488 142616 111552
rect 142680 111488 142696 111552
rect 142760 111488 142768 111552
rect 142448 110464 142768 111488
rect 142448 110400 142456 110464
rect 142520 110400 142536 110464
rect 142600 110400 142616 110464
rect 142680 110400 142696 110464
rect 142760 110400 142768 110464
rect 142448 109376 142768 110400
rect 142448 109312 142456 109376
rect 142520 109312 142536 109376
rect 142600 109312 142616 109376
rect 142680 109312 142696 109376
rect 142760 109312 142768 109376
rect 142448 108288 142768 109312
rect 142448 108224 142456 108288
rect 142520 108224 142536 108288
rect 142600 108224 142616 108288
rect 142680 108224 142696 108288
rect 142760 108224 142768 108288
rect 142448 107200 142768 108224
rect 142448 107136 142456 107200
rect 142520 107136 142536 107200
rect 142600 107136 142616 107200
rect 142680 107136 142696 107200
rect 142760 107136 142768 107200
rect 142448 106112 142768 107136
rect 142448 106048 142456 106112
rect 142520 106048 142536 106112
rect 142600 106048 142616 106112
rect 142680 106048 142696 106112
rect 142760 106048 142768 106112
rect 142448 105024 142768 106048
rect 142448 104960 142456 105024
rect 142520 104960 142536 105024
rect 142600 104960 142616 105024
rect 142680 104960 142696 105024
rect 142760 104960 142768 105024
rect 142448 103936 142768 104960
rect 142448 103872 142456 103936
rect 142520 103872 142536 103936
rect 142600 103872 142616 103936
rect 142680 103872 142696 103936
rect 142760 103872 142768 103936
rect 142448 102848 142768 103872
rect 142448 102784 142456 102848
rect 142520 102784 142536 102848
rect 142600 102784 142616 102848
rect 142680 102784 142696 102848
rect 142760 102784 142768 102848
rect 142448 101760 142768 102784
rect 142448 101696 142456 101760
rect 142520 101696 142536 101760
rect 142600 101696 142616 101760
rect 142680 101696 142696 101760
rect 142760 101696 142768 101760
rect 142448 100672 142768 101696
rect 142448 100608 142456 100672
rect 142520 100608 142536 100672
rect 142600 100608 142616 100672
rect 142680 100608 142696 100672
rect 142760 100608 142768 100672
rect 142448 99584 142768 100608
rect 142448 99520 142456 99584
rect 142520 99520 142536 99584
rect 142600 99520 142616 99584
rect 142680 99520 142696 99584
rect 142760 99520 142768 99584
rect 142448 98496 142768 99520
rect 142448 98432 142456 98496
rect 142520 98432 142536 98496
rect 142600 98432 142616 98496
rect 142680 98432 142696 98496
rect 142760 98432 142768 98496
rect 142448 97408 142768 98432
rect 142448 97344 142456 97408
rect 142520 97344 142536 97408
rect 142600 97344 142616 97408
rect 142680 97344 142696 97408
rect 142760 97344 142768 97408
rect 142448 96320 142768 97344
rect 142448 96256 142456 96320
rect 142520 96256 142536 96320
rect 142600 96256 142616 96320
rect 142680 96256 142696 96320
rect 142760 96256 142768 96320
rect 142448 95232 142768 96256
rect 142448 95168 142456 95232
rect 142520 95168 142536 95232
rect 142600 95168 142616 95232
rect 142680 95168 142696 95232
rect 142760 95168 142768 95232
rect 142448 94144 142768 95168
rect 142448 94080 142456 94144
rect 142520 94080 142536 94144
rect 142600 94080 142616 94144
rect 142680 94080 142696 94144
rect 142760 94080 142768 94144
rect 142448 93056 142768 94080
rect 142448 92992 142456 93056
rect 142520 92992 142536 93056
rect 142600 92992 142616 93056
rect 142680 92992 142696 93056
rect 142760 92992 142768 93056
rect 142448 91968 142768 92992
rect 142448 91904 142456 91968
rect 142520 91904 142536 91968
rect 142600 91904 142616 91968
rect 142680 91904 142696 91968
rect 142760 91904 142768 91968
rect 142448 90880 142768 91904
rect 142448 90816 142456 90880
rect 142520 90816 142536 90880
rect 142600 90816 142616 90880
rect 142680 90816 142696 90880
rect 142760 90816 142768 90880
rect 142448 89792 142768 90816
rect 142448 89728 142456 89792
rect 142520 89728 142536 89792
rect 142600 89728 142616 89792
rect 142680 89728 142696 89792
rect 142760 89728 142768 89792
rect 142448 88704 142768 89728
rect 142448 88640 142456 88704
rect 142520 88640 142536 88704
rect 142600 88640 142616 88704
rect 142680 88640 142696 88704
rect 142760 88640 142768 88704
rect 142448 87616 142768 88640
rect 142448 87552 142456 87616
rect 142520 87552 142536 87616
rect 142600 87552 142616 87616
rect 142680 87552 142696 87616
rect 142760 87552 142768 87616
rect 142448 86528 142768 87552
rect 142448 86464 142456 86528
rect 142520 86464 142536 86528
rect 142600 86464 142616 86528
rect 142680 86464 142696 86528
rect 142760 86464 142768 86528
rect 142448 85440 142768 86464
rect 142448 85376 142456 85440
rect 142520 85376 142536 85440
rect 142600 85376 142616 85440
rect 142680 85376 142696 85440
rect 142760 85376 142768 85440
rect 142448 84352 142768 85376
rect 142448 84288 142456 84352
rect 142520 84288 142536 84352
rect 142600 84288 142616 84352
rect 142680 84288 142696 84352
rect 142760 84288 142768 84352
rect 142448 83264 142768 84288
rect 142448 83200 142456 83264
rect 142520 83200 142536 83264
rect 142600 83200 142616 83264
rect 142680 83200 142696 83264
rect 142760 83200 142768 83264
rect 142448 82176 142768 83200
rect 142448 82112 142456 82176
rect 142520 82112 142536 82176
rect 142600 82112 142616 82176
rect 142680 82112 142696 82176
rect 142760 82112 142768 82176
rect 142448 81088 142768 82112
rect 142448 81024 142456 81088
rect 142520 81024 142536 81088
rect 142600 81024 142616 81088
rect 142680 81024 142696 81088
rect 142760 81024 142768 81088
rect 142448 80000 142768 81024
rect 142448 79936 142456 80000
rect 142520 79936 142536 80000
rect 142600 79936 142616 80000
rect 142680 79936 142696 80000
rect 142760 79936 142768 80000
rect 142448 78912 142768 79936
rect 142448 78848 142456 78912
rect 142520 78848 142536 78912
rect 142600 78848 142616 78912
rect 142680 78848 142696 78912
rect 142760 78848 142768 78912
rect 142448 77824 142768 78848
rect 142448 77760 142456 77824
rect 142520 77760 142536 77824
rect 142600 77760 142616 77824
rect 142680 77760 142696 77824
rect 142760 77760 142768 77824
rect 142448 76736 142768 77760
rect 142448 76672 142456 76736
rect 142520 76672 142536 76736
rect 142600 76672 142616 76736
rect 142680 76672 142696 76736
rect 142760 76672 142768 76736
rect 142448 75648 142768 76672
rect 142448 75584 142456 75648
rect 142520 75584 142536 75648
rect 142600 75584 142616 75648
rect 142680 75584 142696 75648
rect 142760 75584 142768 75648
rect 142448 74560 142768 75584
rect 142448 74496 142456 74560
rect 142520 74496 142536 74560
rect 142600 74496 142616 74560
rect 142680 74496 142696 74560
rect 142760 74496 142768 74560
rect 142448 73472 142768 74496
rect 142448 73408 142456 73472
rect 142520 73408 142536 73472
rect 142600 73408 142616 73472
rect 142680 73408 142696 73472
rect 142760 73408 142768 73472
rect 142448 72384 142768 73408
rect 142448 72320 142456 72384
rect 142520 72320 142536 72384
rect 142600 72320 142616 72384
rect 142680 72320 142696 72384
rect 142760 72320 142768 72384
rect 142448 71296 142768 72320
rect 142448 71232 142456 71296
rect 142520 71232 142536 71296
rect 142600 71232 142616 71296
rect 142680 71232 142696 71296
rect 142760 71232 142768 71296
rect 142448 70208 142768 71232
rect 142448 70144 142456 70208
rect 142520 70144 142536 70208
rect 142600 70144 142616 70208
rect 142680 70144 142696 70208
rect 142760 70144 142768 70208
rect 142448 69120 142768 70144
rect 142448 69056 142456 69120
rect 142520 69056 142536 69120
rect 142600 69056 142616 69120
rect 142680 69056 142696 69120
rect 142760 69056 142768 69120
rect 142448 68032 142768 69056
rect 142448 67968 142456 68032
rect 142520 67968 142536 68032
rect 142600 67968 142616 68032
rect 142680 67968 142696 68032
rect 142760 67968 142768 68032
rect 142448 66944 142768 67968
rect 142448 66880 142456 66944
rect 142520 66880 142536 66944
rect 142600 66880 142616 66944
rect 142680 66880 142696 66944
rect 142760 66880 142768 66944
rect 142448 65856 142768 66880
rect 142448 65792 142456 65856
rect 142520 65792 142536 65856
rect 142600 65792 142616 65856
rect 142680 65792 142696 65856
rect 142760 65792 142768 65856
rect 142448 64768 142768 65792
rect 142448 64704 142456 64768
rect 142520 64704 142536 64768
rect 142600 64704 142616 64768
rect 142680 64704 142696 64768
rect 142760 64704 142768 64768
rect 142448 63680 142768 64704
rect 142448 63616 142456 63680
rect 142520 63616 142536 63680
rect 142600 63616 142616 63680
rect 142680 63616 142696 63680
rect 142760 63616 142768 63680
rect 142448 62592 142768 63616
rect 142448 62528 142456 62592
rect 142520 62528 142536 62592
rect 142600 62528 142616 62592
rect 142680 62528 142696 62592
rect 142760 62528 142768 62592
rect 142448 61504 142768 62528
rect 142448 61440 142456 61504
rect 142520 61440 142536 61504
rect 142600 61440 142616 61504
rect 142680 61440 142696 61504
rect 142760 61440 142768 61504
rect 142448 60416 142768 61440
rect 142448 60352 142456 60416
rect 142520 60352 142536 60416
rect 142600 60352 142616 60416
rect 142680 60352 142696 60416
rect 142760 60352 142768 60416
rect 142448 59328 142768 60352
rect 142448 59264 142456 59328
rect 142520 59264 142536 59328
rect 142600 59264 142616 59328
rect 142680 59264 142696 59328
rect 142760 59264 142768 59328
rect 142448 58240 142768 59264
rect 142448 58176 142456 58240
rect 142520 58176 142536 58240
rect 142600 58176 142616 58240
rect 142680 58176 142696 58240
rect 142760 58176 142768 58240
rect 142448 57152 142768 58176
rect 142448 57088 142456 57152
rect 142520 57088 142536 57152
rect 142600 57088 142616 57152
rect 142680 57088 142696 57152
rect 142760 57088 142768 57152
rect 142448 56064 142768 57088
rect 142448 56000 142456 56064
rect 142520 56000 142536 56064
rect 142600 56000 142616 56064
rect 142680 56000 142696 56064
rect 142760 56000 142768 56064
rect 142448 54976 142768 56000
rect 142448 54912 142456 54976
rect 142520 54912 142536 54976
rect 142600 54912 142616 54976
rect 142680 54912 142696 54976
rect 142760 54912 142768 54976
rect 142448 53888 142768 54912
rect 142448 53824 142456 53888
rect 142520 53824 142536 53888
rect 142600 53824 142616 53888
rect 142680 53824 142696 53888
rect 142760 53824 142768 53888
rect 142448 52800 142768 53824
rect 142448 52736 142456 52800
rect 142520 52736 142536 52800
rect 142600 52736 142616 52800
rect 142680 52736 142696 52800
rect 142760 52736 142768 52800
rect 142448 51712 142768 52736
rect 142448 51648 142456 51712
rect 142520 51648 142536 51712
rect 142600 51648 142616 51712
rect 142680 51648 142696 51712
rect 142760 51648 142768 51712
rect 142448 50624 142768 51648
rect 142448 50560 142456 50624
rect 142520 50560 142536 50624
rect 142600 50560 142616 50624
rect 142680 50560 142696 50624
rect 142760 50560 142768 50624
rect 142448 49536 142768 50560
rect 142448 49472 142456 49536
rect 142520 49472 142536 49536
rect 142600 49472 142616 49536
rect 142680 49472 142696 49536
rect 142760 49472 142768 49536
rect 142448 48448 142768 49472
rect 142448 48384 142456 48448
rect 142520 48384 142536 48448
rect 142600 48384 142616 48448
rect 142680 48384 142696 48448
rect 142760 48384 142768 48448
rect 142448 47360 142768 48384
rect 142448 47296 142456 47360
rect 142520 47296 142536 47360
rect 142600 47296 142616 47360
rect 142680 47296 142696 47360
rect 142760 47296 142768 47360
rect 142448 46272 142768 47296
rect 142448 46208 142456 46272
rect 142520 46208 142536 46272
rect 142600 46208 142616 46272
rect 142680 46208 142696 46272
rect 142760 46208 142768 46272
rect 142448 45184 142768 46208
rect 142448 45120 142456 45184
rect 142520 45120 142536 45184
rect 142600 45120 142616 45184
rect 142680 45120 142696 45184
rect 142760 45120 142768 45184
rect 142448 44096 142768 45120
rect 142448 44032 142456 44096
rect 142520 44032 142536 44096
rect 142600 44032 142616 44096
rect 142680 44032 142696 44096
rect 142760 44032 142768 44096
rect 142448 43008 142768 44032
rect 142448 42944 142456 43008
rect 142520 42944 142536 43008
rect 142600 42944 142616 43008
rect 142680 42944 142696 43008
rect 142760 42944 142768 43008
rect 142448 41920 142768 42944
rect 142448 41856 142456 41920
rect 142520 41856 142536 41920
rect 142600 41856 142616 41920
rect 142680 41856 142696 41920
rect 142760 41856 142768 41920
rect 142448 40832 142768 41856
rect 142448 40768 142456 40832
rect 142520 40768 142536 40832
rect 142600 40768 142616 40832
rect 142680 40768 142696 40832
rect 142760 40768 142768 40832
rect 142448 39744 142768 40768
rect 142448 39680 142456 39744
rect 142520 39680 142536 39744
rect 142600 39680 142616 39744
rect 142680 39680 142696 39744
rect 142760 39680 142768 39744
rect 142448 38656 142768 39680
rect 142448 38592 142456 38656
rect 142520 38592 142536 38656
rect 142600 38592 142616 38656
rect 142680 38592 142696 38656
rect 142760 38592 142768 38656
rect 142448 37568 142768 38592
rect 142448 37504 142456 37568
rect 142520 37504 142536 37568
rect 142600 37504 142616 37568
rect 142680 37504 142696 37568
rect 142760 37504 142768 37568
rect 142448 36480 142768 37504
rect 142448 36416 142456 36480
rect 142520 36416 142536 36480
rect 142600 36416 142616 36480
rect 142680 36416 142696 36480
rect 142760 36416 142768 36480
rect 142448 35392 142768 36416
rect 142448 35328 142456 35392
rect 142520 35328 142536 35392
rect 142600 35328 142616 35392
rect 142680 35328 142696 35392
rect 142760 35328 142768 35392
rect 142448 34304 142768 35328
rect 142448 34240 142456 34304
rect 142520 34240 142536 34304
rect 142600 34240 142616 34304
rect 142680 34240 142696 34304
rect 142760 34240 142768 34304
rect 142448 33216 142768 34240
rect 142448 33152 142456 33216
rect 142520 33152 142536 33216
rect 142600 33152 142616 33216
rect 142680 33152 142696 33216
rect 142760 33152 142768 33216
rect 142448 32128 142768 33152
rect 142448 32064 142456 32128
rect 142520 32064 142536 32128
rect 142600 32064 142616 32128
rect 142680 32064 142696 32128
rect 142760 32064 142768 32128
rect 142448 31040 142768 32064
rect 142448 30976 142456 31040
rect 142520 30976 142536 31040
rect 142600 30976 142616 31040
rect 142680 30976 142696 31040
rect 142760 30976 142768 31040
rect 142448 29952 142768 30976
rect 142448 29888 142456 29952
rect 142520 29888 142536 29952
rect 142600 29888 142616 29952
rect 142680 29888 142696 29952
rect 142760 29888 142768 29952
rect 142448 28864 142768 29888
rect 142448 28800 142456 28864
rect 142520 28800 142536 28864
rect 142600 28800 142616 28864
rect 142680 28800 142696 28864
rect 142760 28800 142768 28864
rect 142448 27776 142768 28800
rect 142448 27712 142456 27776
rect 142520 27712 142536 27776
rect 142600 27712 142616 27776
rect 142680 27712 142696 27776
rect 142760 27712 142768 27776
rect 142448 26688 142768 27712
rect 142448 26624 142456 26688
rect 142520 26624 142536 26688
rect 142600 26624 142616 26688
rect 142680 26624 142696 26688
rect 142760 26624 142768 26688
rect 142448 25600 142768 26624
rect 142448 25536 142456 25600
rect 142520 25536 142536 25600
rect 142600 25536 142616 25600
rect 142680 25536 142696 25600
rect 142760 25536 142768 25600
rect 142448 24512 142768 25536
rect 142448 24448 142456 24512
rect 142520 24448 142536 24512
rect 142600 24448 142616 24512
rect 142680 24448 142696 24512
rect 142760 24448 142768 24512
rect 142448 23424 142768 24448
rect 142448 23360 142456 23424
rect 142520 23360 142536 23424
rect 142600 23360 142616 23424
rect 142680 23360 142696 23424
rect 142760 23360 142768 23424
rect 142448 22336 142768 23360
rect 142448 22272 142456 22336
rect 142520 22272 142536 22336
rect 142600 22272 142616 22336
rect 142680 22272 142696 22336
rect 142760 22272 142768 22336
rect 142448 21248 142768 22272
rect 142448 21184 142456 21248
rect 142520 21184 142536 21248
rect 142600 21184 142616 21248
rect 142680 21184 142696 21248
rect 142760 21184 142768 21248
rect 142448 20160 142768 21184
rect 142448 20096 142456 20160
rect 142520 20096 142536 20160
rect 142600 20096 142616 20160
rect 142680 20096 142696 20160
rect 142760 20096 142768 20160
rect 142448 19072 142768 20096
rect 142448 19008 142456 19072
rect 142520 19008 142536 19072
rect 142600 19008 142616 19072
rect 142680 19008 142696 19072
rect 142760 19008 142768 19072
rect 142448 17984 142768 19008
rect 142448 17920 142456 17984
rect 142520 17920 142536 17984
rect 142600 17920 142616 17984
rect 142680 17920 142696 17984
rect 142760 17920 142768 17984
rect 142448 16896 142768 17920
rect 142448 16832 142456 16896
rect 142520 16832 142536 16896
rect 142600 16832 142616 16896
rect 142680 16832 142696 16896
rect 142760 16832 142768 16896
rect 142448 15808 142768 16832
rect 142448 15744 142456 15808
rect 142520 15744 142536 15808
rect 142600 15744 142616 15808
rect 142680 15744 142696 15808
rect 142760 15744 142768 15808
rect 142448 14720 142768 15744
rect 142448 14656 142456 14720
rect 142520 14656 142536 14720
rect 142600 14656 142616 14720
rect 142680 14656 142696 14720
rect 142760 14656 142768 14720
rect 142448 13632 142768 14656
rect 142448 13568 142456 13632
rect 142520 13568 142536 13632
rect 142600 13568 142616 13632
rect 142680 13568 142696 13632
rect 142760 13568 142768 13632
rect 142448 12544 142768 13568
rect 142448 12480 142456 12544
rect 142520 12480 142536 12544
rect 142600 12480 142616 12544
rect 142680 12480 142696 12544
rect 142760 12480 142768 12544
rect 142448 11456 142768 12480
rect 142448 11392 142456 11456
rect 142520 11392 142536 11456
rect 142600 11392 142616 11456
rect 142680 11392 142696 11456
rect 142760 11392 142768 11456
rect 142448 10368 142768 11392
rect 142448 10304 142456 10368
rect 142520 10304 142536 10368
rect 142600 10304 142616 10368
rect 142680 10304 142696 10368
rect 142760 10304 142768 10368
rect 142448 9280 142768 10304
rect 142448 9216 142456 9280
rect 142520 9216 142536 9280
rect 142600 9216 142616 9280
rect 142680 9216 142696 9280
rect 142760 9216 142768 9280
rect 142448 8192 142768 9216
rect 142448 8128 142456 8192
rect 142520 8128 142536 8192
rect 142600 8128 142616 8192
rect 142680 8128 142696 8192
rect 142760 8128 142768 8192
rect 142448 7104 142768 8128
rect 142448 7040 142456 7104
rect 142520 7040 142536 7104
rect 142600 7040 142616 7104
rect 142680 7040 142696 7104
rect 142760 7040 142768 7104
rect 142448 6016 142768 7040
rect 142448 5952 142456 6016
rect 142520 5952 142536 6016
rect 142600 5952 142616 6016
rect 142680 5952 142696 6016
rect 142760 5952 142768 6016
rect 142448 4928 142768 5952
rect 142448 4864 142456 4928
rect 142520 4864 142536 4928
rect 142600 4864 142616 4928
rect 142680 4864 142696 4928
rect 142760 4864 142768 4928
rect 142448 3840 142768 4864
rect 142448 3776 142456 3840
rect 142520 3776 142536 3840
rect 142600 3776 142616 3840
rect 142680 3776 142696 3840
rect 142760 3776 142768 3840
rect 142448 2752 142768 3776
rect 142448 2688 142456 2752
rect 142520 2688 142536 2752
rect 142600 2688 142616 2752
rect 142680 2688 142696 2752
rect 142760 2688 142768 2752
rect 127088 2128 127408 2144
rect 142448 2128 142768 2688
rect 143108 2176 143428 117504
rect 143768 2176 144088 117504
rect 144428 2176 144748 117504
rect 157808 117472 157816 117536
rect 157880 117472 157896 117536
rect 157960 117472 157976 117536
rect 158040 117472 158056 117536
rect 158120 117472 158128 117536
rect 157808 116448 158128 117472
rect 157808 116384 157816 116448
rect 157880 116384 157896 116448
rect 157960 116384 157976 116448
rect 158040 116384 158056 116448
rect 158120 116384 158128 116448
rect 157808 115360 158128 116384
rect 157808 115296 157816 115360
rect 157880 115296 157896 115360
rect 157960 115296 157976 115360
rect 158040 115296 158056 115360
rect 158120 115296 158128 115360
rect 157808 114272 158128 115296
rect 157808 114208 157816 114272
rect 157880 114208 157896 114272
rect 157960 114208 157976 114272
rect 158040 114208 158056 114272
rect 158120 114208 158128 114272
rect 157808 113184 158128 114208
rect 157808 113120 157816 113184
rect 157880 113120 157896 113184
rect 157960 113120 157976 113184
rect 158040 113120 158056 113184
rect 158120 113120 158128 113184
rect 157808 112096 158128 113120
rect 157808 112032 157816 112096
rect 157880 112032 157896 112096
rect 157960 112032 157976 112096
rect 158040 112032 158056 112096
rect 158120 112032 158128 112096
rect 157808 111008 158128 112032
rect 157808 110944 157816 111008
rect 157880 110944 157896 111008
rect 157960 110944 157976 111008
rect 158040 110944 158056 111008
rect 158120 110944 158128 111008
rect 157808 109920 158128 110944
rect 157808 109856 157816 109920
rect 157880 109856 157896 109920
rect 157960 109856 157976 109920
rect 158040 109856 158056 109920
rect 158120 109856 158128 109920
rect 157808 108832 158128 109856
rect 157808 108768 157816 108832
rect 157880 108768 157896 108832
rect 157960 108768 157976 108832
rect 158040 108768 158056 108832
rect 158120 108768 158128 108832
rect 157808 107744 158128 108768
rect 157808 107680 157816 107744
rect 157880 107680 157896 107744
rect 157960 107680 157976 107744
rect 158040 107680 158056 107744
rect 158120 107680 158128 107744
rect 157808 106656 158128 107680
rect 157808 106592 157816 106656
rect 157880 106592 157896 106656
rect 157960 106592 157976 106656
rect 158040 106592 158056 106656
rect 158120 106592 158128 106656
rect 157808 105568 158128 106592
rect 157808 105504 157816 105568
rect 157880 105504 157896 105568
rect 157960 105504 157976 105568
rect 158040 105504 158056 105568
rect 158120 105504 158128 105568
rect 157808 104480 158128 105504
rect 157808 104416 157816 104480
rect 157880 104416 157896 104480
rect 157960 104416 157976 104480
rect 158040 104416 158056 104480
rect 158120 104416 158128 104480
rect 157808 103392 158128 104416
rect 157808 103328 157816 103392
rect 157880 103328 157896 103392
rect 157960 103328 157976 103392
rect 158040 103328 158056 103392
rect 158120 103328 158128 103392
rect 157808 102304 158128 103328
rect 157808 102240 157816 102304
rect 157880 102240 157896 102304
rect 157960 102240 157976 102304
rect 158040 102240 158056 102304
rect 158120 102240 158128 102304
rect 157808 101216 158128 102240
rect 157808 101152 157816 101216
rect 157880 101152 157896 101216
rect 157960 101152 157976 101216
rect 158040 101152 158056 101216
rect 158120 101152 158128 101216
rect 157808 100128 158128 101152
rect 157808 100064 157816 100128
rect 157880 100064 157896 100128
rect 157960 100064 157976 100128
rect 158040 100064 158056 100128
rect 158120 100064 158128 100128
rect 157808 99040 158128 100064
rect 157808 98976 157816 99040
rect 157880 98976 157896 99040
rect 157960 98976 157976 99040
rect 158040 98976 158056 99040
rect 158120 98976 158128 99040
rect 157808 97952 158128 98976
rect 157808 97888 157816 97952
rect 157880 97888 157896 97952
rect 157960 97888 157976 97952
rect 158040 97888 158056 97952
rect 158120 97888 158128 97952
rect 157808 96864 158128 97888
rect 157808 96800 157816 96864
rect 157880 96800 157896 96864
rect 157960 96800 157976 96864
rect 158040 96800 158056 96864
rect 158120 96800 158128 96864
rect 157808 95776 158128 96800
rect 157808 95712 157816 95776
rect 157880 95712 157896 95776
rect 157960 95712 157976 95776
rect 158040 95712 158056 95776
rect 158120 95712 158128 95776
rect 157808 94688 158128 95712
rect 157808 94624 157816 94688
rect 157880 94624 157896 94688
rect 157960 94624 157976 94688
rect 158040 94624 158056 94688
rect 158120 94624 158128 94688
rect 157808 93600 158128 94624
rect 157808 93536 157816 93600
rect 157880 93536 157896 93600
rect 157960 93536 157976 93600
rect 158040 93536 158056 93600
rect 158120 93536 158128 93600
rect 157808 92512 158128 93536
rect 157808 92448 157816 92512
rect 157880 92448 157896 92512
rect 157960 92448 157976 92512
rect 158040 92448 158056 92512
rect 158120 92448 158128 92512
rect 157808 91424 158128 92448
rect 157808 91360 157816 91424
rect 157880 91360 157896 91424
rect 157960 91360 157976 91424
rect 158040 91360 158056 91424
rect 158120 91360 158128 91424
rect 157808 90336 158128 91360
rect 157808 90272 157816 90336
rect 157880 90272 157896 90336
rect 157960 90272 157976 90336
rect 158040 90272 158056 90336
rect 158120 90272 158128 90336
rect 157808 89248 158128 90272
rect 157808 89184 157816 89248
rect 157880 89184 157896 89248
rect 157960 89184 157976 89248
rect 158040 89184 158056 89248
rect 158120 89184 158128 89248
rect 157808 88160 158128 89184
rect 157808 88096 157816 88160
rect 157880 88096 157896 88160
rect 157960 88096 157976 88160
rect 158040 88096 158056 88160
rect 158120 88096 158128 88160
rect 157808 87072 158128 88096
rect 157808 87008 157816 87072
rect 157880 87008 157896 87072
rect 157960 87008 157976 87072
rect 158040 87008 158056 87072
rect 158120 87008 158128 87072
rect 157808 85984 158128 87008
rect 157808 85920 157816 85984
rect 157880 85920 157896 85984
rect 157960 85920 157976 85984
rect 158040 85920 158056 85984
rect 158120 85920 158128 85984
rect 157808 84896 158128 85920
rect 157808 84832 157816 84896
rect 157880 84832 157896 84896
rect 157960 84832 157976 84896
rect 158040 84832 158056 84896
rect 158120 84832 158128 84896
rect 157808 83808 158128 84832
rect 157808 83744 157816 83808
rect 157880 83744 157896 83808
rect 157960 83744 157976 83808
rect 158040 83744 158056 83808
rect 158120 83744 158128 83808
rect 157808 82720 158128 83744
rect 157808 82656 157816 82720
rect 157880 82656 157896 82720
rect 157960 82656 157976 82720
rect 158040 82656 158056 82720
rect 158120 82656 158128 82720
rect 157808 81632 158128 82656
rect 157808 81568 157816 81632
rect 157880 81568 157896 81632
rect 157960 81568 157976 81632
rect 158040 81568 158056 81632
rect 158120 81568 158128 81632
rect 157808 80544 158128 81568
rect 157808 80480 157816 80544
rect 157880 80480 157896 80544
rect 157960 80480 157976 80544
rect 158040 80480 158056 80544
rect 158120 80480 158128 80544
rect 157808 79456 158128 80480
rect 157808 79392 157816 79456
rect 157880 79392 157896 79456
rect 157960 79392 157976 79456
rect 158040 79392 158056 79456
rect 158120 79392 158128 79456
rect 157808 78368 158128 79392
rect 157808 78304 157816 78368
rect 157880 78304 157896 78368
rect 157960 78304 157976 78368
rect 158040 78304 158056 78368
rect 158120 78304 158128 78368
rect 157808 77280 158128 78304
rect 157808 77216 157816 77280
rect 157880 77216 157896 77280
rect 157960 77216 157976 77280
rect 158040 77216 158056 77280
rect 158120 77216 158128 77280
rect 157808 76192 158128 77216
rect 157808 76128 157816 76192
rect 157880 76128 157896 76192
rect 157960 76128 157976 76192
rect 158040 76128 158056 76192
rect 158120 76128 158128 76192
rect 157808 75104 158128 76128
rect 157808 75040 157816 75104
rect 157880 75040 157896 75104
rect 157960 75040 157976 75104
rect 158040 75040 158056 75104
rect 158120 75040 158128 75104
rect 157808 74016 158128 75040
rect 157808 73952 157816 74016
rect 157880 73952 157896 74016
rect 157960 73952 157976 74016
rect 158040 73952 158056 74016
rect 158120 73952 158128 74016
rect 157808 72928 158128 73952
rect 157808 72864 157816 72928
rect 157880 72864 157896 72928
rect 157960 72864 157976 72928
rect 158040 72864 158056 72928
rect 158120 72864 158128 72928
rect 157808 71840 158128 72864
rect 157808 71776 157816 71840
rect 157880 71776 157896 71840
rect 157960 71776 157976 71840
rect 158040 71776 158056 71840
rect 158120 71776 158128 71840
rect 157808 70752 158128 71776
rect 157808 70688 157816 70752
rect 157880 70688 157896 70752
rect 157960 70688 157976 70752
rect 158040 70688 158056 70752
rect 158120 70688 158128 70752
rect 157808 69664 158128 70688
rect 157808 69600 157816 69664
rect 157880 69600 157896 69664
rect 157960 69600 157976 69664
rect 158040 69600 158056 69664
rect 158120 69600 158128 69664
rect 157808 68576 158128 69600
rect 157808 68512 157816 68576
rect 157880 68512 157896 68576
rect 157960 68512 157976 68576
rect 158040 68512 158056 68576
rect 158120 68512 158128 68576
rect 157808 67488 158128 68512
rect 157808 67424 157816 67488
rect 157880 67424 157896 67488
rect 157960 67424 157976 67488
rect 158040 67424 158056 67488
rect 158120 67424 158128 67488
rect 157808 66400 158128 67424
rect 157808 66336 157816 66400
rect 157880 66336 157896 66400
rect 157960 66336 157976 66400
rect 158040 66336 158056 66400
rect 158120 66336 158128 66400
rect 157808 65312 158128 66336
rect 157808 65248 157816 65312
rect 157880 65248 157896 65312
rect 157960 65248 157976 65312
rect 158040 65248 158056 65312
rect 158120 65248 158128 65312
rect 157808 64224 158128 65248
rect 157808 64160 157816 64224
rect 157880 64160 157896 64224
rect 157960 64160 157976 64224
rect 158040 64160 158056 64224
rect 158120 64160 158128 64224
rect 157808 63136 158128 64160
rect 157808 63072 157816 63136
rect 157880 63072 157896 63136
rect 157960 63072 157976 63136
rect 158040 63072 158056 63136
rect 158120 63072 158128 63136
rect 157808 62048 158128 63072
rect 157808 61984 157816 62048
rect 157880 61984 157896 62048
rect 157960 61984 157976 62048
rect 158040 61984 158056 62048
rect 158120 61984 158128 62048
rect 157808 60960 158128 61984
rect 157808 60896 157816 60960
rect 157880 60896 157896 60960
rect 157960 60896 157976 60960
rect 158040 60896 158056 60960
rect 158120 60896 158128 60960
rect 157808 59872 158128 60896
rect 157808 59808 157816 59872
rect 157880 59808 157896 59872
rect 157960 59808 157976 59872
rect 158040 59808 158056 59872
rect 158120 59808 158128 59872
rect 157808 58784 158128 59808
rect 157808 58720 157816 58784
rect 157880 58720 157896 58784
rect 157960 58720 157976 58784
rect 158040 58720 158056 58784
rect 158120 58720 158128 58784
rect 157808 57696 158128 58720
rect 157808 57632 157816 57696
rect 157880 57632 157896 57696
rect 157960 57632 157976 57696
rect 158040 57632 158056 57696
rect 158120 57632 158128 57696
rect 157808 56608 158128 57632
rect 157808 56544 157816 56608
rect 157880 56544 157896 56608
rect 157960 56544 157976 56608
rect 158040 56544 158056 56608
rect 158120 56544 158128 56608
rect 157808 55520 158128 56544
rect 157808 55456 157816 55520
rect 157880 55456 157896 55520
rect 157960 55456 157976 55520
rect 158040 55456 158056 55520
rect 158120 55456 158128 55520
rect 157808 54432 158128 55456
rect 157808 54368 157816 54432
rect 157880 54368 157896 54432
rect 157960 54368 157976 54432
rect 158040 54368 158056 54432
rect 158120 54368 158128 54432
rect 157808 53344 158128 54368
rect 157808 53280 157816 53344
rect 157880 53280 157896 53344
rect 157960 53280 157976 53344
rect 158040 53280 158056 53344
rect 158120 53280 158128 53344
rect 157808 52256 158128 53280
rect 157808 52192 157816 52256
rect 157880 52192 157896 52256
rect 157960 52192 157976 52256
rect 158040 52192 158056 52256
rect 158120 52192 158128 52256
rect 157808 51168 158128 52192
rect 157808 51104 157816 51168
rect 157880 51104 157896 51168
rect 157960 51104 157976 51168
rect 158040 51104 158056 51168
rect 158120 51104 158128 51168
rect 157808 50080 158128 51104
rect 157808 50016 157816 50080
rect 157880 50016 157896 50080
rect 157960 50016 157976 50080
rect 158040 50016 158056 50080
rect 158120 50016 158128 50080
rect 157808 48992 158128 50016
rect 157808 48928 157816 48992
rect 157880 48928 157896 48992
rect 157960 48928 157976 48992
rect 158040 48928 158056 48992
rect 158120 48928 158128 48992
rect 157808 47904 158128 48928
rect 157808 47840 157816 47904
rect 157880 47840 157896 47904
rect 157960 47840 157976 47904
rect 158040 47840 158056 47904
rect 158120 47840 158128 47904
rect 157808 46816 158128 47840
rect 157808 46752 157816 46816
rect 157880 46752 157896 46816
rect 157960 46752 157976 46816
rect 158040 46752 158056 46816
rect 158120 46752 158128 46816
rect 157808 45728 158128 46752
rect 157808 45664 157816 45728
rect 157880 45664 157896 45728
rect 157960 45664 157976 45728
rect 158040 45664 158056 45728
rect 158120 45664 158128 45728
rect 157808 44640 158128 45664
rect 157808 44576 157816 44640
rect 157880 44576 157896 44640
rect 157960 44576 157976 44640
rect 158040 44576 158056 44640
rect 158120 44576 158128 44640
rect 157808 43552 158128 44576
rect 157808 43488 157816 43552
rect 157880 43488 157896 43552
rect 157960 43488 157976 43552
rect 158040 43488 158056 43552
rect 158120 43488 158128 43552
rect 157808 42464 158128 43488
rect 157808 42400 157816 42464
rect 157880 42400 157896 42464
rect 157960 42400 157976 42464
rect 158040 42400 158056 42464
rect 158120 42400 158128 42464
rect 157808 41376 158128 42400
rect 157808 41312 157816 41376
rect 157880 41312 157896 41376
rect 157960 41312 157976 41376
rect 158040 41312 158056 41376
rect 158120 41312 158128 41376
rect 157808 40288 158128 41312
rect 157808 40224 157816 40288
rect 157880 40224 157896 40288
rect 157960 40224 157976 40288
rect 158040 40224 158056 40288
rect 158120 40224 158128 40288
rect 157808 39200 158128 40224
rect 157808 39136 157816 39200
rect 157880 39136 157896 39200
rect 157960 39136 157976 39200
rect 158040 39136 158056 39200
rect 158120 39136 158128 39200
rect 157808 38112 158128 39136
rect 157808 38048 157816 38112
rect 157880 38048 157896 38112
rect 157960 38048 157976 38112
rect 158040 38048 158056 38112
rect 158120 38048 158128 38112
rect 157808 37024 158128 38048
rect 157808 36960 157816 37024
rect 157880 36960 157896 37024
rect 157960 36960 157976 37024
rect 158040 36960 158056 37024
rect 158120 36960 158128 37024
rect 157808 35936 158128 36960
rect 157808 35872 157816 35936
rect 157880 35872 157896 35936
rect 157960 35872 157976 35936
rect 158040 35872 158056 35936
rect 158120 35872 158128 35936
rect 157808 34848 158128 35872
rect 157808 34784 157816 34848
rect 157880 34784 157896 34848
rect 157960 34784 157976 34848
rect 158040 34784 158056 34848
rect 158120 34784 158128 34848
rect 157808 33760 158128 34784
rect 157808 33696 157816 33760
rect 157880 33696 157896 33760
rect 157960 33696 157976 33760
rect 158040 33696 158056 33760
rect 158120 33696 158128 33760
rect 157808 32672 158128 33696
rect 157808 32608 157816 32672
rect 157880 32608 157896 32672
rect 157960 32608 157976 32672
rect 158040 32608 158056 32672
rect 158120 32608 158128 32672
rect 157808 31584 158128 32608
rect 157808 31520 157816 31584
rect 157880 31520 157896 31584
rect 157960 31520 157976 31584
rect 158040 31520 158056 31584
rect 158120 31520 158128 31584
rect 157808 30496 158128 31520
rect 157808 30432 157816 30496
rect 157880 30432 157896 30496
rect 157960 30432 157976 30496
rect 158040 30432 158056 30496
rect 158120 30432 158128 30496
rect 157808 29408 158128 30432
rect 157808 29344 157816 29408
rect 157880 29344 157896 29408
rect 157960 29344 157976 29408
rect 158040 29344 158056 29408
rect 158120 29344 158128 29408
rect 157808 28320 158128 29344
rect 157808 28256 157816 28320
rect 157880 28256 157896 28320
rect 157960 28256 157976 28320
rect 158040 28256 158056 28320
rect 158120 28256 158128 28320
rect 157808 27232 158128 28256
rect 157808 27168 157816 27232
rect 157880 27168 157896 27232
rect 157960 27168 157976 27232
rect 158040 27168 158056 27232
rect 158120 27168 158128 27232
rect 157808 26144 158128 27168
rect 157808 26080 157816 26144
rect 157880 26080 157896 26144
rect 157960 26080 157976 26144
rect 158040 26080 158056 26144
rect 158120 26080 158128 26144
rect 157808 25056 158128 26080
rect 157808 24992 157816 25056
rect 157880 24992 157896 25056
rect 157960 24992 157976 25056
rect 158040 24992 158056 25056
rect 158120 24992 158128 25056
rect 157808 23968 158128 24992
rect 157808 23904 157816 23968
rect 157880 23904 157896 23968
rect 157960 23904 157976 23968
rect 158040 23904 158056 23968
rect 158120 23904 158128 23968
rect 157808 22880 158128 23904
rect 157808 22816 157816 22880
rect 157880 22816 157896 22880
rect 157960 22816 157976 22880
rect 158040 22816 158056 22880
rect 158120 22816 158128 22880
rect 157808 21792 158128 22816
rect 157808 21728 157816 21792
rect 157880 21728 157896 21792
rect 157960 21728 157976 21792
rect 158040 21728 158056 21792
rect 158120 21728 158128 21792
rect 157808 20704 158128 21728
rect 157808 20640 157816 20704
rect 157880 20640 157896 20704
rect 157960 20640 157976 20704
rect 158040 20640 158056 20704
rect 158120 20640 158128 20704
rect 157808 19616 158128 20640
rect 157808 19552 157816 19616
rect 157880 19552 157896 19616
rect 157960 19552 157976 19616
rect 158040 19552 158056 19616
rect 158120 19552 158128 19616
rect 157808 18528 158128 19552
rect 157808 18464 157816 18528
rect 157880 18464 157896 18528
rect 157960 18464 157976 18528
rect 158040 18464 158056 18528
rect 158120 18464 158128 18528
rect 157808 17440 158128 18464
rect 157808 17376 157816 17440
rect 157880 17376 157896 17440
rect 157960 17376 157976 17440
rect 158040 17376 158056 17440
rect 158120 17376 158128 17440
rect 157808 16352 158128 17376
rect 157808 16288 157816 16352
rect 157880 16288 157896 16352
rect 157960 16288 157976 16352
rect 158040 16288 158056 16352
rect 158120 16288 158128 16352
rect 157808 15264 158128 16288
rect 157808 15200 157816 15264
rect 157880 15200 157896 15264
rect 157960 15200 157976 15264
rect 158040 15200 158056 15264
rect 158120 15200 158128 15264
rect 157808 14176 158128 15200
rect 157808 14112 157816 14176
rect 157880 14112 157896 14176
rect 157960 14112 157976 14176
rect 158040 14112 158056 14176
rect 158120 14112 158128 14176
rect 157808 13088 158128 14112
rect 157808 13024 157816 13088
rect 157880 13024 157896 13088
rect 157960 13024 157976 13088
rect 158040 13024 158056 13088
rect 158120 13024 158128 13088
rect 157808 12000 158128 13024
rect 157808 11936 157816 12000
rect 157880 11936 157896 12000
rect 157960 11936 157976 12000
rect 158040 11936 158056 12000
rect 158120 11936 158128 12000
rect 157808 10912 158128 11936
rect 157808 10848 157816 10912
rect 157880 10848 157896 10912
rect 157960 10848 157976 10912
rect 158040 10848 158056 10912
rect 158120 10848 158128 10912
rect 157808 9824 158128 10848
rect 157808 9760 157816 9824
rect 157880 9760 157896 9824
rect 157960 9760 157976 9824
rect 158040 9760 158056 9824
rect 158120 9760 158128 9824
rect 157808 8736 158128 9760
rect 157808 8672 157816 8736
rect 157880 8672 157896 8736
rect 157960 8672 157976 8736
rect 158040 8672 158056 8736
rect 158120 8672 158128 8736
rect 157808 7648 158128 8672
rect 157808 7584 157816 7648
rect 157880 7584 157896 7648
rect 157960 7584 157976 7648
rect 158040 7584 158056 7648
rect 158120 7584 158128 7648
rect 157808 6560 158128 7584
rect 157808 6496 157816 6560
rect 157880 6496 157896 6560
rect 157960 6496 157976 6560
rect 158040 6496 158056 6560
rect 158120 6496 158128 6560
rect 157808 5472 158128 6496
rect 157808 5408 157816 5472
rect 157880 5408 157896 5472
rect 157960 5408 157976 5472
rect 158040 5408 158056 5472
rect 158120 5408 158128 5472
rect 157808 4384 158128 5408
rect 157808 4320 157816 4384
rect 157880 4320 157896 4384
rect 157960 4320 157976 4384
rect 158040 4320 158056 4384
rect 158120 4320 158128 4384
rect 157808 3296 158128 4320
rect 157808 3232 157816 3296
rect 157880 3232 157896 3296
rect 157960 3232 157976 3296
rect 158040 3232 158056 3296
rect 158120 3232 158128 3296
rect 157808 2208 158128 3232
rect 157808 2144 157816 2208
rect 157880 2144 157896 2208
rect 157960 2144 157976 2208
rect 158040 2144 158056 2208
rect 158120 2144 158128 2208
rect 158468 2176 158788 117504
rect 159128 2176 159448 117504
rect 159788 2176 160108 117504
rect 173168 116992 173488 117552
rect 173168 116928 173176 116992
rect 173240 116928 173256 116992
rect 173320 116928 173336 116992
rect 173400 116928 173416 116992
rect 173480 116928 173488 116992
rect 173168 115904 173488 116928
rect 173168 115840 173176 115904
rect 173240 115840 173256 115904
rect 173320 115840 173336 115904
rect 173400 115840 173416 115904
rect 173480 115840 173488 115904
rect 173168 114816 173488 115840
rect 173168 114752 173176 114816
rect 173240 114752 173256 114816
rect 173320 114752 173336 114816
rect 173400 114752 173416 114816
rect 173480 114752 173488 114816
rect 173168 113728 173488 114752
rect 173168 113664 173176 113728
rect 173240 113664 173256 113728
rect 173320 113664 173336 113728
rect 173400 113664 173416 113728
rect 173480 113664 173488 113728
rect 173168 112640 173488 113664
rect 173168 112576 173176 112640
rect 173240 112576 173256 112640
rect 173320 112576 173336 112640
rect 173400 112576 173416 112640
rect 173480 112576 173488 112640
rect 173168 111552 173488 112576
rect 173168 111488 173176 111552
rect 173240 111488 173256 111552
rect 173320 111488 173336 111552
rect 173400 111488 173416 111552
rect 173480 111488 173488 111552
rect 173168 110464 173488 111488
rect 173168 110400 173176 110464
rect 173240 110400 173256 110464
rect 173320 110400 173336 110464
rect 173400 110400 173416 110464
rect 173480 110400 173488 110464
rect 173168 109376 173488 110400
rect 173168 109312 173176 109376
rect 173240 109312 173256 109376
rect 173320 109312 173336 109376
rect 173400 109312 173416 109376
rect 173480 109312 173488 109376
rect 173168 108288 173488 109312
rect 173168 108224 173176 108288
rect 173240 108224 173256 108288
rect 173320 108224 173336 108288
rect 173400 108224 173416 108288
rect 173480 108224 173488 108288
rect 173168 107200 173488 108224
rect 173168 107136 173176 107200
rect 173240 107136 173256 107200
rect 173320 107136 173336 107200
rect 173400 107136 173416 107200
rect 173480 107136 173488 107200
rect 173168 106112 173488 107136
rect 173168 106048 173176 106112
rect 173240 106048 173256 106112
rect 173320 106048 173336 106112
rect 173400 106048 173416 106112
rect 173480 106048 173488 106112
rect 173168 105024 173488 106048
rect 173168 104960 173176 105024
rect 173240 104960 173256 105024
rect 173320 104960 173336 105024
rect 173400 104960 173416 105024
rect 173480 104960 173488 105024
rect 173168 103936 173488 104960
rect 173168 103872 173176 103936
rect 173240 103872 173256 103936
rect 173320 103872 173336 103936
rect 173400 103872 173416 103936
rect 173480 103872 173488 103936
rect 173168 102848 173488 103872
rect 173168 102784 173176 102848
rect 173240 102784 173256 102848
rect 173320 102784 173336 102848
rect 173400 102784 173416 102848
rect 173480 102784 173488 102848
rect 173168 101760 173488 102784
rect 173168 101696 173176 101760
rect 173240 101696 173256 101760
rect 173320 101696 173336 101760
rect 173400 101696 173416 101760
rect 173480 101696 173488 101760
rect 173168 100672 173488 101696
rect 173168 100608 173176 100672
rect 173240 100608 173256 100672
rect 173320 100608 173336 100672
rect 173400 100608 173416 100672
rect 173480 100608 173488 100672
rect 173168 99584 173488 100608
rect 173168 99520 173176 99584
rect 173240 99520 173256 99584
rect 173320 99520 173336 99584
rect 173400 99520 173416 99584
rect 173480 99520 173488 99584
rect 173168 98496 173488 99520
rect 173168 98432 173176 98496
rect 173240 98432 173256 98496
rect 173320 98432 173336 98496
rect 173400 98432 173416 98496
rect 173480 98432 173488 98496
rect 173168 97408 173488 98432
rect 173168 97344 173176 97408
rect 173240 97344 173256 97408
rect 173320 97344 173336 97408
rect 173400 97344 173416 97408
rect 173480 97344 173488 97408
rect 173168 96320 173488 97344
rect 173168 96256 173176 96320
rect 173240 96256 173256 96320
rect 173320 96256 173336 96320
rect 173400 96256 173416 96320
rect 173480 96256 173488 96320
rect 173168 95232 173488 96256
rect 173168 95168 173176 95232
rect 173240 95168 173256 95232
rect 173320 95168 173336 95232
rect 173400 95168 173416 95232
rect 173480 95168 173488 95232
rect 173168 94144 173488 95168
rect 173168 94080 173176 94144
rect 173240 94080 173256 94144
rect 173320 94080 173336 94144
rect 173400 94080 173416 94144
rect 173480 94080 173488 94144
rect 173168 93056 173488 94080
rect 173168 92992 173176 93056
rect 173240 92992 173256 93056
rect 173320 92992 173336 93056
rect 173400 92992 173416 93056
rect 173480 92992 173488 93056
rect 173168 91968 173488 92992
rect 173168 91904 173176 91968
rect 173240 91904 173256 91968
rect 173320 91904 173336 91968
rect 173400 91904 173416 91968
rect 173480 91904 173488 91968
rect 173168 90880 173488 91904
rect 173168 90816 173176 90880
rect 173240 90816 173256 90880
rect 173320 90816 173336 90880
rect 173400 90816 173416 90880
rect 173480 90816 173488 90880
rect 173168 89792 173488 90816
rect 173168 89728 173176 89792
rect 173240 89728 173256 89792
rect 173320 89728 173336 89792
rect 173400 89728 173416 89792
rect 173480 89728 173488 89792
rect 173168 88704 173488 89728
rect 173168 88640 173176 88704
rect 173240 88640 173256 88704
rect 173320 88640 173336 88704
rect 173400 88640 173416 88704
rect 173480 88640 173488 88704
rect 173168 87616 173488 88640
rect 173168 87552 173176 87616
rect 173240 87552 173256 87616
rect 173320 87552 173336 87616
rect 173400 87552 173416 87616
rect 173480 87552 173488 87616
rect 173168 86528 173488 87552
rect 173168 86464 173176 86528
rect 173240 86464 173256 86528
rect 173320 86464 173336 86528
rect 173400 86464 173416 86528
rect 173480 86464 173488 86528
rect 173168 85440 173488 86464
rect 173168 85376 173176 85440
rect 173240 85376 173256 85440
rect 173320 85376 173336 85440
rect 173400 85376 173416 85440
rect 173480 85376 173488 85440
rect 173168 84352 173488 85376
rect 173168 84288 173176 84352
rect 173240 84288 173256 84352
rect 173320 84288 173336 84352
rect 173400 84288 173416 84352
rect 173480 84288 173488 84352
rect 173168 83264 173488 84288
rect 173168 83200 173176 83264
rect 173240 83200 173256 83264
rect 173320 83200 173336 83264
rect 173400 83200 173416 83264
rect 173480 83200 173488 83264
rect 173168 82176 173488 83200
rect 173168 82112 173176 82176
rect 173240 82112 173256 82176
rect 173320 82112 173336 82176
rect 173400 82112 173416 82176
rect 173480 82112 173488 82176
rect 173168 81088 173488 82112
rect 173168 81024 173176 81088
rect 173240 81024 173256 81088
rect 173320 81024 173336 81088
rect 173400 81024 173416 81088
rect 173480 81024 173488 81088
rect 173168 80000 173488 81024
rect 173168 79936 173176 80000
rect 173240 79936 173256 80000
rect 173320 79936 173336 80000
rect 173400 79936 173416 80000
rect 173480 79936 173488 80000
rect 173168 78912 173488 79936
rect 173168 78848 173176 78912
rect 173240 78848 173256 78912
rect 173320 78848 173336 78912
rect 173400 78848 173416 78912
rect 173480 78848 173488 78912
rect 173168 77824 173488 78848
rect 173168 77760 173176 77824
rect 173240 77760 173256 77824
rect 173320 77760 173336 77824
rect 173400 77760 173416 77824
rect 173480 77760 173488 77824
rect 173168 76736 173488 77760
rect 173168 76672 173176 76736
rect 173240 76672 173256 76736
rect 173320 76672 173336 76736
rect 173400 76672 173416 76736
rect 173480 76672 173488 76736
rect 173168 75648 173488 76672
rect 173168 75584 173176 75648
rect 173240 75584 173256 75648
rect 173320 75584 173336 75648
rect 173400 75584 173416 75648
rect 173480 75584 173488 75648
rect 173168 74560 173488 75584
rect 173168 74496 173176 74560
rect 173240 74496 173256 74560
rect 173320 74496 173336 74560
rect 173400 74496 173416 74560
rect 173480 74496 173488 74560
rect 173168 73472 173488 74496
rect 173168 73408 173176 73472
rect 173240 73408 173256 73472
rect 173320 73408 173336 73472
rect 173400 73408 173416 73472
rect 173480 73408 173488 73472
rect 173168 72384 173488 73408
rect 173168 72320 173176 72384
rect 173240 72320 173256 72384
rect 173320 72320 173336 72384
rect 173400 72320 173416 72384
rect 173480 72320 173488 72384
rect 173168 71296 173488 72320
rect 173168 71232 173176 71296
rect 173240 71232 173256 71296
rect 173320 71232 173336 71296
rect 173400 71232 173416 71296
rect 173480 71232 173488 71296
rect 173168 70208 173488 71232
rect 173168 70144 173176 70208
rect 173240 70144 173256 70208
rect 173320 70144 173336 70208
rect 173400 70144 173416 70208
rect 173480 70144 173488 70208
rect 173168 69120 173488 70144
rect 173168 69056 173176 69120
rect 173240 69056 173256 69120
rect 173320 69056 173336 69120
rect 173400 69056 173416 69120
rect 173480 69056 173488 69120
rect 173168 68032 173488 69056
rect 173168 67968 173176 68032
rect 173240 67968 173256 68032
rect 173320 67968 173336 68032
rect 173400 67968 173416 68032
rect 173480 67968 173488 68032
rect 173168 66944 173488 67968
rect 173168 66880 173176 66944
rect 173240 66880 173256 66944
rect 173320 66880 173336 66944
rect 173400 66880 173416 66944
rect 173480 66880 173488 66944
rect 173168 65856 173488 66880
rect 173168 65792 173176 65856
rect 173240 65792 173256 65856
rect 173320 65792 173336 65856
rect 173400 65792 173416 65856
rect 173480 65792 173488 65856
rect 173168 64768 173488 65792
rect 173168 64704 173176 64768
rect 173240 64704 173256 64768
rect 173320 64704 173336 64768
rect 173400 64704 173416 64768
rect 173480 64704 173488 64768
rect 173168 63680 173488 64704
rect 173168 63616 173176 63680
rect 173240 63616 173256 63680
rect 173320 63616 173336 63680
rect 173400 63616 173416 63680
rect 173480 63616 173488 63680
rect 173168 62592 173488 63616
rect 173168 62528 173176 62592
rect 173240 62528 173256 62592
rect 173320 62528 173336 62592
rect 173400 62528 173416 62592
rect 173480 62528 173488 62592
rect 173168 61504 173488 62528
rect 173168 61440 173176 61504
rect 173240 61440 173256 61504
rect 173320 61440 173336 61504
rect 173400 61440 173416 61504
rect 173480 61440 173488 61504
rect 173168 60416 173488 61440
rect 173168 60352 173176 60416
rect 173240 60352 173256 60416
rect 173320 60352 173336 60416
rect 173400 60352 173416 60416
rect 173480 60352 173488 60416
rect 173168 59328 173488 60352
rect 173168 59264 173176 59328
rect 173240 59264 173256 59328
rect 173320 59264 173336 59328
rect 173400 59264 173416 59328
rect 173480 59264 173488 59328
rect 173168 58240 173488 59264
rect 173168 58176 173176 58240
rect 173240 58176 173256 58240
rect 173320 58176 173336 58240
rect 173400 58176 173416 58240
rect 173480 58176 173488 58240
rect 173168 57152 173488 58176
rect 173168 57088 173176 57152
rect 173240 57088 173256 57152
rect 173320 57088 173336 57152
rect 173400 57088 173416 57152
rect 173480 57088 173488 57152
rect 173168 56064 173488 57088
rect 173168 56000 173176 56064
rect 173240 56000 173256 56064
rect 173320 56000 173336 56064
rect 173400 56000 173416 56064
rect 173480 56000 173488 56064
rect 173168 54976 173488 56000
rect 173168 54912 173176 54976
rect 173240 54912 173256 54976
rect 173320 54912 173336 54976
rect 173400 54912 173416 54976
rect 173480 54912 173488 54976
rect 173168 53888 173488 54912
rect 173168 53824 173176 53888
rect 173240 53824 173256 53888
rect 173320 53824 173336 53888
rect 173400 53824 173416 53888
rect 173480 53824 173488 53888
rect 173168 52800 173488 53824
rect 173168 52736 173176 52800
rect 173240 52736 173256 52800
rect 173320 52736 173336 52800
rect 173400 52736 173416 52800
rect 173480 52736 173488 52800
rect 173168 51712 173488 52736
rect 173168 51648 173176 51712
rect 173240 51648 173256 51712
rect 173320 51648 173336 51712
rect 173400 51648 173416 51712
rect 173480 51648 173488 51712
rect 173168 50624 173488 51648
rect 173168 50560 173176 50624
rect 173240 50560 173256 50624
rect 173320 50560 173336 50624
rect 173400 50560 173416 50624
rect 173480 50560 173488 50624
rect 173168 49536 173488 50560
rect 173168 49472 173176 49536
rect 173240 49472 173256 49536
rect 173320 49472 173336 49536
rect 173400 49472 173416 49536
rect 173480 49472 173488 49536
rect 173168 48448 173488 49472
rect 173168 48384 173176 48448
rect 173240 48384 173256 48448
rect 173320 48384 173336 48448
rect 173400 48384 173416 48448
rect 173480 48384 173488 48448
rect 173168 47360 173488 48384
rect 173168 47296 173176 47360
rect 173240 47296 173256 47360
rect 173320 47296 173336 47360
rect 173400 47296 173416 47360
rect 173480 47296 173488 47360
rect 173168 46272 173488 47296
rect 173168 46208 173176 46272
rect 173240 46208 173256 46272
rect 173320 46208 173336 46272
rect 173400 46208 173416 46272
rect 173480 46208 173488 46272
rect 173168 45184 173488 46208
rect 173168 45120 173176 45184
rect 173240 45120 173256 45184
rect 173320 45120 173336 45184
rect 173400 45120 173416 45184
rect 173480 45120 173488 45184
rect 173168 44096 173488 45120
rect 173168 44032 173176 44096
rect 173240 44032 173256 44096
rect 173320 44032 173336 44096
rect 173400 44032 173416 44096
rect 173480 44032 173488 44096
rect 173168 43008 173488 44032
rect 173168 42944 173176 43008
rect 173240 42944 173256 43008
rect 173320 42944 173336 43008
rect 173400 42944 173416 43008
rect 173480 42944 173488 43008
rect 173168 41920 173488 42944
rect 173168 41856 173176 41920
rect 173240 41856 173256 41920
rect 173320 41856 173336 41920
rect 173400 41856 173416 41920
rect 173480 41856 173488 41920
rect 173168 40832 173488 41856
rect 173168 40768 173176 40832
rect 173240 40768 173256 40832
rect 173320 40768 173336 40832
rect 173400 40768 173416 40832
rect 173480 40768 173488 40832
rect 173168 39744 173488 40768
rect 173168 39680 173176 39744
rect 173240 39680 173256 39744
rect 173320 39680 173336 39744
rect 173400 39680 173416 39744
rect 173480 39680 173488 39744
rect 173168 38656 173488 39680
rect 173168 38592 173176 38656
rect 173240 38592 173256 38656
rect 173320 38592 173336 38656
rect 173400 38592 173416 38656
rect 173480 38592 173488 38656
rect 173168 37568 173488 38592
rect 173168 37504 173176 37568
rect 173240 37504 173256 37568
rect 173320 37504 173336 37568
rect 173400 37504 173416 37568
rect 173480 37504 173488 37568
rect 173168 36480 173488 37504
rect 173168 36416 173176 36480
rect 173240 36416 173256 36480
rect 173320 36416 173336 36480
rect 173400 36416 173416 36480
rect 173480 36416 173488 36480
rect 173168 35392 173488 36416
rect 173168 35328 173176 35392
rect 173240 35328 173256 35392
rect 173320 35328 173336 35392
rect 173400 35328 173416 35392
rect 173480 35328 173488 35392
rect 173168 34304 173488 35328
rect 173168 34240 173176 34304
rect 173240 34240 173256 34304
rect 173320 34240 173336 34304
rect 173400 34240 173416 34304
rect 173480 34240 173488 34304
rect 173168 33216 173488 34240
rect 173168 33152 173176 33216
rect 173240 33152 173256 33216
rect 173320 33152 173336 33216
rect 173400 33152 173416 33216
rect 173480 33152 173488 33216
rect 173168 32128 173488 33152
rect 173168 32064 173176 32128
rect 173240 32064 173256 32128
rect 173320 32064 173336 32128
rect 173400 32064 173416 32128
rect 173480 32064 173488 32128
rect 173168 31040 173488 32064
rect 173168 30976 173176 31040
rect 173240 30976 173256 31040
rect 173320 30976 173336 31040
rect 173400 30976 173416 31040
rect 173480 30976 173488 31040
rect 173168 29952 173488 30976
rect 173168 29888 173176 29952
rect 173240 29888 173256 29952
rect 173320 29888 173336 29952
rect 173400 29888 173416 29952
rect 173480 29888 173488 29952
rect 173168 28864 173488 29888
rect 173168 28800 173176 28864
rect 173240 28800 173256 28864
rect 173320 28800 173336 28864
rect 173400 28800 173416 28864
rect 173480 28800 173488 28864
rect 173168 27776 173488 28800
rect 173168 27712 173176 27776
rect 173240 27712 173256 27776
rect 173320 27712 173336 27776
rect 173400 27712 173416 27776
rect 173480 27712 173488 27776
rect 173168 26688 173488 27712
rect 173168 26624 173176 26688
rect 173240 26624 173256 26688
rect 173320 26624 173336 26688
rect 173400 26624 173416 26688
rect 173480 26624 173488 26688
rect 173168 25600 173488 26624
rect 173168 25536 173176 25600
rect 173240 25536 173256 25600
rect 173320 25536 173336 25600
rect 173400 25536 173416 25600
rect 173480 25536 173488 25600
rect 173168 24512 173488 25536
rect 173168 24448 173176 24512
rect 173240 24448 173256 24512
rect 173320 24448 173336 24512
rect 173400 24448 173416 24512
rect 173480 24448 173488 24512
rect 173168 23424 173488 24448
rect 173168 23360 173176 23424
rect 173240 23360 173256 23424
rect 173320 23360 173336 23424
rect 173400 23360 173416 23424
rect 173480 23360 173488 23424
rect 173168 22336 173488 23360
rect 173168 22272 173176 22336
rect 173240 22272 173256 22336
rect 173320 22272 173336 22336
rect 173400 22272 173416 22336
rect 173480 22272 173488 22336
rect 173168 21248 173488 22272
rect 173168 21184 173176 21248
rect 173240 21184 173256 21248
rect 173320 21184 173336 21248
rect 173400 21184 173416 21248
rect 173480 21184 173488 21248
rect 173168 20160 173488 21184
rect 173168 20096 173176 20160
rect 173240 20096 173256 20160
rect 173320 20096 173336 20160
rect 173400 20096 173416 20160
rect 173480 20096 173488 20160
rect 173168 19072 173488 20096
rect 173168 19008 173176 19072
rect 173240 19008 173256 19072
rect 173320 19008 173336 19072
rect 173400 19008 173416 19072
rect 173480 19008 173488 19072
rect 173168 17984 173488 19008
rect 173168 17920 173176 17984
rect 173240 17920 173256 17984
rect 173320 17920 173336 17984
rect 173400 17920 173416 17984
rect 173480 17920 173488 17984
rect 173168 16896 173488 17920
rect 173168 16832 173176 16896
rect 173240 16832 173256 16896
rect 173320 16832 173336 16896
rect 173400 16832 173416 16896
rect 173480 16832 173488 16896
rect 173168 15808 173488 16832
rect 173168 15744 173176 15808
rect 173240 15744 173256 15808
rect 173320 15744 173336 15808
rect 173400 15744 173416 15808
rect 173480 15744 173488 15808
rect 173168 14720 173488 15744
rect 173168 14656 173176 14720
rect 173240 14656 173256 14720
rect 173320 14656 173336 14720
rect 173400 14656 173416 14720
rect 173480 14656 173488 14720
rect 173168 13632 173488 14656
rect 173168 13568 173176 13632
rect 173240 13568 173256 13632
rect 173320 13568 173336 13632
rect 173400 13568 173416 13632
rect 173480 13568 173488 13632
rect 173168 12544 173488 13568
rect 173168 12480 173176 12544
rect 173240 12480 173256 12544
rect 173320 12480 173336 12544
rect 173400 12480 173416 12544
rect 173480 12480 173488 12544
rect 173168 11456 173488 12480
rect 173168 11392 173176 11456
rect 173240 11392 173256 11456
rect 173320 11392 173336 11456
rect 173400 11392 173416 11456
rect 173480 11392 173488 11456
rect 173168 10368 173488 11392
rect 173168 10304 173176 10368
rect 173240 10304 173256 10368
rect 173320 10304 173336 10368
rect 173400 10304 173416 10368
rect 173480 10304 173488 10368
rect 173168 9280 173488 10304
rect 173168 9216 173176 9280
rect 173240 9216 173256 9280
rect 173320 9216 173336 9280
rect 173400 9216 173416 9280
rect 173480 9216 173488 9280
rect 173168 8192 173488 9216
rect 173168 8128 173176 8192
rect 173240 8128 173256 8192
rect 173320 8128 173336 8192
rect 173400 8128 173416 8192
rect 173480 8128 173488 8192
rect 173168 7104 173488 8128
rect 173168 7040 173176 7104
rect 173240 7040 173256 7104
rect 173320 7040 173336 7104
rect 173400 7040 173416 7104
rect 173480 7040 173488 7104
rect 173168 6016 173488 7040
rect 173168 5952 173176 6016
rect 173240 5952 173256 6016
rect 173320 5952 173336 6016
rect 173400 5952 173416 6016
rect 173480 5952 173488 6016
rect 173168 4928 173488 5952
rect 173168 4864 173176 4928
rect 173240 4864 173256 4928
rect 173320 4864 173336 4928
rect 173400 4864 173416 4928
rect 173480 4864 173488 4928
rect 173168 3840 173488 4864
rect 173168 3776 173176 3840
rect 173240 3776 173256 3840
rect 173320 3776 173336 3840
rect 173400 3776 173416 3840
rect 173480 3776 173488 3840
rect 173168 2752 173488 3776
rect 173168 2688 173176 2752
rect 173240 2688 173256 2752
rect 173320 2688 173336 2752
rect 173400 2688 173416 2752
rect 173480 2688 173488 2752
rect 157808 2128 158128 2144
rect 173168 2128 173488 2688
rect 173828 2176 174148 117504
rect 174488 2176 174808 117504
rect 175148 2176 175468 117504
rect 86723 2004 86789 2005
rect 86723 1940 86724 2004
rect 86788 1940 86789 2004
rect 86723 1939 86789 1940
<< via4 >>
rect 2550 3092 2786 3178
rect 2550 3028 2636 3092
rect 2636 3028 2700 3092
rect 2700 3028 2786 3092
rect 2550 2942 2786 3028
rect 102094 3092 102330 3178
rect 102094 3028 102180 3092
rect 102180 3028 102244 3092
rect 102244 3028 102330 3092
rect 102094 2942 102330 3028
<< metal5 >>
rect 2508 3178 102372 3220
rect 2508 2942 2550 3178
rect 2786 2942 102094 3178
rect 102330 2942 102372 3178
rect 2508 2900 102372 2942
<< labels >>
rlabel metal2 s 754 119200 810 120000 6 io_in[0]
port 0 nsew signal input
rlabel metal2 s 47674 119200 47730 120000 6 io_in[10]
port 1 nsew signal input
rlabel metal2 s 52366 119200 52422 120000 6 io_in[11]
port 2 nsew signal input
rlabel metal2 s 57058 119200 57114 120000 6 io_in[12]
port 3 nsew signal input
rlabel metal2 s 61750 119200 61806 120000 6 io_in[13]
port 4 nsew signal input
rlabel metal2 s 66442 119200 66498 120000 6 io_in[14]
port 5 nsew signal input
rlabel metal2 s 71134 119200 71190 120000 6 io_in[15]
port 6 nsew signal input
rlabel metal2 s 75826 119200 75882 120000 6 io_in[16]
port 7 nsew signal input
rlabel metal2 s 80518 119200 80574 120000 6 io_in[17]
port 8 nsew signal input
rlabel metal2 s 85210 119200 85266 120000 6 io_in[18]
port 9 nsew signal input
rlabel metal2 s 89902 119200 89958 120000 6 io_in[19]
port 10 nsew signal input
rlabel metal2 s 5446 119200 5502 120000 6 io_in[1]
port 11 nsew signal input
rlabel metal2 s 94686 119200 94742 120000 6 io_in[20]
port 12 nsew signal input
rlabel metal2 s 99378 119200 99434 120000 6 io_in[21]
port 13 nsew signal input
rlabel metal2 s 104070 119200 104126 120000 6 io_in[22]
port 14 nsew signal input
rlabel metal2 s 108762 119200 108818 120000 6 io_in[23]
port 15 nsew signal input
rlabel metal2 s 113454 119200 113510 120000 6 io_in[24]
port 16 nsew signal input
rlabel metal2 s 118146 119200 118202 120000 6 io_in[25]
port 17 nsew signal input
rlabel metal2 s 122838 119200 122894 120000 6 io_in[26]
port 18 nsew signal input
rlabel metal2 s 127530 119200 127586 120000 6 io_in[27]
port 19 nsew signal input
rlabel metal2 s 132222 119200 132278 120000 6 io_in[28]
port 20 nsew signal input
rlabel metal2 s 136914 119200 136970 120000 6 io_in[29]
port 21 nsew signal input
rlabel metal2 s 10138 119200 10194 120000 6 io_in[2]
port 22 nsew signal input
rlabel metal2 s 141606 119200 141662 120000 6 io_in[30]
port 23 nsew signal input
rlabel metal2 s 146298 119200 146354 120000 6 io_in[31]
port 24 nsew signal input
rlabel metal2 s 150990 119200 151046 120000 6 io_in[32]
port 25 nsew signal input
rlabel metal2 s 155682 119200 155738 120000 6 io_in[33]
port 26 nsew signal input
rlabel metal2 s 160374 119200 160430 120000 6 io_in[34]
port 27 nsew signal input
rlabel metal2 s 165066 119200 165122 120000 6 io_in[35]
port 28 nsew signal input
rlabel metal2 s 169758 119200 169814 120000 6 io_in[36]
port 29 nsew signal input
rlabel metal2 s 174450 119200 174506 120000 6 io_in[37]
port 30 nsew signal input
rlabel metal2 s 14830 119200 14886 120000 6 io_in[3]
port 31 nsew signal input
rlabel metal2 s 19522 119200 19578 120000 6 io_in[4]
port 32 nsew signal input
rlabel metal2 s 24214 119200 24270 120000 6 io_in[5]
port 33 nsew signal input
rlabel metal2 s 28906 119200 28962 120000 6 io_in[6]
port 34 nsew signal input
rlabel metal2 s 33598 119200 33654 120000 6 io_in[7]
port 35 nsew signal input
rlabel metal2 s 38290 119200 38346 120000 6 io_in[8]
port 36 nsew signal input
rlabel metal2 s 42982 119200 43038 120000 6 io_in[9]
port 37 nsew signal input
rlabel metal2 s 2318 119200 2374 120000 6 io_oeb[0]
port 38 nsew signal tristate
rlabel metal2 s 49238 119200 49294 120000 6 io_oeb[10]
port 39 nsew signal tristate
rlabel metal2 s 53930 119200 53986 120000 6 io_oeb[11]
port 40 nsew signal tristate
rlabel metal2 s 58622 119200 58678 120000 6 io_oeb[12]
port 41 nsew signal tristate
rlabel metal2 s 63314 119200 63370 120000 6 io_oeb[13]
port 42 nsew signal tristate
rlabel metal2 s 68006 119200 68062 120000 6 io_oeb[14]
port 43 nsew signal tristate
rlabel metal2 s 72698 119200 72754 120000 6 io_oeb[15]
port 44 nsew signal tristate
rlabel metal2 s 77390 119200 77446 120000 6 io_oeb[16]
port 45 nsew signal tristate
rlabel metal2 s 82082 119200 82138 120000 6 io_oeb[17]
port 46 nsew signal tristate
rlabel metal2 s 86774 119200 86830 120000 6 io_oeb[18]
port 47 nsew signal tristate
rlabel metal2 s 91558 119200 91614 120000 6 io_oeb[19]
port 48 nsew signal tristate
rlabel metal2 s 7010 119200 7066 120000 6 io_oeb[1]
port 49 nsew signal tristate
rlabel metal2 s 96250 119200 96306 120000 6 io_oeb[20]
port 50 nsew signal tristate
rlabel metal2 s 100942 119200 100998 120000 6 io_oeb[21]
port 51 nsew signal tristate
rlabel metal2 s 105634 119200 105690 120000 6 io_oeb[22]
port 52 nsew signal tristate
rlabel metal2 s 110326 119200 110382 120000 6 io_oeb[23]
port 53 nsew signal tristate
rlabel metal2 s 115018 119200 115074 120000 6 io_oeb[24]
port 54 nsew signal tristate
rlabel metal2 s 119710 119200 119766 120000 6 io_oeb[25]
port 55 nsew signal tristate
rlabel metal2 s 124402 119200 124458 120000 6 io_oeb[26]
port 56 nsew signal tristate
rlabel metal2 s 129094 119200 129150 120000 6 io_oeb[27]
port 57 nsew signal tristate
rlabel metal2 s 133786 119200 133842 120000 6 io_oeb[28]
port 58 nsew signal tristate
rlabel metal2 s 138478 119200 138534 120000 6 io_oeb[29]
port 59 nsew signal tristate
rlabel metal2 s 11702 119200 11758 120000 6 io_oeb[2]
port 60 nsew signal tristate
rlabel metal2 s 143170 119200 143226 120000 6 io_oeb[30]
port 61 nsew signal tristate
rlabel metal2 s 147862 119200 147918 120000 6 io_oeb[31]
port 62 nsew signal tristate
rlabel metal2 s 152554 119200 152610 120000 6 io_oeb[32]
port 63 nsew signal tristate
rlabel metal2 s 157246 119200 157302 120000 6 io_oeb[33]
port 64 nsew signal tristate
rlabel metal2 s 161938 119200 161994 120000 6 io_oeb[34]
port 65 nsew signal tristate
rlabel metal2 s 166630 119200 166686 120000 6 io_oeb[35]
port 66 nsew signal tristate
rlabel metal2 s 171322 119200 171378 120000 6 io_oeb[36]
port 67 nsew signal tristate
rlabel metal2 s 176014 119200 176070 120000 6 io_oeb[37]
port 68 nsew signal tristate
rlabel metal2 s 16394 119200 16450 120000 6 io_oeb[3]
port 69 nsew signal tristate
rlabel metal2 s 21086 119200 21142 120000 6 io_oeb[4]
port 70 nsew signal tristate
rlabel metal2 s 25778 119200 25834 120000 6 io_oeb[5]
port 71 nsew signal tristate
rlabel metal2 s 30470 119200 30526 120000 6 io_oeb[6]
port 72 nsew signal tristate
rlabel metal2 s 35162 119200 35218 120000 6 io_oeb[7]
port 73 nsew signal tristate
rlabel metal2 s 39854 119200 39910 120000 6 io_oeb[8]
port 74 nsew signal tristate
rlabel metal2 s 44546 119200 44602 120000 6 io_oeb[9]
port 75 nsew signal tristate
rlabel metal2 s 3882 119200 3938 120000 6 io_out[0]
port 76 nsew signal tristate
rlabel metal2 s 50802 119200 50858 120000 6 io_out[10]
port 77 nsew signal tristate
rlabel metal2 s 55494 119200 55550 120000 6 io_out[11]
port 78 nsew signal tristate
rlabel metal2 s 60186 119200 60242 120000 6 io_out[12]
port 79 nsew signal tristate
rlabel metal2 s 64878 119200 64934 120000 6 io_out[13]
port 80 nsew signal tristate
rlabel metal2 s 69570 119200 69626 120000 6 io_out[14]
port 81 nsew signal tristate
rlabel metal2 s 74262 119200 74318 120000 6 io_out[15]
port 82 nsew signal tristate
rlabel metal2 s 78954 119200 79010 120000 6 io_out[16]
port 83 nsew signal tristate
rlabel metal2 s 83646 119200 83702 120000 6 io_out[17]
port 84 nsew signal tristate
rlabel metal2 s 88338 119200 88394 120000 6 io_out[18]
port 85 nsew signal tristate
rlabel metal2 s 93122 119200 93178 120000 6 io_out[19]
port 86 nsew signal tristate
rlabel metal2 s 8574 119200 8630 120000 6 io_out[1]
port 87 nsew signal tristate
rlabel metal2 s 97814 119200 97870 120000 6 io_out[20]
port 88 nsew signal tristate
rlabel metal2 s 102506 119200 102562 120000 6 io_out[21]
port 89 nsew signal tristate
rlabel metal2 s 107198 119200 107254 120000 6 io_out[22]
port 90 nsew signal tristate
rlabel metal2 s 111890 119200 111946 120000 6 io_out[23]
port 91 nsew signal tristate
rlabel metal2 s 116582 119200 116638 120000 6 io_out[24]
port 92 nsew signal tristate
rlabel metal2 s 121274 119200 121330 120000 6 io_out[25]
port 93 nsew signal tristate
rlabel metal2 s 125966 119200 126022 120000 6 io_out[26]
port 94 nsew signal tristate
rlabel metal2 s 130658 119200 130714 120000 6 io_out[27]
port 95 nsew signal tristate
rlabel metal2 s 135350 119200 135406 120000 6 io_out[28]
port 96 nsew signal tristate
rlabel metal2 s 140042 119200 140098 120000 6 io_out[29]
port 97 nsew signal tristate
rlabel metal2 s 13266 119200 13322 120000 6 io_out[2]
port 98 nsew signal tristate
rlabel metal2 s 144734 119200 144790 120000 6 io_out[30]
port 99 nsew signal tristate
rlabel metal2 s 149426 119200 149482 120000 6 io_out[31]
port 100 nsew signal tristate
rlabel metal2 s 154118 119200 154174 120000 6 io_out[32]
port 101 nsew signal tristate
rlabel metal2 s 158810 119200 158866 120000 6 io_out[33]
port 102 nsew signal tristate
rlabel metal2 s 163502 119200 163558 120000 6 io_out[34]
port 103 nsew signal tristate
rlabel metal2 s 168194 119200 168250 120000 6 io_out[35]
port 104 nsew signal tristate
rlabel metal2 s 172886 119200 172942 120000 6 io_out[36]
port 105 nsew signal tristate
rlabel metal2 s 177578 119200 177634 120000 6 io_out[37]
port 106 nsew signal tristate
rlabel metal2 s 17958 119200 18014 120000 6 io_out[3]
port 107 nsew signal tristate
rlabel metal2 s 22650 119200 22706 120000 6 io_out[4]
port 108 nsew signal tristate
rlabel metal2 s 27342 119200 27398 120000 6 io_out[5]
port 109 nsew signal tristate
rlabel metal2 s 32034 119200 32090 120000 6 io_out[6]
port 110 nsew signal tristate
rlabel metal2 s 36726 119200 36782 120000 6 io_out[7]
port 111 nsew signal tristate
rlabel metal2 s 41418 119200 41474 120000 6 io_out[8]
port 112 nsew signal tristate
rlabel metal2 s 46110 119200 46166 120000 6 io_out[9]
port 113 nsew signal tristate
rlabel metal3 s 179200 59984 180000 60104 6 irq[0]
port 114 nsew signal tristate
rlabel metal3 s 0 59984 800 60104 6 irq[1]
port 115 nsew signal tristate
rlabel metal2 s 179142 119200 179198 120000 6 irq[2]
port 116 nsew signal tristate
rlabel metal2 s 39026 0 39082 800 6 la_data_in[0]
port 117 nsew signal input
rlabel metal2 s 149242 0 149298 800 6 la_data_in[100]
port 118 nsew signal input
rlabel metal2 s 150346 0 150402 800 6 la_data_in[101]
port 119 nsew signal input
rlabel metal2 s 151450 0 151506 800 6 la_data_in[102]
port 120 nsew signal input
rlabel metal2 s 152554 0 152610 800 6 la_data_in[103]
port 121 nsew signal input
rlabel metal2 s 153658 0 153714 800 6 la_data_in[104]
port 122 nsew signal input
rlabel metal2 s 154762 0 154818 800 6 la_data_in[105]
port 123 nsew signal input
rlabel metal2 s 155866 0 155922 800 6 la_data_in[106]
port 124 nsew signal input
rlabel metal2 s 156970 0 157026 800 6 la_data_in[107]
port 125 nsew signal input
rlabel metal2 s 158074 0 158130 800 6 la_data_in[108]
port 126 nsew signal input
rlabel metal2 s 159178 0 159234 800 6 la_data_in[109]
port 127 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 la_data_in[10]
port 128 nsew signal input
rlabel metal2 s 160282 0 160338 800 6 la_data_in[110]
port 129 nsew signal input
rlabel metal2 s 161386 0 161442 800 6 la_data_in[111]
port 130 nsew signal input
rlabel metal2 s 162490 0 162546 800 6 la_data_in[112]
port 131 nsew signal input
rlabel metal2 s 163594 0 163650 800 6 la_data_in[113]
port 132 nsew signal input
rlabel metal2 s 164698 0 164754 800 6 la_data_in[114]
port 133 nsew signal input
rlabel metal2 s 165802 0 165858 800 6 la_data_in[115]
port 134 nsew signal input
rlabel metal2 s 166906 0 166962 800 6 la_data_in[116]
port 135 nsew signal input
rlabel metal2 s 168010 0 168066 800 6 la_data_in[117]
port 136 nsew signal input
rlabel metal2 s 169114 0 169170 800 6 la_data_in[118]
port 137 nsew signal input
rlabel metal2 s 170218 0 170274 800 6 la_data_in[119]
port 138 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 la_data_in[11]
port 139 nsew signal input
rlabel metal2 s 171322 0 171378 800 6 la_data_in[120]
port 140 nsew signal input
rlabel metal2 s 172426 0 172482 800 6 la_data_in[121]
port 141 nsew signal input
rlabel metal2 s 173530 0 173586 800 6 la_data_in[122]
port 142 nsew signal input
rlabel metal2 s 174634 0 174690 800 6 la_data_in[123]
port 143 nsew signal input
rlabel metal2 s 175738 0 175794 800 6 la_data_in[124]
port 144 nsew signal input
rlabel metal2 s 176842 0 176898 800 6 la_data_in[125]
port 145 nsew signal input
rlabel metal2 s 177946 0 178002 800 6 la_data_in[126]
port 146 nsew signal input
rlabel metal2 s 179050 0 179106 800 6 la_data_in[127]
port 147 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 la_data_in[12]
port 148 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 la_data_in[13]
port 149 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 la_data_in[14]
port 150 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 la_data_in[15]
port 151 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 la_data_in[16]
port 152 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 la_data_in[17]
port 153 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 la_data_in[18]
port 154 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 la_data_in[19]
port 155 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 la_data_in[1]
port 156 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 la_data_in[20]
port 157 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 la_data_in[21]
port 158 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 la_data_in[22]
port 159 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 la_data_in[23]
port 160 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_data_in[24]
port 161 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_data_in[25]
port 162 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_data_in[26]
port 163 nsew signal input
rlabel metal2 s 68742 0 68798 800 6 la_data_in[27]
port 164 nsew signal input
rlabel metal2 s 69846 0 69902 800 6 la_data_in[28]
port 165 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 la_data_in[29]
port 166 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 la_data_in[2]
port 167 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_data_in[30]
port 168 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 la_data_in[31]
port 169 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 la_data_in[32]
port 170 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 la_data_in[33]
port 171 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 la_data_in[34]
port 172 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 la_data_in[35]
port 173 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 la_data_in[36]
port 174 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 la_data_in[37]
port 175 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 la_data_in[38]
port 176 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_data_in[39]
port 177 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 la_data_in[3]
port 178 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 la_data_in[40]
port 179 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 la_data_in[41]
port 180 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 la_data_in[42]
port 181 nsew signal input
rlabel metal2 s 86406 0 86462 800 6 la_data_in[43]
port 182 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_data_in[44]
port 183 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 la_data_in[45]
port 184 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_data_in[46]
port 185 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 la_data_in[47]
port 186 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 la_data_in[48]
port 187 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 la_data_in[49]
port 188 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 la_data_in[4]
port 189 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 la_data_in[50]
port 190 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 la_data_in[51]
port 191 nsew signal input
rlabel metal2 s 96342 0 96398 800 6 la_data_in[52]
port 192 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_data_in[53]
port 193 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 la_data_in[54]
port 194 nsew signal input
rlabel metal2 s 99654 0 99710 800 6 la_data_in[55]
port 195 nsew signal input
rlabel metal2 s 100758 0 100814 800 6 la_data_in[56]
port 196 nsew signal input
rlabel metal2 s 101862 0 101918 800 6 la_data_in[57]
port 197 nsew signal input
rlabel metal2 s 102966 0 103022 800 6 la_data_in[58]
port 198 nsew signal input
rlabel metal2 s 104070 0 104126 800 6 la_data_in[59]
port 199 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 la_data_in[5]
port 200 nsew signal input
rlabel metal2 s 105174 0 105230 800 6 la_data_in[60]
port 201 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 la_data_in[61]
port 202 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 la_data_in[62]
port 203 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 la_data_in[63]
port 204 nsew signal input
rlabel metal2 s 109590 0 109646 800 6 la_data_in[64]
port 205 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 la_data_in[65]
port 206 nsew signal input
rlabel metal2 s 111798 0 111854 800 6 la_data_in[66]
port 207 nsew signal input
rlabel metal2 s 112902 0 112958 800 6 la_data_in[67]
port 208 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 la_data_in[68]
port 209 nsew signal input
rlabel metal2 s 115110 0 115166 800 6 la_data_in[69]
port 210 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 la_data_in[6]
port 211 nsew signal input
rlabel metal2 s 116214 0 116270 800 6 la_data_in[70]
port 212 nsew signal input
rlabel metal2 s 117318 0 117374 800 6 la_data_in[71]
port 213 nsew signal input
rlabel metal2 s 118422 0 118478 800 6 la_data_in[72]
port 214 nsew signal input
rlabel metal2 s 119526 0 119582 800 6 la_data_in[73]
port 215 nsew signal input
rlabel metal2 s 120538 0 120594 800 6 la_data_in[74]
port 216 nsew signal input
rlabel metal2 s 121642 0 121698 800 6 la_data_in[75]
port 217 nsew signal input
rlabel metal2 s 122746 0 122802 800 6 la_data_in[76]
port 218 nsew signal input
rlabel metal2 s 123850 0 123906 800 6 la_data_in[77]
port 219 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 la_data_in[78]
port 220 nsew signal input
rlabel metal2 s 126058 0 126114 800 6 la_data_in[79]
port 221 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 la_data_in[7]
port 222 nsew signal input
rlabel metal2 s 127162 0 127218 800 6 la_data_in[80]
port 223 nsew signal input
rlabel metal2 s 128266 0 128322 800 6 la_data_in[81]
port 224 nsew signal input
rlabel metal2 s 129370 0 129426 800 6 la_data_in[82]
port 225 nsew signal input
rlabel metal2 s 130474 0 130530 800 6 la_data_in[83]
port 226 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 la_data_in[84]
port 227 nsew signal input
rlabel metal2 s 132682 0 132738 800 6 la_data_in[85]
port 228 nsew signal input
rlabel metal2 s 133786 0 133842 800 6 la_data_in[86]
port 229 nsew signal input
rlabel metal2 s 134890 0 134946 800 6 la_data_in[87]
port 230 nsew signal input
rlabel metal2 s 135994 0 136050 800 6 la_data_in[88]
port 231 nsew signal input
rlabel metal2 s 137098 0 137154 800 6 la_data_in[89]
port 232 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 la_data_in[8]
port 233 nsew signal input
rlabel metal2 s 138202 0 138258 800 6 la_data_in[90]
port 234 nsew signal input
rlabel metal2 s 139306 0 139362 800 6 la_data_in[91]
port 235 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 la_data_in[92]
port 236 nsew signal input
rlabel metal2 s 141514 0 141570 800 6 la_data_in[93]
port 237 nsew signal input
rlabel metal2 s 142618 0 142674 800 6 la_data_in[94]
port 238 nsew signal input
rlabel metal2 s 143722 0 143778 800 6 la_data_in[95]
port 239 nsew signal input
rlabel metal2 s 144826 0 144882 800 6 la_data_in[96]
port 240 nsew signal input
rlabel metal2 s 145930 0 145986 800 6 la_data_in[97]
port 241 nsew signal input
rlabel metal2 s 147034 0 147090 800 6 la_data_in[98]
port 242 nsew signal input
rlabel metal2 s 148138 0 148194 800 6 la_data_in[99]
port 243 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 la_data_in[9]
port 244 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 la_data_out[0]
port 245 nsew signal tristate
rlabel metal2 s 149610 0 149666 800 6 la_data_out[100]
port 246 nsew signal tristate
rlabel metal2 s 150714 0 150770 800 6 la_data_out[101]
port 247 nsew signal tristate
rlabel metal2 s 151818 0 151874 800 6 la_data_out[102]
port 248 nsew signal tristate
rlabel metal2 s 152922 0 152978 800 6 la_data_out[103]
port 249 nsew signal tristate
rlabel metal2 s 154026 0 154082 800 6 la_data_out[104]
port 250 nsew signal tristate
rlabel metal2 s 155130 0 155186 800 6 la_data_out[105]
port 251 nsew signal tristate
rlabel metal2 s 156234 0 156290 800 6 la_data_out[106]
port 252 nsew signal tristate
rlabel metal2 s 157338 0 157394 800 6 la_data_out[107]
port 253 nsew signal tristate
rlabel metal2 s 158442 0 158498 800 6 la_data_out[108]
port 254 nsew signal tristate
rlabel metal2 s 159546 0 159602 800 6 la_data_out[109]
port 255 nsew signal tristate
rlabel metal2 s 50434 0 50490 800 6 la_data_out[10]
port 256 nsew signal tristate
rlabel metal2 s 160650 0 160706 800 6 la_data_out[110]
port 257 nsew signal tristate
rlabel metal2 s 161754 0 161810 800 6 la_data_out[111]
port 258 nsew signal tristate
rlabel metal2 s 162858 0 162914 800 6 la_data_out[112]
port 259 nsew signal tristate
rlabel metal2 s 163962 0 164018 800 6 la_data_out[113]
port 260 nsew signal tristate
rlabel metal2 s 165066 0 165122 800 6 la_data_out[114]
port 261 nsew signal tristate
rlabel metal2 s 166170 0 166226 800 6 la_data_out[115]
port 262 nsew signal tristate
rlabel metal2 s 167274 0 167330 800 6 la_data_out[116]
port 263 nsew signal tristate
rlabel metal2 s 168378 0 168434 800 6 la_data_out[117]
port 264 nsew signal tristate
rlabel metal2 s 169482 0 169538 800 6 la_data_out[118]
port 265 nsew signal tristate
rlabel metal2 s 170586 0 170642 800 6 la_data_out[119]
port 266 nsew signal tristate
rlabel metal2 s 51538 0 51594 800 6 la_data_out[11]
port 267 nsew signal tristate
rlabel metal2 s 171690 0 171746 800 6 la_data_out[120]
port 268 nsew signal tristate
rlabel metal2 s 172794 0 172850 800 6 la_data_out[121]
port 269 nsew signal tristate
rlabel metal2 s 173898 0 173954 800 6 la_data_out[122]
port 270 nsew signal tristate
rlabel metal2 s 175002 0 175058 800 6 la_data_out[123]
port 271 nsew signal tristate
rlabel metal2 s 176106 0 176162 800 6 la_data_out[124]
port 272 nsew signal tristate
rlabel metal2 s 177210 0 177266 800 6 la_data_out[125]
port 273 nsew signal tristate
rlabel metal2 s 178314 0 178370 800 6 la_data_out[126]
port 274 nsew signal tristate
rlabel metal2 s 179418 0 179474 800 6 la_data_out[127]
port 275 nsew signal tristate
rlabel metal2 s 52642 0 52698 800 6 la_data_out[12]
port 276 nsew signal tristate
rlabel metal2 s 53746 0 53802 800 6 la_data_out[13]
port 277 nsew signal tristate
rlabel metal2 s 54850 0 54906 800 6 la_data_out[14]
port 278 nsew signal tristate
rlabel metal2 s 55954 0 56010 800 6 la_data_out[15]
port 279 nsew signal tristate
rlabel metal2 s 57058 0 57114 800 6 la_data_out[16]
port 280 nsew signal tristate
rlabel metal2 s 58162 0 58218 800 6 la_data_out[17]
port 281 nsew signal tristate
rlabel metal2 s 59266 0 59322 800 6 la_data_out[18]
port 282 nsew signal tristate
rlabel metal2 s 60278 0 60334 800 6 la_data_out[19]
port 283 nsew signal tristate
rlabel metal2 s 40498 0 40554 800 6 la_data_out[1]
port 284 nsew signal tristate
rlabel metal2 s 61382 0 61438 800 6 la_data_out[20]
port 285 nsew signal tristate
rlabel metal2 s 62486 0 62542 800 6 la_data_out[21]
port 286 nsew signal tristate
rlabel metal2 s 63590 0 63646 800 6 la_data_out[22]
port 287 nsew signal tristate
rlabel metal2 s 64694 0 64750 800 6 la_data_out[23]
port 288 nsew signal tristate
rlabel metal2 s 65798 0 65854 800 6 la_data_out[24]
port 289 nsew signal tristate
rlabel metal2 s 66902 0 66958 800 6 la_data_out[25]
port 290 nsew signal tristate
rlabel metal2 s 68006 0 68062 800 6 la_data_out[26]
port 291 nsew signal tristate
rlabel metal2 s 69110 0 69166 800 6 la_data_out[27]
port 292 nsew signal tristate
rlabel metal2 s 70214 0 70270 800 6 la_data_out[28]
port 293 nsew signal tristate
rlabel metal2 s 71318 0 71374 800 6 la_data_out[29]
port 294 nsew signal tristate
rlabel metal2 s 41602 0 41658 800 6 la_data_out[2]
port 295 nsew signal tristate
rlabel metal2 s 72422 0 72478 800 6 la_data_out[30]
port 296 nsew signal tristate
rlabel metal2 s 73526 0 73582 800 6 la_data_out[31]
port 297 nsew signal tristate
rlabel metal2 s 74630 0 74686 800 6 la_data_out[32]
port 298 nsew signal tristate
rlabel metal2 s 75734 0 75790 800 6 la_data_out[33]
port 299 nsew signal tristate
rlabel metal2 s 76838 0 76894 800 6 la_data_out[34]
port 300 nsew signal tristate
rlabel metal2 s 77942 0 77998 800 6 la_data_out[35]
port 301 nsew signal tristate
rlabel metal2 s 79046 0 79102 800 6 la_data_out[36]
port 302 nsew signal tristate
rlabel metal2 s 80150 0 80206 800 6 la_data_out[37]
port 303 nsew signal tristate
rlabel metal2 s 81254 0 81310 800 6 la_data_out[38]
port 304 nsew signal tristate
rlabel metal2 s 82358 0 82414 800 6 la_data_out[39]
port 305 nsew signal tristate
rlabel metal2 s 42706 0 42762 800 6 la_data_out[3]
port 306 nsew signal tristate
rlabel metal2 s 83462 0 83518 800 6 la_data_out[40]
port 307 nsew signal tristate
rlabel metal2 s 84566 0 84622 800 6 la_data_out[41]
port 308 nsew signal tristate
rlabel metal2 s 85670 0 85726 800 6 la_data_out[42]
port 309 nsew signal tristate
rlabel metal2 s 86774 0 86830 800 6 la_data_out[43]
port 310 nsew signal tristate
rlabel metal2 s 87878 0 87934 800 6 la_data_out[44]
port 311 nsew signal tristate
rlabel metal2 s 88982 0 89038 800 6 la_data_out[45]
port 312 nsew signal tristate
rlabel metal2 s 90086 0 90142 800 6 la_data_out[46]
port 313 nsew signal tristate
rlabel metal2 s 91190 0 91246 800 6 la_data_out[47]
port 314 nsew signal tristate
rlabel metal2 s 92294 0 92350 800 6 la_data_out[48]
port 315 nsew signal tristate
rlabel metal2 s 93398 0 93454 800 6 la_data_out[49]
port 316 nsew signal tristate
rlabel metal2 s 43810 0 43866 800 6 la_data_out[4]
port 317 nsew signal tristate
rlabel metal2 s 94502 0 94558 800 6 la_data_out[50]
port 318 nsew signal tristate
rlabel metal2 s 95606 0 95662 800 6 la_data_out[51]
port 319 nsew signal tristate
rlabel metal2 s 96710 0 96766 800 6 la_data_out[52]
port 320 nsew signal tristate
rlabel metal2 s 97814 0 97870 800 6 la_data_out[53]
port 321 nsew signal tristate
rlabel metal2 s 98918 0 98974 800 6 la_data_out[54]
port 322 nsew signal tristate
rlabel metal2 s 100022 0 100078 800 6 la_data_out[55]
port 323 nsew signal tristate
rlabel metal2 s 101126 0 101182 800 6 la_data_out[56]
port 324 nsew signal tristate
rlabel metal2 s 102230 0 102286 800 6 la_data_out[57]
port 325 nsew signal tristate
rlabel metal2 s 103334 0 103390 800 6 la_data_out[58]
port 326 nsew signal tristate
rlabel metal2 s 104438 0 104494 800 6 la_data_out[59]
port 327 nsew signal tristate
rlabel metal2 s 44914 0 44970 800 6 la_data_out[5]
port 328 nsew signal tristate
rlabel metal2 s 105542 0 105598 800 6 la_data_out[60]
port 329 nsew signal tristate
rlabel metal2 s 106646 0 106702 800 6 la_data_out[61]
port 330 nsew signal tristate
rlabel metal2 s 107750 0 107806 800 6 la_data_out[62]
port 331 nsew signal tristate
rlabel metal2 s 108854 0 108910 800 6 la_data_out[63]
port 332 nsew signal tristate
rlabel metal2 s 109958 0 110014 800 6 la_data_out[64]
port 333 nsew signal tristate
rlabel metal2 s 111062 0 111118 800 6 la_data_out[65]
port 334 nsew signal tristate
rlabel metal2 s 112166 0 112222 800 6 la_data_out[66]
port 335 nsew signal tristate
rlabel metal2 s 113270 0 113326 800 6 la_data_out[67]
port 336 nsew signal tristate
rlabel metal2 s 114374 0 114430 800 6 la_data_out[68]
port 337 nsew signal tristate
rlabel metal2 s 115478 0 115534 800 6 la_data_out[69]
port 338 nsew signal tristate
rlabel metal2 s 46018 0 46074 800 6 la_data_out[6]
port 339 nsew signal tristate
rlabel metal2 s 116582 0 116638 800 6 la_data_out[70]
port 340 nsew signal tristate
rlabel metal2 s 117686 0 117742 800 6 la_data_out[71]
port 341 nsew signal tristate
rlabel metal2 s 118790 0 118846 800 6 la_data_out[72]
port 342 nsew signal tristate
rlabel metal2 s 119894 0 119950 800 6 la_data_out[73]
port 343 nsew signal tristate
rlabel metal2 s 120906 0 120962 800 6 la_data_out[74]
port 344 nsew signal tristate
rlabel metal2 s 122010 0 122066 800 6 la_data_out[75]
port 345 nsew signal tristate
rlabel metal2 s 123114 0 123170 800 6 la_data_out[76]
port 346 nsew signal tristate
rlabel metal2 s 124218 0 124274 800 6 la_data_out[77]
port 347 nsew signal tristate
rlabel metal2 s 125322 0 125378 800 6 la_data_out[78]
port 348 nsew signal tristate
rlabel metal2 s 126426 0 126482 800 6 la_data_out[79]
port 349 nsew signal tristate
rlabel metal2 s 47122 0 47178 800 6 la_data_out[7]
port 350 nsew signal tristate
rlabel metal2 s 127530 0 127586 800 6 la_data_out[80]
port 351 nsew signal tristate
rlabel metal2 s 128634 0 128690 800 6 la_data_out[81]
port 352 nsew signal tristate
rlabel metal2 s 129738 0 129794 800 6 la_data_out[82]
port 353 nsew signal tristate
rlabel metal2 s 130842 0 130898 800 6 la_data_out[83]
port 354 nsew signal tristate
rlabel metal2 s 131946 0 132002 800 6 la_data_out[84]
port 355 nsew signal tristate
rlabel metal2 s 133050 0 133106 800 6 la_data_out[85]
port 356 nsew signal tristate
rlabel metal2 s 134154 0 134210 800 6 la_data_out[86]
port 357 nsew signal tristate
rlabel metal2 s 135258 0 135314 800 6 la_data_out[87]
port 358 nsew signal tristate
rlabel metal2 s 136362 0 136418 800 6 la_data_out[88]
port 359 nsew signal tristate
rlabel metal2 s 137466 0 137522 800 6 la_data_out[89]
port 360 nsew signal tristate
rlabel metal2 s 48226 0 48282 800 6 la_data_out[8]
port 361 nsew signal tristate
rlabel metal2 s 138570 0 138626 800 6 la_data_out[90]
port 362 nsew signal tristate
rlabel metal2 s 139674 0 139730 800 6 la_data_out[91]
port 363 nsew signal tristate
rlabel metal2 s 140778 0 140834 800 6 la_data_out[92]
port 364 nsew signal tristate
rlabel metal2 s 141882 0 141938 800 6 la_data_out[93]
port 365 nsew signal tristate
rlabel metal2 s 142986 0 143042 800 6 la_data_out[94]
port 366 nsew signal tristate
rlabel metal2 s 144090 0 144146 800 6 la_data_out[95]
port 367 nsew signal tristate
rlabel metal2 s 145194 0 145250 800 6 la_data_out[96]
port 368 nsew signal tristate
rlabel metal2 s 146298 0 146354 800 6 la_data_out[97]
port 369 nsew signal tristate
rlabel metal2 s 147402 0 147458 800 6 la_data_out[98]
port 370 nsew signal tristate
rlabel metal2 s 148506 0 148562 800 6 la_data_out[99]
port 371 nsew signal tristate
rlabel metal2 s 49330 0 49386 800 6 la_data_out[9]
port 372 nsew signal tristate
rlabel metal2 s 39762 0 39818 800 6 la_oenb[0]
port 373 nsew signal input
rlabel metal2 s 149978 0 150034 800 6 la_oenb[100]
port 374 nsew signal input
rlabel metal2 s 151082 0 151138 800 6 la_oenb[101]
port 375 nsew signal input
rlabel metal2 s 152186 0 152242 800 6 la_oenb[102]
port 376 nsew signal input
rlabel metal2 s 153290 0 153346 800 6 la_oenb[103]
port 377 nsew signal input
rlabel metal2 s 154394 0 154450 800 6 la_oenb[104]
port 378 nsew signal input
rlabel metal2 s 155498 0 155554 800 6 la_oenb[105]
port 379 nsew signal input
rlabel metal2 s 156602 0 156658 800 6 la_oenb[106]
port 380 nsew signal input
rlabel metal2 s 157706 0 157762 800 6 la_oenb[107]
port 381 nsew signal input
rlabel metal2 s 158810 0 158866 800 6 la_oenb[108]
port 382 nsew signal input
rlabel metal2 s 159914 0 159970 800 6 la_oenb[109]
port 383 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 la_oenb[10]
port 384 nsew signal input
rlabel metal2 s 161018 0 161074 800 6 la_oenb[110]
port 385 nsew signal input
rlabel metal2 s 162122 0 162178 800 6 la_oenb[111]
port 386 nsew signal input
rlabel metal2 s 163226 0 163282 800 6 la_oenb[112]
port 387 nsew signal input
rlabel metal2 s 164330 0 164386 800 6 la_oenb[113]
port 388 nsew signal input
rlabel metal2 s 165434 0 165490 800 6 la_oenb[114]
port 389 nsew signal input
rlabel metal2 s 166538 0 166594 800 6 la_oenb[115]
port 390 nsew signal input
rlabel metal2 s 167642 0 167698 800 6 la_oenb[116]
port 391 nsew signal input
rlabel metal2 s 168746 0 168802 800 6 la_oenb[117]
port 392 nsew signal input
rlabel metal2 s 169850 0 169906 800 6 la_oenb[118]
port 393 nsew signal input
rlabel metal2 s 170954 0 171010 800 6 la_oenb[119]
port 394 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 la_oenb[11]
port 395 nsew signal input
rlabel metal2 s 172058 0 172114 800 6 la_oenb[120]
port 396 nsew signal input
rlabel metal2 s 173162 0 173218 800 6 la_oenb[121]
port 397 nsew signal input
rlabel metal2 s 174266 0 174322 800 6 la_oenb[122]
port 398 nsew signal input
rlabel metal2 s 175370 0 175426 800 6 la_oenb[123]
port 399 nsew signal input
rlabel metal2 s 176474 0 176530 800 6 la_oenb[124]
port 400 nsew signal input
rlabel metal2 s 177578 0 177634 800 6 la_oenb[125]
port 401 nsew signal input
rlabel metal2 s 178682 0 178738 800 6 la_oenb[126]
port 402 nsew signal input
rlabel metal2 s 179786 0 179842 800 6 la_oenb[127]
port 403 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 la_oenb[12]
port 404 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 la_oenb[13]
port 405 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 la_oenb[14]
port 406 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 la_oenb[15]
port 407 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 la_oenb[16]
port 408 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 la_oenb[17]
port 409 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 la_oenb[18]
port 410 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 la_oenb[19]
port 411 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 la_oenb[1]
port 412 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 la_oenb[20]
port 413 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_oenb[21]
port 414 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 la_oenb[22]
port 415 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 la_oenb[23]
port 416 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 la_oenb[24]
port 417 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 la_oenb[25]
port 418 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_oenb[26]
port 419 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 la_oenb[27]
port 420 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 la_oenb[28]
port 421 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 la_oenb[29]
port 422 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 la_oenb[2]
port 423 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 la_oenb[30]
port 424 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 la_oenb[31]
port 425 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_oenb[32]
port 426 nsew signal input
rlabel metal2 s 76102 0 76158 800 6 la_oenb[33]
port 427 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_oenb[34]
port 428 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 la_oenb[35]
port 429 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 la_oenb[36]
port 430 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_oenb[37]
port 431 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 la_oenb[38]
port 432 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 la_oenb[39]
port 433 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 la_oenb[3]
port 434 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 la_oenb[40]
port 435 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 la_oenb[41]
port 436 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 la_oenb[42]
port 437 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 la_oenb[43]
port 438 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 la_oenb[44]
port 439 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 la_oenb[45]
port 440 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 la_oenb[46]
port 441 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_oenb[47]
port 442 nsew signal input
rlabel metal2 s 92662 0 92718 800 6 la_oenb[48]
port 443 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 la_oenb[49]
port 444 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 la_oenb[4]
port 445 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 la_oenb[50]
port 446 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 la_oenb[51]
port 447 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 la_oenb[52]
port 448 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 la_oenb[53]
port 449 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 la_oenb[54]
port 450 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 la_oenb[55]
port 451 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 la_oenb[56]
port 452 nsew signal input
rlabel metal2 s 102598 0 102654 800 6 la_oenb[57]
port 453 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 la_oenb[58]
port 454 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 la_oenb[59]
port 455 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 la_oenb[5]
port 456 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 la_oenb[60]
port 457 nsew signal input
rlabel metal2 s 107014 0 107070 800 6 la_oenb[61]
port 458 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 la_oenb[62]
port 459 nsew signal input
rlabel metal2 s 109222 0 109278 800 6 la_oenb[63]
port 460 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 la_oenb[64]
port 461 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 la_oenb[65]
port 462 nsew signal input
rlabel metal2 s 112534 0 112590 800 6 la_oenb[66]
port 463 nsew signal input
rlabel metal2 s 113638 0 113694 800 6 la_oenb[67]
port 464 nsew signal input
rlabel metal2 s 114742 0 114798 800 6 la_oenb[68]
port 465 nsew signal input
rlabel metal2 s 115846 0 115902 800 6 la_oenb[69]
port 466 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 la_oenb[6]
port 467 nsew signal input
rlabel metal2 s 116950 0 117006 800 6 la_oenb[70]
port 468 nsew signal input
rlabel metal2 s 118054 0 118110 800 6 la_oenb[71]
port 469 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 la_oenb[72]
port 470 nsew signal input
rlabel metal2 s 120170 0 120226 800 6 la_oenb[73]
port 471 nsew signal input
rlabel metal2 s 121274 0 121330 800 6 la_oenb[74]
port 472 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 la_oenb[75]
port 473 nsew signal input
rlabel metal2 s 123482 0 123538 800 6 la_oenb[76]
port 474 nsew signal input
rlabel metal2 s 124586 0 124642 800 6 la_oenb[77]
port 475 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 la_oenb[78]
port 476 nsew signal input
rlabel metal2 s 126794 0 126850 800 6 la_oenb[79]
port 477 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 la_oenb[7]
port 478 nsew signal input
rlabel metal2 s 127898 0 127954 800 6 la_oenb[80]
port 479 nsew signal input
rlabel metal2 s 129002 0 129058 800 6 la_oenb[81]
port 480 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 la_oenb[82]
port 481 nsew signal input
rlabel metal2 s 131210 0 131266 800 6 la_oenb[83]
port 482 nsew signal input
rlabel metal2 s 132314 0 132370 800 6 la_oenb[84]
port 483 nsew signal input
rlabel metal2 s 133418 0 133474 800 6 la_oenb[85]
port 484 nsew signal input
rlabel metal2 s 134522 0 134578 800 6 la_oenb[86]
port 485 nsew signal input
rlabel metal2 s 135626 0 135682 800 6 la_oenb[87]
port 486 nsew signal input
rlabel metal2 s 136730 0 136786 800 6 la_oenb[88]
port 487 nsew signal input
rlabel metal2 s 137834 0 137890 800 6 la_oenb[89]
port 488 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 la_oenb[8]
port 489 nsew signal input
rlabel metal2 s 138938 0 138994 800 6 la_oenb[90]
port 490 nsew signal input
rlabel metal2 s 140042 0 140098 800 6 la_oenb[91]
port 491 nsew signal input
rlabel metal2 s 141146 0 141202 800 6 la_oenb[92]
port 492 nsew signal input
rlabel metal2 s 142250 0 142306 800 6 la_oenb[93]
port 493 nsew signal input
rlabel metal2 s 143354 0 143410 800 6 la_oenb[94]
port 494 nsew signal input
rlabel metal2 s 144458 0 144514 800 6 la_oenb[95]
port 495 nsew signal input
rlabel metal2 s 145562 0 145618 800 6 la_oenb[96]
port 496 nsew signal input
rlabel metal2 s 146666 0 146722 800 6 la_oenb[97]
port 497 nsew signal input
rlabel metal2 s 147770 0 147826 800 6 la_oenb[98]
port 498 nsew signal input
rlabel metal2 s 148874 0 148930 800 6 la_oenb[99]
port 499 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_oenb[9]
port 500 nsew signal input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 501 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 502 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_ack_o
port 503 nsew signal tristate
rlabel metal2 s 2226 0 2282 800 6 wbs_adr_i[0]
port 504 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wbs_adr_i[10]
port 505 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 wbs_adr_i[11]
port 506 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_adr_i[12]
port 507 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_adr_i[13]
port 508 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_adr_i[14]
port 509 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 wbs_adr_i[15]
port 510 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_adr_i[16]
port 511 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_adr_i[17]
port 512 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 wbs_adr_i[18]
port 513 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 wbs_adr_i[19]
port 514 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[1]
port 515 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 wbs_adr_i[20]
port 516 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 wbs_adr_i[21]
port 517 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 wbs_adr_i[22]
port 518 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 wbs_adr_i[23]
port 519 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 wbs_adr_i[24]
port 520 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 wbs_adr_i[25]
port 521 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 wbs_adr_i[26]
port 522 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 wbs_adr_i[27]
port 523 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 wbs_adr_i[28]
port 524 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 wbs_adr_i[29]
port 525 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[2]
port 526 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 wbs_adr_i[30]
port 527 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 wbs_adr_i[31]
port 528 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_adr_i[3]
port 529 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_adr_i[4]
port 530 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_adr_i[5]
port 531 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_adr_i[6]
port 532 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_adr_i[7]
port 533 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_adr_i[8]
port 534 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_adr_i[9]
port 535 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_cyc_i
port 536 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_i[0]
port 537 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 wbs_dat_i[10]
port 538 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_i[11]
port 539 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 wbs_dat_i[12]
port 540 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 wbs_dat_i[13]
port 541 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_i[14]
port 542 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_i[15]
port 543 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wbs_dat_i[16]
port 544 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 wbs_dat_i[17]
port 545 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_i[18]
port 546 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wbs_dat_i[19]
port 547 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_dat_i[1]
port 548 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 wbs_dat_i[20]
port 549 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 wbs_dat_i[21]
port 550 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 wbs_dat_i[22]
port 551 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 wbs_dat_i[23]
port 552 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 wbs_dat_i[24]
port 553 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 wbs_dat_i[25]
port 554 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 wbs_dat_i[26]
port 555 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 wbs_dat_i[27]
port 556 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 wbs_dat_i[28]
port 557 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_i[29]
port 558 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_i[2]
port 559 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 wbs_dat_i[30]
port 560 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 wbs_dat_i[31]
port 561 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_dat_i[3]
port 562 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_i[4]
port 563 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_i[5]
port 564 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 wbs_dat_i[6]
port 565 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 wbs_dat_i[7]
port 566 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_i[8]
port 567 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_dat_i[9]
port 568 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_o[0]
port 569 nsew signal tristate
rlabel metal2 s 15474 0 15530 800 6 wbs_dat_o[10]
port 570 nsew signal tristate
rlabel metal2 s 16578 0 16634 800 6 wbs_dat_o[11]
port 571 nsew signal tristate
rlabel metal2 s 17682 0 17738 800 6 wbs_dat_o[12]
port 572 nsew signal tristate
rlabel metal2 s 18786 0 18842 800 6 wbs_dat_o[13]
port 573 nsew signal tristate
rlabel metal2 s 19890 0 19946 800 6 wbs_dat_o[14]
port 574 nsew signal tristate
rlabel metal2 s 20994 0 21050 800 6 wbs_dat_o[15]
port 575 nsew signal tristate
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_o[16]
port 576 nsew signal tristate
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_o[17]
port 577 nsew signal tristate
rlabel metal2 s 24306 0 24362 800 6 wbs_dat_o[18]
port 578 nsew signal tristate
rlabel metal2 s 25410 0 25466 800 6 wbs_dat_o[19]
port 579 nsew signal tristate
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_o[1]
port 580 nsew signal tristate
rlabel metal2 s 26514 0 26570 800 6 wbs_dat_o[20]
port 581 nsew signal tristate
rlabel metal2 s 27618 0 27674 800 6 wbs_dat_o[21]
port 582 nsew signal tristate
rlabel metal2 s 28722 0 28778 800 6 wbs_dat_o[22]
port 583 nsew signal tristate
rlabel metal2 s 29826 0 29882 800 6 wbs_dat_o[23]
port 584 nsew signal tristate
rlabel metal2 s 30930 0 30986 800 6 wbs_dat_o[24]
port 585 nsew signal tristate
rlabel metal2 s 32034 0 32090 800 6 wbs_dat_o[25]
port 586 nsew signal tristate
rlabel metal2 s 33138 0 33194 800 6 wbs_dat_o[26]
port 587 nsew signal tristate
rlabel metal2 s 34242 0 34298 800 6 wbs_dat_o[27]
port 588 nsew signal tristate
rlabel metal2 s 35346 0 35402 800 6 wbs_dat_o[28]
port 589 nsew signal tristate
rlabel metal2 s 36450 0 36506 800 6 wbs_dat_o[29]
port 590 nsew signal tristate
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_o[2]
port 591 nsew signal tristate
rlabel metal2 s 37554 0 37610 800 6 wbs_dat_o[30]
port 592 nsew signal tristate
rlabel metal2 s 38658 0 38714 800 6 wbs_dat_o[31]
port 593 nsew signal tristate
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_o[3]
port 594 nsew signal tristate
rlabel metal2 s 8850 0 8906 800 6 wbs_dat_o[4]
port 595 nsew signal tristate
rlabel metal2 s 9954 0 10010 800 6 wbs_dat_o[5]
port 596 nsew signal tristate
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_o[6]
port 597 nsew signal tristate
rlabel metal2 s 12162 0 12218 800 6 wbs_dat_o[7]
port 598 nsew signal tristate
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_o[8]
port 599 nsew signal tristate
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_o[9]
port 600 nsew signal tristate
rlabel metal2 s 3330 0 3386 800 6 wbs_sel_i[0]
port 601 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wbs_sel_i[1]
port 602 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_sel_i[2]
port 603 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_sel_i[3]
port 604 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_stb_i
port 605 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wbs_we_i
port 606 nsew signal input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 607 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 608 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 610 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 611 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 612 nsew power bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 613 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 614 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 615 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 616 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 617 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 618 nsew ground bidirectional
rlabel metal4 s 158468 2176 158788 117504 6 vccd2
port 619 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 117504 6 vccd2
port 620 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 117504 6 vccd2
port 621 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 117504 6 vccd2
port 622 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 117504 6 vccd2
port 623 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 117504 6 vccd2
port 624 nsew power bidirectional
rlabel metal4 s 173828 2176 174148 117504 6 vssd2
port 625 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 117504 6 vssd2
port 626 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 117504 6 vssd2
port 627 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 117504 6 vssd2
port 628 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 117504 6 vssd2
port 629 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 117504 6 vssd2
port 630 nsew ground bidirectional
rlabel metal4 s 159128 2176 159448 117504 6 vdda1
port 631 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 117504 6 vdda1
port 632 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 117504 6 vdda1
port 633 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 117504 6 vdda1
port 634 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 117504 6 vdda1
port 635 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 117504 6 vdda1
port 636 nsew power bidirectional
rlabel metal4 s 174488 2176 174808 117504 6 vssa1
port 637 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 117504 6 vssa1
port 638 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 117504 6 vssa1
port 639 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 117504 6 vssa1
port 640 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 117504 6 vssa1
port 641 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 117504 6 vssa1
port 642 nsew ground bidirectional
rlabel metal4 s 159788 2176 160108 117504 6 vdda2
port 643 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 117504 6 vdda2
port 644 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 117504 6 vdda2
port 645 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 117504 6 vdda2
port 646 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 117504 6 vdda2
port 647 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 117504 6 vdda2
port 648 nsew power bidirectional
rlabel metal4 s 175148 2176 175468 117504 6 vssa2
port 649 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 117504 6 vssa2
port 650 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 117504 6 vssa2
port 651 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 117504 6 vssa2
port 652 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 117504 6 vssa2
port 653 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 117504 6 vssa2
port 654 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 180000 120000
<< end >>
