VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO darkuart
  CLASS BLOCK ;
  FOREIGN darkuart ;
  ORIGIN 0.000 0.000 ;
  SIZE 113.430 BY 128.550 ;
  PIN BE[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.270 4.000 59.870 ;
    END
  END BE[0]
  PIN BE[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.670 4.000 30.270 ;
    END
  END BE[1]
  PIN BE[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.300 124.550 31.580 128.550 ;
    END
  END BE[2]
  PIN BE[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.300 0.000 103.580 4.000 ;
    END
  END BE[3]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.100 0.000 60.380 4.000 ;
    END
  END CLK
  PIN DATAI[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.270 4.000 96.870 ;
    END
  END DATAI[0]
  PIN DATAI[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.300 0.000 7.580 4.000 ;
    END
  END DATAI[10]
  PIN DATAI[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.700 0.000 45.980 4.000 ;
    END
  END DATAI[11]
  PIN DATAI[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.700 0.000 93.980 4.000 ;
    END
  END DATAI[12]
  PIN DATAI[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.430 11.170 113.430 11.770 ;
    END
  END DATAI[13]
  PIN DATAI[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.500 124.550 26.780 128.550 ;
    END
  END DATAI[14]
  PIN DATAI[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.300 124.550 7.580 128.550 ;
    END
  END DATAI[15]
  PIN DATAI[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.430 33.370 113.430 33.970 ;
    END
  END DATAI[16]
  PIN DATAI[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.430 25.970 113.430 26.570 ;
    END
  END DATAI[17]
  PIN DATAI[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.500 0.000 26.780 4.000 ;
    END
  END DATAI[18]
  PIN DATAI[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.430 85.170 113.430 85.770 ;
    END
  END DATAI[19]
  PIN DATAI[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.500 0.000 74.780 4.000 ;
    END
  END DATAI[1]
  PIN DATAI[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.100 0.000 12.380 4.000 ;
    END
  END DATAI[20]
  PIN DATAI[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.300 0.000 55.580 4.000 ;
    END
  END DATAI[21]
  PIN DATAI[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.500 0.000 98.780 4.000 ;
    END
  END DATAI[22]
  PIN DATAI[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.670 4.000 104.270 ;
    END
  END DATAI[23]
  PIN DATAI[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.900 124.550 89.180 128.550 ;
    END
  END DATAI[24]
  PIN DATAI[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.870 4.000 15.470 ;
    END
  END DATAI[25]
  PIN DATAI[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.500 124.550 2.780 128.550 ;
    END
  END DATAI[26]
  PIN DATAI[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.430 40.770 113.430 41.370 ;
    END
  END DATAI[27]
  PIN DATAI[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.900 124.550 41.180 128.550 ;
    END
  END DATAI[28]
  PIN DATAI[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.430 122.170 113.430 122.770 ;
    END
  END DATAI[29]
  PIN DATAI[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.900 0.000 41.180 4.000 ;
    END
  END DATAI[2]
  PIN DATAI[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.300 124.550 79.580 128.550 ;
    END
  END DATAI[30]
  PIN DATAI[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.100 0.000 36.380 4.000 ;
    END
  END DATAI[31]
  PIN DATAI[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.430 55.570 113.430 56.170 ;
    END
  END DATAI[3]
  PIN DATAI[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.470 4.000 45.070 ;
    END
  END DATAI[4]
  PIN DATAI[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.100 124.550 12.380 128.550 ;
    END
  END DATAI[5]
  PIN DATAI[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.070 4.000 111.670 ;
    END
  END DATAI[6]
  PIN DATAI[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.500 124.550 74.780 128.550 ;
    END
  END DATAI[7]
  PIN DATAI[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.430 114.770 113.430 115.370 ;
    END
  END DATAI[8]
  PIN DATAI[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.070 4.000 74.670 ;
    END
  END DATAI[9]
  PIN DATAO[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.870 4.000 52.470 ;
    END
  END DATAO[0]
  PIN DATAO[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.700 0.000 69.980 4.000 ;
    END
  END DATAO[10]
  PIN DATAO[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.470 4.000 119.070 ;
    END
  END DATAO[11]
  PIN DATAO[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.470 4.000 82.070 ;
    END
  END DATAO[12]
  PIN DATAO[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.870 4.000 89.470 ;
    END
  END DATAO[13]
  PIN DATAO[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.500 124.550 50.780 128.550 ;
    END
  END DATAO[14]
  PIN DATAO[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.430 3.770 113.430 4.370 ;
    END
  END DATAO[15]
  PIN DATAO[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.100 124.550 84.380 128.550 ;
    END
  END DATAO[16]
  PIN DATAO[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.500 0.000 50.780 4.000 ;
    END
  END DATAO[17]
  PIN DATAO[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.100 0.000 108.380 4.000 ;
    END
  END DATAO[18]
  PIN DATAO[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.900 0.000 89.180 4.000 ;
    END
  END DATAO[19]
  PIN DATAO[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.300 124.550 55.580 128.550 ;
    END
  END DATAO[1]
  PIN DATAO[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.700 0.000 21.980 4.000 ;
    END
  END DATAO[20]
  PIN DATAO[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.900 0.000 17.180 4.000 ;
    END
  END DATAO[21]
  PIN DATAO[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.300 0.000 79.580 4.000 ;
    END
  END DATAO[22]
  PIN DATAO[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.670 4.000 67.270 ;
    END
  END DATAO[23]
  PIN DATAO[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.500 0.000 2.780 4.000 ;
    END
  END DATAO[24]
  PIN DATAO[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.430 48.170 113.430 48.770 ;
    END
  END DATAO[25]
  PIN DATAO[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.300 124.550 103.580 128.550 ;
    END
  END DATAO[26]
  PIN DATAO[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.470 4.000 8.070 ;
    END
  END DATAO[27]
  PIN DATAO[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.270 4.000 22.870 ;
    END
  END DATAO[28]
  PIN DATAO[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.700 124.550 69.980 128.550 ;
    END
  END DATAO[29]
  PIN DATAO[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.900 124.550 17.180 128.550 ;
    END
  END DATAO[2]
  PIN DATAO[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.700 124.550 21.980 128.550 ;
    END
  END DATAO[30]
  PIN DATAO[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.700 124.550 45.980 128.550 ;
    END
  END DATAO[31]
  PIN DATAO[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.100 0.000 84.380 4.000 ;
    END
  END DATAO[3]
  PIN DATAO[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.430 107.370 113.430 107.970 ;
    END
  END DATAO[4]
  PIN DATAO[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.900 0.000 65.180 4.000 ;
    END
  END DATAO[5]
  PIN DATAO[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.430 77.770 113.430 78.370 ;
    END
  END DATAO[6]
  PIN DATAO[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.430 99.970 113.430 100.570 ;
    END
  END DATAO[7]
  PIN DATAO[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.900 124.550 65.180 128.550 ;
    END
  END DATAO[8]
  PIN DATAO[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.430 18.570 113.430 19.170 ;
    END
  END DATAO[9]
  PIN DEBUG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.430 92.570 113.430 93.170 ;
    END
  END DEBUG[0]
  PIN DEBUG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.300 0.000 31.580 4.000 ;
    END
  END DEBUG[1]
  PIN DEBUG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.100 124.550 36.380 128.550 ;
    END
  END DEBUG[2]
  PIN DEBUG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.070 4.000 37.670 ;
    END
  END DEBUG[3]
  PIN IRQ
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.100 124.550 60.380 128.550 ;
    END
  END IRQ
  PIN RD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.500 124.550 98.780 128.550 ;
    END
  END RD
  PIN RES
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.100 124.550 108.380 128.550 ;
    END
  END RES
  PIN RXD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.430 62.970 113.430 63.570 ;
    END
  END RXD
  PIN TXD
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.430 70.370 113.430 70.970 ;
    END
  END TXD
  PIN WR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.700 124.550 93.980 128.550 ;
    END
  END WR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 89.760 13.080 91.360 113.460 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 55.840 13.080 57.440 113.460 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.920 13.080 23.520 113.460 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 95.530 107.520 97.130 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 62.230 107.520 63.830 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 28.930 107.520 30.530 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 72.800 13.080 74.400 113.460 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 38.880 13.080 40.480 113.460 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 78.880 107.520 80.480 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 45.580 107.520 47.180 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.760 13.235 107.520 113.305 ;
      LAYER met1 ;
        RECT 2.480 13.075 108.400 113.465 ;
      LAYER met2 ;
        RECT 3.060 124.270 7.020 124.550 ;
        RECT 7.860 124.270 11.820 124.550 ;
        RECT 12.660 124.270 16.620 124.550 ;
        RECT 17.460 124.270 21.420 124.550 ;
        RECT 22.260 124.270 26.220 124.550 ;
        RECT 27.060 124.270 31.020 124.550 ;
        RECT 31.860 124.270 35.820 124.550 ;
        RECT 36.660 124.270 40.620 124.550 ;
        RECT 41.460 124.270 45.420 124.550 ;
        RECT 46.260 124.270 50.220 124.550 ;
        RECT 51.060 124.270 55.020 124.550 ;
        RECT 55.860 124.270 59.820 124.550 ;
        RECT 60.660 124.270 64.620 124.550 ;
        RECT 65.460 124.270 69.420 124.550 ;
        RECT 70.260 124.270 74.220 124.550 ;
        RECT 75.060 124.270 79.020 124.550 ;
        RECT 79.860 124.270 83.820 124.550 ;
        RECT 84.660 124.270 88.620 124.550 ;
        RECT 89.460 124.270 93.420 124.550 ;
        RECT 94.260 124.270 98.220 124.550 ;
        RECT 99.060 124.270 103.020 124.550 ;
        RECT 103.860 124.270 107.820 124.550 ;
        RECT 2.510 4.280 108.370 124.270 ;
        RECT 3.060 0.300 7.020 4.280 ;
        RECT 7.860 0.300 11.820 4.280 ;
        RECT 12.660 0.300 16.620 4.280 ;
        RECT 17.460 0.300 21.420 4.280 ;
        RECT 22.260 0.300 26.220 4.280 ;
        RECT 27.060 0.300 31.020 4.280 ;
        RECT 31.860 0.300 35.820 4.280 ;
        RECT 36.660 0.300 40.620 4.280 ;
        RECT 41.460 0.300 45.420 4.280 ;
        RECT 46.260 0.300 50.220 4.280 ;
        RECT 51.060 0.300 55.020 4.280 ;
        RECT 55.860 0.300 59.820 4.280 ;
        RECT 60.660 0.300 64.620 4.280 ;
        RECT 65.460 0.300 69.420 4.280 ;
        RECT 70.260 0.300 74.220 4.280 ;
        RECT 75.060 0.300 79.020 4.280 ;
        RECT 79.860 0.300 83.820 4.280 ;
        RECT 84.660 0.300 88.620 4.280 ;
        RECT 89.460 0.300 93.420 4.280 ;
        RECT 94.260 0.300 98.220 4.280 ;
        RECT 99.060 0.300 103.020 4.280 ;
        RECT 103.860 0.300 107.820 4.280 ;
      LAYER met3 ;
        RECT 4.000 121.770 109.030 122.635 ;
        RECT 4.000 119.470 109.430 121.770 ;
        RECT 4.400 118.070 109.430 119.470 ;
        RECT 4.000 115.770 109.430 118.070 ;
        RECT 4.000 114.370 109.030 115.770 ;
        RECT 4.000 112.070 109.430 114.370 ;
        RECT 4.400 110.670 109.430 112.070 ;
        RECT 4.000 108.370 109.430 110.670 ;
        RECT 4.000 106.970 109.030 108.370 ;
        RECT 4.000 104.670 109.430 106.970 ;
        RECT 4.400 103.270 109.430 104.670 ;
        RECT 4.000 100.970 109.430 103.270 ;
        RECT 4.000 99.570 109.030 100.970 ;
        RECT 4.000 97.270 109.430 99.570 ;
        RECT 4.400 95.870 109.430 97.270 ;
        RECT 4.000 93.570 109.430 95.870 ;
        RECT 4.000 92.170 109.030 93.570 ;
        RECT 4.000 89.870 109.430 92.170 ;
        RECT 4.400 88.470 109.430 89.870 ;
        RECT 4.000 86.170 109.430 88.470 ;
        RECT 4.000 84.770 109.030 86.170 ;
        RECT 4.000 82.470 109.430 84.770 ;
        RECT 4.400 81.070 109.430 82.470 ;
        RECT 4.000 78.770 109.430 81.070 ;
        RECT 4.000 77.370 109.030 78.770 ;
        RECT 4.000 75.070 109.430 77.370 ;
        RECT 4.400 73.670 109.430 75.070 ;
        RECT 4.000 71.370 109.430 73.670 ;
        RECT 4.000 69.970 109.030 71.370 ;
        RECT 4.000 67.670 109.430 69.970 ;
        RECT 4.400 66.270 109.430 67.670 ;
        RECT 4.000 63.970 109.430 66.270 ;
        RECT 4.000 62.570 109.030 63.970 ;
        RECT 4.000 60.270 109.430 62.570 ;
        RECT 4.400 58.870 109.430 60.270 ;
        RECT 4.000 56.570 109.430 58.870 ;
        RECT 4.000 55.170 109.030 56.570 ;
        RECT 4.000 52.870 109.430 55.170 ;
        RECT 4.400 51.470 109.430 52.870 ;
        RECT 4.000 49.170 109.430 51.470 ;
        RECT 4.000 47.770 109.030 49.170 ;
        RECT 4.000 45.470 109.430 47.770 ;
        RECT 4.400 44.070 109.430 45.470 ;
        RECT 4.000 41.770 109.430 44.070 ;
        RECT 4.000 40.370 109.030 41.770 ;
        RECT 4.000 38.070 109.430 40.370 ;
        RECT 4.400 36.670 109.430 38.070 ;
        RECT 4.000 34.370 109.430 36.670 ;
        RECT 4.000 32.970 109.030 34.370 ;
        RECT 4.000 30.670 109.430 32.970 ;
        RECT 4.400 29.270 109.430 30.670 ;
        RECT 4.000 26.970 109.430 29.270 ;
        RECT 4.000 25.570 109.030 26.970 ;
        RECT 4.000 23.270 109.430 25.570 ;
        RECT 4.400 21.870 109.430 23.270 ;
        RECT 4.000 19.570 109.430 21.870 ;
        RECT 4.000 18.170 109.030 19.570 ;
        RECT 4.000 15.870 109.430 18.170 ;
        RECT 4.400 14.470 109.430 15.870 ;
        RECT 4.000 12.170 109.430 14.470 ;
        RECT 4.000 10.770 109.030 12.170 ;
        RECT 4.000 8.470 109.430 10.770 ;
        RECT 4.400 7.070 109.430 8.470 ;
        RECT 4.000 4.770 109.430 7.070 ;
        RECT 4.000 3.905 109.030 4.770 ;
  END
END darkuart
END LIBRARY

